magic
tech sky130B
magscale 1 2
timestamp 1668086266
<< viali >>
rect 5273 57409 5307 57443
rect 15209 57409 15243 57443
rect 25145 57409 25179 57443
rect 35081 57409 35115 57443
rect 45017 57409 45051 57443
rect 55321 57409 55355 57443
rect 64889 57409 64923 57443
rect 67005 57409 67039 57443
rect 67649 57409 67683 57443
rect 68109 56797 68143 56831
rect 67649 55097 67683 55131
rect 67649 53941 67683 53975
rect 68109 52445 68143 52479
rect 68109 51357 68143 51391
rect 67649 49725 67683 49759
rect 67649 48501 67683 48535
rect 68109 47005 68143 47039
rect 68109 45917 68143 45951
rect 67649 44217 67683 44251
rect 67649 43061 67683 43095
rect 68109 41565 68143 41599
rect 68109 40477 68143 40511
rect 67649 38777 67683 38811
rect 67649 37621 67683 37655
rect 68109 36125 68143 36159
rect 68109 35037 68143 35071
rect 67649 33337 67683 33371
rect 67649 32181 67683 32215
rect 15761 31705 15795 31739
rect 17785 31637 17819 31671
rect 8769 31365 8803 31399
rect 12449 31365 12483 31399
rect 15025 31365 15059 31399
rect 21833 31365 21867 31399
rect 23489 31365 23523 31399
rect 23673 31365 23707 31399
rect 8585 31297 8619 31331
rect 12081 31297 12115 31331
rect 12265 31297 12299 31331
rect 12909 31297 12943 31331
rect 13072 31300 13106 31334
rect 13185 31297 13219 31331
rect 13323 31297 13357 31331
rect 15209 31297 15243 31331
rect 15945 31297 15979 31331
rect 17049 31297 17083 31331
rect 17233 31297 17267 31331
rect 17325 31297 17359 31331
rect 17417 31297 17451 31331
rect 20545 31297 20579 31331
rect 20637 31297 20671 31331
rect 20729 31297 20763 31331
rect 20913 31297 20947 31331
rect 23305 31297 23339 31331
rect 24133 31297 24167 31331
rect 24317 31297 24351 31331
rect 24409 31297 24443 31331
rect 24501 31297 24535 31331
rect 14105 31161 14139 31195
rect 18153 31161 18187 31195
rect 8953 31093 8987 31127
rect 13553 31093 13587 31127
rect 15393 31093 15427 31127
rect 17693 31093 17727 31127
rect 20269 31093 20303 31127
rect 24777 31093 24811 31127
rect 10333 30889 10367 30923
rect 17509 30889 17543 30923
rect 20269 30889 20303 30923
rect 16681 30753 16715 30787
rect 8401 30685 8435 30719
rect 9367 30685 9401 30719
rect 9505 30685 9539 30719
rect 9602 30682 9636 30716
rect 9781 30685 9815 30719
rect 11601 30685 11635 30719
rect 11713 30685 11747 30719
rect 11810 30685 11844 30719
rect 11989 30685 12023 30719
rect 15209 30685 15243 30719
rect 15301 30685 15335 30719
rect 15393 30685 15427 30719
rect 15577 30685 15611 30719
rect 16037 30685 16071 30719
rect 16221 30685 16255 30719
rect 16313 30685 16347 30719
rect 16405 30685 16439 30719
rect 20453 30685 20487 30719
rect 68109 30685 68143 30719
rect 8217 30617 8251 30651
rect 17141 30617 17175 30651
rect 17325 30617 17359 30651
rect 20637 30617 20671 30651
rect 8033 30549 8067 30583
rect 9137 30549 9171 30583
rect 11345 30549 11379 30583
rect 12449 30549 12483 30583
rect 14933 30549 14967 30583
rect 18061 30549 18095 30583
rect 24409 30549 24443 30583
rect 5825 30345 5859 30379
rect 11897 30345 11931 30379
rect 15669 30345 15703 30379
rect 7104 30277 7138 30311
rect 11713 30277 11747 30311
rect 13746 30277 13780 30311
rect 15485 30277 15519 30311
rect 18622 30277 18656 30311
rect 19616 30277 19650 30311
rect 23673 30277 23707 30311
rect 4445 30209 4479 30243
rect 4712 30209 4746 30243
rect 9229 30209 9263 30243
rect 9318 30212 9352 30246
rect 9413 30209 9447 30243
rect 9597 30209 9631 30243
rect 11529 30209 11563 30243
rect 15301 30209 15335 30243
rect 18889 30209 18923 30243
rect 19349 30209 19383 30243
rect 22089 30209 22123 30243
rect 23857 30209 23891 30243
rect 26166 30209 26200 30243
rect 26433 30209 26467 30243
rect 28181 30209 28215 30243
rect 28437 30209 28471 30243
rect 6837 30141 6871 30175
rect 14013 30141 14047 30175
rect 21833 30141 21867 30175
rect 8953 30073 8987 30107
rect 10149 30073 10183 30107
rect 17049 30073 17083 30107
rect 25053 30073 25087 30107
rect 8217 30005 8251 30039
rect 12633 30005 12667 30039
rect 17509 30005 17543 30039
rect 20729 30005 20763 30039
rect 23213 30005 23247 30039
rect 24041 30005 24075 30039
rect 29561 30005 29595 30039
rect 10425 29801 10459 29835
rect 17325 29801 17359 29835
rect 20729 29801 20763 29835
rect 21833 29801 21867 29835
rect 3801 29665 3835 29699
rect 22293 29665 22327 29699
rect 11805 29597 11839 29631
rect 12541 29597 12575 29631
rect 12633 29597 12667 29631
rect 12725 29597 12759 29631
rect 12909 29597 12943 29631
rect 16589 29597 16623 29631
rect 18705 29597 18739 29631
rect 21189 29597 21223 29631
rect 21352 29597 21386 29631
rect 21452 29597 21486 29631
rect 21557 29597 21591 29631
rect 22477 29597 22511 29631
rect 22661 29597 22695 29631
rect 23489 29597 23523 29631
rect 23594 29591 23628 29625
rect 23694 29597 23728 29631
rect 23857 29597 23891 29631
rect 24961 29597 24995 29631
rect 28181 29597 28215 29631
rect 68109 29597 68143 29631
rect 4046 29529 4080 29563
rect 11538 29529 11572 29563
rect 13461 29529 13495 29563
rect 16322 29529 16356 29563
rect 18438 29529 18472 29563
rect 25228 29529 25262 29563
rect 27914 29529 27948 29563
rect 5181 29461 5215 29495
rect 12265 29461 12299 29495
rect 15209 29461 15243 29495
rect 23213 29461 23247 29495
rect 24409 29461 24443 29495
rect 26341 29461 26375 29495
rect 26801 29461 26835 29495
rect 7757 29257 7791 29291
rect 12173 29257 12207 29291
rect 13001 29257 13035 29291
rect 15025 29257 15059 29291
rect 17601 29257 17635 29291
rect 11805 29189 11839 29223
rect 12817 29189 12851 29223
rect 16681 29189 16715 29223
rect 20637 29189 20671 29223
rect 28917 29189 28951 29223
rect 6377 29121 6411 29155
rect 6644 29121 6678 29155
rect 10793 29121 10827 29155
rect 11529 29121 11563 29155
rect 11677 29121 11711 29155
rect 11897 29121 11931 29155
rect 11994 29121 12028 29155
rect 12633 29121 12667 29155
rect 13645 29121 13679 29155
rect 13912 29121 13946 29155
rect 16865 29121 16899 29155
rect 20821 29121 20855 29155
rect 23213 29121 23247 29155
rect 23469 29121 23503 29155
rect 29101 29121 29135 29155
rect 30858 29121 30892 29155
rect 31125 29121 31159 29155
rect 33250 29121 33284 29155
rect 33517 29121 33551 29155
rect 9505 28985 9539 29019
rect 21925 28985 21959 29019
rect 24593 28985 24627 29019
rect 27905 28985 27939 29019
rect 29745 28985 29779 29019
rect 8217 28917 8251 28951
rect 17049 28917 17083 28951
rect 21005 28917 21039 28951
rect 28733 28917 28767 28951
rect 32137 28917 32171 28951
rect 6561 28713 6595 28747
rect 8401 28713 8435 28747
rect 16221 28713 16255 28747
rect 22201 28713 22235 28747
rect 27537 28713 27571 28747
rect 28273 28713 28307 28747
rect 30941 28713 30975 28747
rect 9505 28645 9539 28679
rect 17325 28645 17359 28679
rect 15761 28577 15795 28611
rect 21097 28577 21131 28611
rect 22753 28577 22787 28611
rect 4077 28509 4111 28543
rect 6837 28509 6871 28543
rect 6929 28509 6963 28543
rect 7021 28509 7055 28543
rect 7205 28509 7239 28543
rect 7849 28509 7883 28543
rect 8125 28509 8159 28543
rect 8217 28509 8251 28543
rect 10885 28509 10919 28543
rect 12173 28509 12207 28543
rect 12266 28509 12300 28543
rect 12403 28509 12437 28543
rect 12541 28509 12575 28543
rect 12679 28509 12713 28543
rect 15393 28509 15427 28543
rect 16451 28509 16485 28543
rect 16589 28509 16623 28543
rect 16681 28509 16715 28543
rect 16865 28509 16899 28543
rect 18705 28509 18739 28543
rect 22017 28509 22051 28543
rect 23489 28509 23523 28543
rect 23594 28506 23628 28540
rect 23694 28506 23728 28540
rect 23857 28509 23891 28543
rect 28549 28509 28583 28543
rect 28641 28509 28675 28543
rect 28733 28509 28767 28543
rect 28917 28509 28951 28543
rect 30297 28509 30331 28543
rect 30481 28509 30515 28543
rect 30573 28509 30607 28543
rect 30711 28509 30745 28543
rect 1961 28441 1995 28475
rect 2145 28441 2179 28475
rect 4322 28441 4356 28475
rect 8033 28441 8067 28475
rect 10640 28441 10674 28475
rect 15577 28441 15611 28475
rect 18438 28441 18472 28475
rect 20830 28441 20864 28475
rect 25237 28441 25271 28475
rect 25421 28441 25455 28475
rect 26065 28441 26099 28475
rect 2329 28373 2363 28407
rect 5457 28373 5491 28407
rect 8953 28373 8987 28407
rect 11345 28373 11379 28407
rect 12817 28373 12851 28407
rect 19717 28373 19751 28407
rect 23213 28373 23247 28407
rect 25605 28373 25639 28407
rect 29745 28373 29779 28407
rect 3249 28169 3283 28203
rect 6837 28169 6871 28203
rect 9505 28169 9539 28203
rect 10701 28169 10735 28203
rect 16037 28169 16071 28203
rect 17877 28169 17911 28203
rect 20637 28169 20671 28203
rect 25237 28169 25271 28203
rect 26341 28169 26375 28203
rect 27629 28169 27663 28203
rect 28181 28169 28215 28203
rect 30481 28169 30515 28203
rect 1961 28101 1995 28135
rect 9229 28101 9263 28135
rect 10333 28101 10367 28135
rect 11897 28101 11931 28135
rect 11989 28101 12023 28135
rect 22201 28101 22235 28135
rect 22385 28101 22419 28135
rect 23112 28101 23146 28135
rect 29377 28101 29411 28135
rect 1777 28033 1811 28067
rect 2605 28033 2639 28067
rect 2789 28033 2823 28067
rect 2881 28033 2915 28067
rect 3019 28033 3053 28067
rect 3709 28033 3743 28067
rect 5641 28033 5675 28067
rect 5825 28033 5859 28067
rect 6469 28033 6503 28067
rect 6653 28033 6687 28067
rect 7757 28033 7791 28067
rect 7941 28033 7975 28067
rect 8953 28033 8987 28067
rect 9137 28033 9171 28067
rect 9321 28033 9355 28067
rect 10149 28033 10183 28067
rect 10425 28033 10459 28067
rect 10517 28033 10551 28067
rect 11621 28033 11655 28067
rect 11714 28033 11748 28067
rect 12086 28033 12120 28067
rect 13277 28033 13311 28067
rect 15126 28033 15160 28067
rect 15853 28033 15887 28067
rect 17233 28033 17267 28067
rect 17417 28033 17451 28067
rect 17509 28033 17543 28067
rect 17601 28033 17635 28067
rect 18337 28033 18371 28067
rect 19073 28033 19107 28067
rect 19809 28033 19843 28067
rect 20913 28033 20947 28067
rect 21005 28033 21039 28067
rect 21097 28033 21131 28067
rect 21281 28033 21315 28067
rect 25513 28033 25547 28067
rect 25605 28033 25639 28067
rect 25697 28033 25731 28067
rect 25881 28033 25915 28067
rect 26985 28033 27019 28067
rect 27169 28033 27203 28067
rect 27261 28033 27295 28067
rect 27353 28033 27387 28067
rect 28733 28033 28767 28067
rect 28896 28033 28930 28067
rect 28996 28039 29030 28073
rect 29147 28033 29181 28067
rect 29837 28033 29871 28067
rect 30665 28033 30699 28067
rect 30849 28033 30883 28067
rect 33250 28033 33284 28067
rect 33517 28033 33551 28067
rect 2145 27965 2179 27999
rect 13553 27965 13587 27999
rect 15393 27965 15427 27999
rect 19625 27965 19659 27999
rect 22845 27965 22879 27999
rect 67649 27897 67683 27931
rect 5457 27829 5491 27863
rect 8125 27829 8159 27863
rect 12265 27829 12299 27863
rect 14013 27829 14047 27863
rect 24225 27829 24259 27863
rect 24777 27829 24811 27863
rect 32137 27829 32171 27863
rect 14749 27625 14783 27659
rect 20453 27625 20487 27659
rect 24409 27625 24443 27659
rect 1593 27557 1627 27591
rect 2697 27557 2731 27591
rect 5273 27557 5307 27591
rect 10333 27557 10367 27591
rect 11529 27557 11563 27591
rect 17141 27557 17175 27591
rect 21465 27557 21499 27591
rect 25237 27557 25271 27591
rect 26157 27557 26191 27591
rect 30757 27557 30791 27591
rect 6653 27489 6687 27523
rect 16221 27489 16255 27523
rect 22293 27489 22327 27523
rect 27813 27489 27847 27523
rect 2053 27421 2087 27455
rect 2237 27421 2271 27455
rect 2329 27421 2363 27455
rect 2421 27421 2455 27455
rect 7205 27421 7239 27455
rect 7757 27421 7791 27455
rect 7941 27421 7975 27455
rect 8033 27421 8067 27455
rect 8171 27421 8205 27455
rect 8953 27421 8987 27455
rect 10885 27421 10919 27455
rect 11033 27421 11067 27455
rect 11391 27421 11425 27455
rect 12725 27421 12759 27455
rect 13369 27421 13403 27455
rect 14105 27421 14139 27455
rect 14289 27421 14323 27455
rect 14381 27421 14415 27455
rect 14473 27421 14507 27455
rect 16497 27421 16531 27455
rect 18245 27421 18279 27455
rect 18521 27421 18555 27455
rect 21281 27421 21315 27455
rect 22017 27421 22051 27455
rect 25973 27421 26007 27455
rect 28089 27421 28123 27455
rect 30113 27421 30147 27455
rect 30297 27421 30331 27455
rect 30389 27421 30423 27455
rect 30481 27421 30515 27455
rect 6408 27353 6442 27387
rect 8401 27353 8435 27387
rect 9198 27353 9232 27387
rect 11161 27353 11195 27387
rect 11253 27353 11287 27387
rect 13185 27353 13219 27387
rect 13553 27353 13587 27387
rect 19257 27353 19291 27387
rect 19441 27353 19475 27387
rect 24593 27353 24627 27387
rect 24777 27353 24811 27387
rect 25789 27353 25823 27387
rect 29561 27353 29595 27387
rect 12541 27285 12575 27319
rect 19625 27285 19659 27319
rect 26709 27285 26743 27319
rect 6561 27081 6595 27115
rect 10885 27081 10919 27115
rect 16129 27081 16163 27115
rect 20453 27081 20487 27115
rect 23121 27081 23155 27115
rect 29377 27081 29411 27115
rect 30389 27081 30423 27115
rect 2973 27013 3007 27047
rect 3678 27013 3712 27047
rect 10517 27013 10551 27047
rect 18153 27013 18187 27047
rect 22017 27013 22051 27047
rect 23765 27013 23799 27047
rect 26433 27013 26467 27047
rect 29009 27013 29043 27047
rect 30021 27013 30055 27047
rect 2329 26945 2363 26979
rect 2513 26945 2547 26979
rect 2605 26945 2639 26979
rect 2697 26945 2731 26979
rect 3433 26945 3467 26979
rect 6837 26945 6871 26979
rect 6929 26945 6963 26979
rect 7021 26945 7055 26979
rect 7205 26945 7239 26979
rect 7665 26945 7699 26979
rect 10333 26945 10367 26979
rect 10609 26945 10643 26979
rect 10701 26945 10735 26979
rect 12725 26945 12759 26979
rect 14197 26945 14231 26979
rect 15945 26945 15979 26979
rect 20545 26945 20579 26979
rect 21097 26945 21131 26979
rect 21833 26945 21867 26979
rect 23949 26945 23983 26979
rect 24961 26945 24995 26979
rect 25237 26945 25271 26979
rect 25795 26945 25829 26979
rect 25952 26945 25986 26979
rect 26065 26945 26099 26979
rect 26177 26945 26211 26979
rect 28282 26945 28316 26979
rect 28549 26945 28583 26979
rect 29193 26945 29227 26979
rect 30205 26945 30239 26979
rect 12081 26877 12115 26911
rect 12541 26877 12575 26911
rect 13921 26877 13955 26911
rect 16681 26877 16715 26911
rect 16957 26877 16991 26911
rect 4813 26741 4847 26775
rect 12909 26741 12943 26775
rect 14933 26741 14967 26775
rect 19441 26741 19475 26775
rect 22201 26741 22235 26775
rect 23581 26741 23615 26775
rect 27169 26741 27203 26775
rect 30941 26741 30975 26775
rect 67649 26741 67683 26775
rect 2605 26537 2639 26571
rect 5181 26537 5215 26571
rect 8217 26537 8251 26571
rect 14197 26537 14231 26571
rect 26617 26537 26651 26571
rect 27721 26537 27755 26571
rect 10793 26469 10827 26503
rect 21005 26469 21039 26503
rect 24409 26469 24443 26503
rect 28457 26469 28491 26503
rect 3801 26401 3835 26435
rect 19993 26401 20027 26435
rect 22385 26401 22419 26435
rect 25789 26401 25823 26435
rect 33149 26401 33183 26435
rect 2421 26333 2455 26367
rect 6837 26333 6871 26367
rect 10241 26333 10275 26367
rect 10517 26333 10551 26367
rect 10609 26333 10643 26367
rect 12357 26333 12391 26367
rect 12449 26333 12483 26367
rect 12541 26333 12575 26367
rect 12725 26333 12759 26367
rect 13185 26333 13219 26367
rect 14105 26333 14139 26367
rect 14289 26333 14323 26367
rect 14749 26333 14783 26367
rect 15025 26333 15059 26367
rect 16037 26333 16071 26367
rect 16221 26333 16255 26367
rect 17325 26333 17359 26367
rect 17509 26333 17543 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 18337 26333 18371 26367
rect 18429 26333 18463 26367
rect 19717 26333 19751 26367
rect 23213 26333 23247 26367
rect 23376 26330 23410 26364
rect 23476 26333 23510 26367
rect 23601 26333 23635 26367
rect 29009 26333 29043 26367
rect 29837 26333 29871 26367
rect 29929 26333 29963 26367
rect 30021 26333 30055 26367
rect 30205 26333 30239 26367
rect 30665 26333 30699 26367
rect 30849 26333 30883 26367
rect 30941 26333 30975 26367
rect 31033 26333 31067 26367
rect 2237 26265 2271 26299
rect 4046 26265 4080 26299
rect 7082 26265 7116 26299
rect 10425 26265 10459 26299
rect 12081 26265 12115 26299
rect 16865 26265 16899 26299
rect 18705 26265 18739 26299
rect 22118 26265 22152 26299
rect 23857 26265 23891 26299
rect 25522 26265 25556 26299
rect 26249 26265 26283 26299
rect 26433 26265 26467 26299
rect 27077 26265 27111 26299
rect 28273 26265 28307 26299
rect 31309 26265 31343 26299
rect 32882 26265 32916 26299
rect 13369 26197 13403 26231
rect 16221 26197 16255 26231
rect 29561 26197 29595 26231
rect 31769 26197 31803 26231
rect 3249 25993 3283 26027
rect 12909 25993 12943 26027
rect 22201 25993 22235 26027
rect 25973 25993 26007 26027
rect 31493 25993 31527 26027
rect 34897 25993 34931 26027
rect 1777 25925 1811 25959
rect 1961 25925 1995 25959
rect 8484 25925 8518 25959
rect 11529 25925 11563 25959
rect 15209 25925 15243 25959
rect 15761 25925 15795 25959
rect 29552 25925 29586 25959
rect 2605 25857 2639 25891
rect 2789 25857 2823 25891
rect 2881 25857 2915 25891
rect 3019 25857 3053 25891
rect 3801 25857 3835 25891
rect 5825 25857 5859 25891
rect 6653 25857 6687 25891
rect 6745 25857 6779 25891
rect 6837 25857 6871 25891
rect 7021 25857 7055 25891
rect 8217 25857 8251 25891
rect 11713 25857 11747 25891
rect 13829 25857 13863 25891
rect 15025 25857 15059 25891
rect 15945 25857 15979 25891
rect 18346 25857 18380 25891
rect 19513 25857 19547 25891
rect 21281 25857 21315 25891
rect 22477 25857 22511 25891
rect 22569 25857 22603 25891
rect 22661 25857 22695 25891
rect 22845 25857 22879 25891
rect 23581 25857 23615 25891
rect 24685 25857 24719 25891
rect 27997 25857 28031 25891
rect 29285 25857 29319 25891
rect 31125 25857 31159 25891
rect 31309 25857 31343 25891
rect 32505 25857 32539 25891
rect 32689 25857 32723 25891
rect 32781 25857 32815 25891
rect 32873 25857 32907 25891
rect 33609 25857 33643 25891
rect 2145 25789 2179 25823
rect 11897 25789 11931 25823
rect 13553 25789 13587 25823
rect 14841 25789 14875 25823
rect 18613 25789 18647 25823
rect 19257 25789 19291 25823
rect 23305 25789 23339 25823
rect 28273 25789 28307 25823
rect 9597 25721 9631 25755
rect 17233 25721 17267 25755
rect 6377 25653 6411 25687
rect 16129 25653 16163 25687
rect 20637 25653 20671 25687
rect 27077 25653 27111 25687
rect 30665 25653 30699 25687
rect 33149 25653 33183 25687
rect 5733 25449 5767 25483
rect 6745 25449 6779 25483
rect 16681 25449 16715 25483
rect 20637 25449 20671 25483
rect 21925 25449 21959 25483
rect 31309 25449 31343 25483
rect 32781 25449 32815 25483
rect 18705 25381 18739 25415
rect 26249 25381 26283 25415
rect 26801 25381 26835 25415
rect 4353 25313 4387 25347
rect 10517 25313 10551 25347
rect 28181 25313 28215 25347
rect 29837 25313 29871 25347
rect 35449 25313 35483 25347
rect 2605 25245 2639 25279
rect 2789 25245 2823 25279
rect 2881 25245 2915 25279
rect 3019 25245 3053 25279
rect 3893 25245 3927 25279
rect 6929 25245 6963 25279
rect 14289 25245 14323 25279
rect 16037 25245 16071 25279
rect 16221 25245 16255 25279
rect 16313 25245 16347 25279
rect 16451 25245 16485 25279
rect 17601 25245 17635 25279
rect 17785 25245 17819 25279
rect 19257 25245 19291 25279
rect 21741 25245 21775 25279
rect 22385 25245 22419 25279
rect 22569 25245 22603 25279
rect 22661 25245 22695 25279
rect 22799 25245 22833 25279
rect 25513 25245 25547 25279
rect 25789 25245 25823 25279
rect 29561 25245 29595 25279
rect 31677 25245 31711 25279
rect 35705 25245 35739 25279
rect 68109 25245 68143 25279
rect 3249 25177 3283 25211
rect 4598 25177 4632 25211
rect 7113 25177 7147 25211
rect 10784 25177 10818 25211
rect 14105 25177 14139 25211
rect 14933 25177 14967 25211
rect 19502 25177 19536 25211
rect 21281 25177 21315 25211
rect 23489 25177 23523 25211
rect 23673 25177 23707 25211
rect 27914 25177 27948 25211
rect 31493 25177 31527 25211
rect 32413 25177 32447 25211
rect 32597 25177 32631 25211
rect 11897 25109 11931 25143
rect 13461 25109 13495 25143
rect 14473 25109 14507 25143
rect 17969 25109 18003 25143
rect 23029 25109 23063 25143
rect 23857 25109 23891 25143
rect 33517 25109 33551 25143
rect 36829 25109 36863 25143
rect 2881 24905 2915 24939
rect 22201 24905 22235 24939
rect 24777 24905 24811 24939
rect 31125 24905 31159 24939
rect 32413 24905 32447 24939
rect 2513 24837 2547 24871
rect 19257 24837 19291 24871
rect 2697 24769 2731 24803
rect 4169 24769 4203 24803
rect 6561 24769 6595 24803
rect 8401 24769 8435 24803
rect 8668 24769 8702 24803
rect 11805 24769 11839 24803
rect 11897 24769 11931 24803
rect 11989 24769 12023 24803
rect 12173 24769 12207 24803
rect 13553 24769 13587 24803
rect 13645 24769 13679 24803
rect 13737 24769 13771 24803
rect 13921 24769 13955 24803
rect 15862 24769 15896 24803
rect 16865 24769 16899 24803
rect 17969 24769 18003 24803
rect 18153 24769 18187 24803
rect 18245 24769 18279 24803
rect 18337 24769 18371 24803
rect 19441 24769 19475 24803
rect 19993 24769 20027 24803
rect 20177 24769 20211 24803
rect 21097 24769 21131 24803
rect 21833 24769 21867 24803
rect 22017 24769 22051 24803
rect 23958 24769 23992 24803
rect 24225 24769 24259 24803
rect 25329 24769 25363 24803
rect 25513 24769 25547 24803
rect 25605 24769 25639 24803
rect 25697 24769 25731 24803
rect 26985 24769 27019 24803
rect 27169 24769 27203 24803
rect 27261 24769 27295 24803
rect 27353 24769 27387 24803
rect 28089 24769 28123 24803
rect 30297 24769 30331 24803
rect 30941 24769 30975 24803
rect 33057 24769 33091 24803
rect 33241 24769 33275 24803
rect 33333 24769 33367 24803
rect 33425 24769 33459 24803
rect 34713 24769 34747 24803
rect 34969 24769 35003 24803
rect 7665 24701 7699 24735
rect 7941 24701 7975 24735
rect 11529 24701 11563 24735
rect 13277 24701 13311 24735
rect 16129 24701 16163 24735
rect 18613 24701 18647 24735
rect 25973 24701 26007 24735
rect 33701 24701 33735 24735
rect 4353 24633 4387 24667
rect 6377 24633 6411 24667
rect 12725 24633 12759 24667
rect 21281 24633 21315 24667
rect 30481 24633 30515 24667
rect 4905 24565 4939 24599
rect 9781 24565 9815 24599
rect 14749 24565 14783 24599
rect 22845 24565 22879 24599
rect 27629 24565 27663 24599
rect 36093 24565 36127 24599
rect 1777 24361 1811 24395
rect 3019 24361 3053 24395
rect 9413 24361 9447 24395
rect 13185 24361 13219 24395
rect 14841 24361 14875 24395
rect 23397 24361 23431 24395
rect 25421 24361 25455 24395
rect 31769 24361 31803 24395
rect 33149 24361 33183 24395
rect 25881 24293 25915 24327
rect 33609 24293 33643 24327
rect 21373 24225 21407 24259
rect 22845 24225 22879 24259
rect 27813 24225 27847 24259
rect 1961 24157 1995 24191
rect 3249 24157 3283 24191
rect 3801 24157 3835 24191
rect 3985 24157 4019 24191
rect 4077 24157 4111 24191
rect 4169 24157 4203 24191
rect 4905 24157 4939 24191
rect 9597 24157 9631 24191
rect 10241 24157 10275 24191
rect 10609 24157 10643 24191
rect 13001 24157 13035 24191
rect 14185 24157 14219 24191
rect 14381 24157 14415 24191
rect 14473 24157 14507 24191
rect 14565 24157 14599 24191
rect 17141 24157 17175 24191
rect 19257 24157 19291 24191
rect 19441 24157 19475 24191
rect 19533 24157 19567 24191
rect 19625 24157 19659 24191
rect 21281 24157 21315 24191
rect 21465 24157 21499 24191
rect 22569 24157 22603 24191
rect 23305 24157 23339 24191
rect 23489 24157 23523 24191
rect 25053 24157 25087 24191
rect 27546 24157 27580 24191
rect 28365 24157 28399 24191
rect 28549 24157 28583 24191
rect 28641 24157 28675 24191
rect 28733 24157 28767 24191
rect 29561 24157 29595 24191
rect 68109 24157 68143 24191
rect 5549 24089 5583 24123
rect 7757 24089 7791 24123
rect 9781 24089 9815 24123
rect 10425 24089 10459 24123
rect 10517 24089 10551 24123
rect 12817 24089 12851 24123
rect 15301 24089 15335 24123
rect 16957 24089 16991 24123
rect 25237 24089 25271 24123
rect 29009 24089 29043 24123
rect 29806 24089 29840 24123
rect 31401 24089 31435 24123
rect 31585 24089 31619 24123
rect 32781 24089 32815 24123
rect 32965 24089 32999 24123
rect 4445 24021 4479 24055
rect 6837 24021 6871 24055
rect 10793 24021 10827 24055
rect 11345 24021 11379 24055
rect 17325 24021 17359 24055
rect 18153 24021 18187 24055
rect 18705 24021 18739 24055
rect 19901 24021 19935 24055
rect 20361 24021 20395 24055
rect 24409 24021 24443 24055
rect 26433 24021 26467 24055
rect 30941 24021 30975 24055
rect 32229 24021 32263 24055
rect 5733 23817 5767 23851
rect 8769 23817 8803 23851
rect 14749 23817 14783 23851
rect 18613 23817 18647 23851
rect 20729 23817 20763 23851
rect 22293 23817 22327 23851
rect 28181 23817 28215 23851
rect 36737 23817 36771 23851
rect 4068 23749 4102 23783
rect 6561 23749 6595 23783
rect 6745 23749 6779 23783
rect 15884 23749 15918 23783
rect 17141 23749 17175 23783
rect 18429 23749 18463 23783
rect 19616 23749 19650 23783
rect 22937 23749 22971 23783
rect 31217 23749 31251 23783
rect 33057 23749 33091 23783
rect 35602 23749 35636 23783
rect 2329 23681 2363 23715
rect 3801 23681 3835 23715
rect 7389 23681 7423 23715
rect 7645 23681 7679 23715
rect 9965 23681 9999 23715
rect 10149 23681 10183 23715
rect 10241 23681 10275 23715
rect 10333 23681 10367 23715
rect 11897 23681 11931 23715
rect 12045 23681 12079 23715
rect 12173 23681 12207 23715
rect 12265 23681 12299 23715
rect 12362 23681 12396 23715
rect 13369 23681 13403 23715
rect 13553 23681 13587 23715
rect 13645 23681 13679 23715
rect 13737 23681 13771 23715
rect 17417 23681 17451 23715
rect 17509 23681 17543 23715
rect 17601 23681 17635 23715
rect 17785 23681 17819 23715
rect 18245 23681 18279 23715
rect 22385 23681 22419 23715
rect 23121 23681 23155 23715
rect 23765 23681 23799 23715
rect 23949 23681 23983 23715
rect 24041 23681 24075 23715
rect 24133 23681 24167 23715
rect 25237 23681 25271 23715
rect 25400 23681 25434 23715
rect 25500 23681 25534 23715
rect 25625 23681 25659 23715
rect 29561 23681 29595 23715
rect 29837 23681 29871 23715
rect 31401 23681 31435 23715
rect 32413 23681 32447 23715
rect 32597 23681 32631 23715
rect 32689 23681 32723 23715
rect 32781 23681 32815 23715
rect 34630 23681 34664 23715
rect 34897 23681 34931 23715
rect 35357 23681 35391 23715
rect 2605 23613 2639 23647
rect 16129 23613 16163 23647
rect 19349 23613 19383 23647
rect 23305 23613 23339 23647
rect 5181 23545 5215 23579
rect 14013 23545 14047 23579
rect 3157 23477 3191 23511
rect 6929 23477 6963 23511
rect 10517 23477 10551 23511
rect 12541 23477 12575 23511
rect 21189 23477 21223 23511
rect 24409 23477 24443 23511
rect 25881 23477 25915 23511
rect 31585 23477 31619 23511
rect 33517 23477 33551 23511
rect 5641 23273 5675 23307
rect 6377 23273 6411 23307
rect 11529 23273 11563 23307
rect 19349 23273 19383 23307
rect 21097 23273 21131 23307
rect 21925 23273 21959 23307
rect 25237 23273 25271 23307
rect 28917 23273 28951 23307
rect 29929 23273 29963 23307
rect 33701 23273 33735 23307
rect 9045 23205 9079 23239
rect 23305 23205 23339 23239
rect 32873 23205 32907 23239
rect 4261 23137 4295 23171
rect 9689 23137 9723 23171
rect 13001 23137 13035 23171
rect 15485 23137 15519 23171
rect 20269 23137 20303 23171
rect 25697 23137 25731 23171
rect 26985 23137 27019 23171
rect 31769 23137 31803 23171
rect 2145 23069 2179 23103
rect 2329 23069 2363 23103
rect 2421 23069 2455 23103
rect 2513 23069 2547 23103
rect 6653 23069 6687 23103
rect 6745 23069 6779 23103
rect 6837 23069 6871 23103
rect 7021 23069 7055 23103
rect 7481 23069 7515 23103
rect 7665 23069 7699 23103
rect 7757 23069 7791 23103
rect 7849 23069 7883 23103
rect 8953 23069 8987 23103
rect 9137 23069 9171 23103
rect 10609 23069 10643 23103
rect 10977 23069 11011 23103
rect 12725 23069 12759 23103
rect 15218 23069 15252 23103
rect 17049 23069 17083 23103
rect 17233 23069 17267 23103
rect 17325 23069 17359 23103
rect 17417 23069 17451 23103
rect 18521 23069 18555 23103
rect 20729 23069 20763 23103
rect 20913 23069 20947 23103
rect 21557 23069 21591 23103
rect 21741 23069 21775 23103
rect 24869 23069 24903 23103
rect 27241 23069 27275 23103
rect 28825 23069 28859 23103
rect 29009 23069 29043 23103
rect 29561 23069 29595 23103
rect 29745 23069 29779 23103
rect 32229 23069 32263 23103
rect 32408 23069 32442 23103
rect 32508 23066 32542 23100
rect 32597 23069 32631 23103
rect 33333 23069 33367 23103
rect 2789 23001 2823 23035
rect 4506 23001 4540 23035
rect 10701 23001 10735 23035
rect 10793 23001 10827 23035
rect 11621 23001 11655 23035
rect 18153 23001 18187 23035
rect 18337 23001 18371 23035
rect 22661 23001 22695 23035
rect 23489 23001 23523 23035
rect 25053 23001 25087 23035
rect 31502 23001 31536 23035
rect 33517 23001 33551 23035
rect 8125 22933 8159 22967
rect 10425 22933 10459 22967
rect 14105 22933 14139 22967
rect 17693 22933 17727 22967
rect 22753 22933 22787 22967
rect 28365 22933 28399 22967
rect 30389 22933 30423 22967
rect 2513 22729 2547 22763
rect 4537 22729 4571 22763
rect 5457 22729 5491 22763
rect 13553 22729 13587 22763
rect 18153 22729 18187 22763
rect 29377 22729 29411 22763
rect 31493 22729 31527 22763
rect 12173 22661 12207 22695
rect 13185 22661 13219 22695
rect 13369 22661 13403 22695
rect 19266 22661 19300 22695
rect 22017 22661 22051 22695
rect 30757 22661 30791 22695
rect 32505 22661 32539 22695
rect 2145 22593 2179 22627
rect 2329 22593 2363 22627
rect 3157 22593 3191 22627
rect 3413 22593 3447 22627
rect 5641 22593 5675 22627
rect 7941 22593 7975 22627
rect 8208 22593 8242 22627
rect 10701 22593 10735 22627
rect 11897 22593 11931 22627
rect 11990 22593 12024 22627
rect 12265 22593 12299 22627
rect 12362 22593 12396 22627
rect 14197 22593 14231 22627
rect 17601 22593 17635 22627
rect 24317 22593 24351 22627
rect 24410 22593 24444 22627
rect 24593 22593 24627 22627
rect 24685 22593 24719 22627
rect 24823 22593 24857 22627
rect 30573 22593 30607 22627
rect 32321 22593 32355 22627
rect 37289 22593 37323 22627
rect 37556 22593 37590 22627
rect 5825 22525 5859 22559
rect 7205 22525 7239 22559
rect 7481 22525 7515 22559
rect 10977 22525 11011 22559
rect 19533 22525 19567 22559
rect 23305 22525 23339 22559
rect 9321 22457 9355 22491
rect 12541 22457 12575 22491
rect 21281 22457 21315 22491
rect 67649 22457 67683 22491
rect 20637 22389 20671 22423
rect 23075 22389 23109 22423
rect 23765 22389 23799 22423
rect 24961 22389 24995 22423
rect 30941 22389 30975 22423
rect 32137 22389 32171 22423
rect 32965 22389 32999 22423
rect 38669 22389 38703 22423
rect 2237 22185 2271 22219
rect 17785 22185 17819 22219
rect 19717 22185 19751 22219
rect 27629 22185 27663 22219
rect 9505 22117 9539 22151
rect 12265 22117 12299 22151
rect 4997 22049 5031 22083
rect 6837 22049 6871 22083
rect 11161 22049 11195 22083
rect 14933 22049 14967 22083
rect 22753 22049 22787 22083
rect 25605 22049 25639 22083
rect 34069 22049 34103 22083
rect 1593 21981 1627 22015
rect 2605 21981 2639 22015
rect 7021 21981 7055 22015
rect 7665 21981 7699 22015
rect 7849 21981 7883 22015
rect 10885 21981 10919 22015
rect 11621 21981 11655 22015
rect 11714 21981 11748 22015
rect 11897 21981 11931 22015
rect 12127 21981 12161 22015
rect 13277 21981 13311 22015
rect 13553 21981 13587 22015
rect 14657 21981 14691 22015
rect 15945 21981 15979 22015
rect 16038 21981 16072 22015
rect 16310 21981 16344 22015
rect 16429 21981 16463 22015
rect 19625 21981 19659 22015
rect 20269 21981 20303 22015
rect 20637 21981 20671 22015
rect 22109 21981 22143 22015
rect 22293 21981 22327 22015
rect 22385 21981 22419 22015
rect 22477 21981 22511 22015
rect 23397 21981 23431 22015
rect 24409 21981 24443 22015
rect 24557 21981 24591 22015
rect 24777 21981 24811 22015
rect 24915 21981 24949 22015
rect 25861 21981 25895 22015
rect 28181 21981 28215 22015
rect 28365 21981 28399 22015
rect 28457 21981 28491 22015
rect 28595 21981 28629 22015
rect 30941 21981 30975 22015
rect 31861 21981 31895 22015
rect 32045 21981 32079 22015
rect 32137 21981 32171 22015
rect 32229 21981 32263 22015
rect 32965 21981 32999 22015
rect 33149 21981 33183 22015
rect 33241 21981 33275 22015
rect 33333 21981 33367 22015
rect 36277 21981 36311 22015
rect 1777 21913 1811 21947
rect 2421 21913 2455 21947
rect 5242 21913 5276 21947
rect 7205 21913 7239 21947
rect 9689 21913 9723 21947
rect 11989 21913 12023 21947
rect 16221 21913 16255 21947
rect 20453 21913 20487 21947
rect 20545 21913 20579 21947
rect 24685 21913 24719 21947
rect 28825 21913 28859 21947
rect 30674 21913 30708 21947
rect 33609 21913 33643 21947
rect 36010 21913 36044 21947
rect 1409 21845 1443 21879
rect 3065 21845 3099 21879
rect 6377 21845 6411 21879
rect 7665 21845 7699 21879
rect 16589 21845 16623 21879
rect 18613 21845 18647 21879
rect 20821 21845 20855 21879
rect 21373 21845 21407 21879
rect 23305 21845 23339 21879
rect 25053 21845 25087 21879
rect 26985 21845 27019 21879
rect 29561 21845 29595 21879
rect 32505 21845 32539 21879
rect 34897 21845 34931 21879
rect 2237 21641 2271 21675
rect 4077 21641 4111 21675
rect 10609 21641 10643 21675
rect 13737 21641 13771 21675
rect 16681 21641 16715 21675
rect 20913 21641 20947 21675
rect 28273 21641 28307 21675
rect 30665 21641 30699 21675
rect 32689 21641 32723 21675
rect 33517 21641 33551 21675
rect 36645 21641 36679 21675
rect 6377 21573 6411 21607
rect 9496 21573 9530 21607
rect 13369 21573 13403 21607
rect 14565 21573 14599 21607
rect 15485 21573 15519 21607
rect 19625 21573 19659 21607
rect 19717 21573 19751 21607
rect 20637 21573 20671 21607
rect 23765 21573 23799 21607
rect 28089 21573 28123 21607
rect 32321 21573 32355 21607
rect 32505 21573 32539 21607
rect 34630 21573 34664 21607
rect 35541 21573 35575 21607
rect 1593 21505 1627 21539
rect 1777 21505 1811 21539
rect 1869 21505 1903 21539
rect 1961 21505 1995 21539
rect 6561 21505 6595 21539
rect 13185 21505 13219 21539
rect 13461 21505 13495 21539
rect 13553 21505 13587 21539
rect 14381 21505 14415 21539
rect 15209 21505 15243 21539
rect 15357 21505 15391 21539
rect 15577 21505 15611 21539
rect 15715 21505 15749 21539
rect 17794 21505 17828 21539
rect 18797 21505 18831 21539
rect 19533 21505 19567 21539
rect 19901 21505 19935 21539
rect 20361 21505 20395 21539
rect 20545 21505 20579 21539
rect 20729 21505 20763 21539
rect 22937 21505 22971 21539
rect 23397 21505 23431 21539
rect 23581 21505 23615 21539
rect 25191 21505 25225 21539
rect 25329 21505 25363 21539
rect 25421 21505 25455 21539
rect 25604 21505 25638 21539
rect 25697 21505 25731 21539
rect 27905 21505 27939 21539
rect 29561 21505 29595 21539
rect 30205 21505 30239 21539
rect 30941 21505 30975 21539
rect 31033 21505 31067 21539
rect 31125 21505 31159 21539
rect 31309 21505 31343 21539
rect 36001 21505 36035 21539
rect 36185 21505 36219 21539
rect 36280 21505 36314 21539
rect 36415 21505 36449 21539
rect 37473 21505 37507 21539
rect 37740 21505 37774 21539
rect 2697 21437 2731 21471
rect 2973 21437 3007 21471
rect 9229 21437 9263 21471
rect 18061 21437 18095 21471
rect 22661 21437 22695 21471
rect 34897 21437 34931 21471
rect 6745 21369 6779 21403
rect 18613 21369 18647 21403
rect 5825 21301 5859 21335
rect 14749 21301 14783 21335
rect 15853 21301 15887 21335
rect 19349 21301 19383 21335
rect 25053 21301 25087 21335
rect 38853 21301 38887 21335
rect 67649 21301 67683 21335
rect 5181 21097 5215 21131
rect 15853 21097 15887 21131
rect 22753 21097 22787 21131
rect 34069 21097 34103 21131
rect 35449 21097 35483 21131
rect 37841 21097 37875 21131
rect 8125 21029 8159 21063
rect 24777 21029 24811 21063
rect 26341 21029 26375 21063
rect 6745 20961 6779 20995
rect 14657 20961 14691 20995
rect 35909 20961 35943 20995
rect 2053 20893 2087 20927
rect 2881 20893 2915 20927
rect 3801 20893 3835 20927
rect 9137 20893 9171 20927
rect 9321 20893 9355 20927
rect 10241 20893 10275 20927
rect 11069 20893 11103 20927
rect 11253 20893 11287 20927
rect 11345 20893 11379 20927
rect 11437 20893 11471 20927
rect 12173 20893 12207 20927
rect 13001 20893 13035 20927
rect 13277 20893 13311 20927
rect 13369 20893 13403 20927
rect 15209 20893 15243 20927
rect 15393 20893 15427 20927
rect 15485 20893 15519 20927
rect 15577 20893 15611 20927
rect 16313 20893 16347 20927
rect 16497 20893 16531 20927
rect 16589 20893 16623 20927
rect 16681 20893 16715 20927
rect 17417 20893 17451 20927
rect 18153 20893 18187 20927
rect 19717 20893 19751 20927
rect 25237 20893 25271 20927
rect 25421 20893 25455 20927
rect 25513 20893 25547 20927
rect 25605 20893 25639 20927
rect 27721 20893 27755 20927
rect 31769 20893 31803 20927
rect 32597 20893 32631 20927
rect 32781 20893 32815 20927
rect 32873 20893 32907 20927
rect 32965 20893 32999 20927
rect 35265 20893 35299 20927
rect 36185 20893 36219 20927
rect 37197 20893 37231 20927
rect 37381 20893 37415 20927
rect 37473 20893 37507 20927
rect 37565 20893 37599 20927
rect 1869 20825 1903 20859
rect 4046 20825 4080 20859
rect 7012 20825 7046 20859
rect 10425 20825 10459 20859
rect 10609 20825 10643 20859
rect 13185 20825 13219 20859
rect 16957 20825 16991 20859
rect 20545 20825 20579 20859
rect 25881 20825 25915 20859
rect 27454 20825 27488 20859
rect 31953 20825 31987 20859
rect 32137 20825 32171 20859
rect 35081 20825 35115 20859
rect 2237 20757 2271 20791
rect 2697 20757 2731 20791
rect 8953 20757 8987 20791
rect 11713 20757 11747 20791
rect 13553 20757 13587 20791
rect 18613 20757 18647 20791
rect 19901 20757 19935 20791
rect 21833 20757 21867 20791
rect 30665 20757 30699 20791
rect 31309 20757 31343 20791
rect 33241 20757 33275 20791
rect 2697 20553 2731 20587
rect 3801 20553 3835 20587
rect 7757 20553 7791 20587
rect 9965 20553 9999 20587
rect 14197 20553 14231 20587
rect 17049 20553 17083 20587
rect 19993 20553 20027 20587
rect 21925 20553 21959 20587
rect 26065 20553 26099 20587
rect 33149 20553 33183 20587
rect 36277 20553 36311 20587
rect 7205 20485 7239 20519
rect 9137 20485 9171 20519
rect 9321 20485 9355 20519
rect 13062 20485 13096 20519
rect 22744 20485 22778 20519
rect 25237 20485 25271 20519
rect 26241 20485 26275 20519
rect 31493 20485 31527 20519
rect 2053 20417 2087 20451
rect 2237 20417 2271 20451
rect 2329 20417 2363 20451
rect 2467 20417 2501 20451
rect 3157 20417 3191 20451
rect 3341 20417 3375 20451
rect 3433 20417 3467 20451
rect 3571 20417 3605 20451
rect 7021 20417 7055 20451
rect 7987 20417 8021 20451
rect 8125 20417 8159 20451
rect 8217 20417 8251 20451
rect 8401 20417 8435 20451
rect 16681 20417 16715 20451
rect 16865 20417 16899 20451
rect 17693 20417 17727 20451
rect 17960 20417 17994 20451
rect 21005 20417 21039 20451
rect 22477 20417 22511 20451
rect 25099 20417 25133 20451
rect 25329 20417 25363 20451
rect 25512 20417 25546 20451
rect 25605 20417 25639 20451
rect 26433 20417 26467 20451
rect 27997 20417 28031 20451
rect 28181 20417 28215 20451
rect 29938 20417 29972 20451
rect 30205 20417 30239 20451
rect 34262 20417 34296 20451
rect 34529 20417 34563 20451
rect 34989 20417 35023 20451
rect 12817 20349 12851 20383
rect 21281 20349 21315 20383
rect 19073 20281 19107 20315
rect 24961 20281 24995 20315
rect 28825 20281 28859 20315
rect 1593 20213 1627 20247
rect 4353 20213 4387 20247
rect 5733 20213 5767 20247
rect 6837 20213 6871 20247
rect 9505 20213 9539 20247
rect 11529 20213 11563 20247
rect 23857 20213 23891 20247
rect 28365 20213 28399 20247
rect 32505 20213 32539 20247
rect 37381 20213 37415 20247
rect 9045 20009 9079 20043
rect 13001 20009 13035 20043
rect 18705 20009 18739 20043
rect 21373 20009 21407 20043
rect 24961 20009 24995 20043
rect 27813 20009 27847 20043
rect 29009 20009 29043 20043
rect 34805 20009 34839 20043
rect 36461 20009 36495 20043
rect 17877 19941 17911 19975
rect 31125 19941 31159 19975
rect 35541 19941 35575 19975
rect 7573 19873 7607 19907
rect 11621 19873 11655 19907
rect 15761 19873 15795 19907
rect 20637 19873 20671 19907
rect 21833 19873 21867 19907
rect 37657 19873 37691 19907
rect 1593 19805 1627 19839
rect 2329 19805 2363 19839
rect 2513 19805 2547 19839
rect 2605 19805 2639 19839
rect 2697 19805 2731 19839
rect 3801 19805 3835 19839
rect 4905 19805 4939 19839
rect 5365 19805 5399 19839
rect 6469 19805 6503 19839
rect 6561 19805 6595 19839
rect 6653 19805 6687 19839
rect 6837 19805 6871 19839
rect 7297 19805 7331 19839
rect 9321 19805 9355 19839
rect 9413 19805 9447 19839
rect 9505 19805 9539 19839
rect 9689 19805 9723 19839
rect 10517 19805 10551 19839
rect 10701 19805 10735 19839
rect 10793 19805 10827 19839
rect 10885 19805 10919 19839
rect 14657 19805 14691 19839
rect 14841 19805 14875 19839
rect 14933 19805 14967 19839
rect 15025 19805 15059 19839
rect 22109 19805 22143 19839
rect 23305 19805 23339 19839
rect 23581 19805 23615 19839
rect 23673 19805 23707 19839
rect 24409 19805 24443 19839
rect 24685 19805 24719 19839
rect 24777 19805 24811 19839
rect 25881 19805 25915 19839
rect 25974 19805 26008 19839
rect 26346 19805 26380 19839
rect 28365 19805 28399 19839
rect 28549 19805 28583 19839
rect 28641 19805 28675 19839
rect 28733 19805 28767 19839
rect 30481 19805 30515 19839
rect 32505 19805 32539 19839
rect 36093 19805 36127 19839
rect 68109 19805 68143 19839
rect 11161 19737 11195 19771
rect 11866 19737 11900 19771
rect 14105 19737 14139 19771
rect 15301 19737 15335 19771
rect 16006 19737 16040 19771
rect 18061 19737 18095 19771
rect 20392 19737 20426 19771
rect 23489 19737 23523 19771
rect 24593 19737 24627 19771
rect 26157 19737 26191 19771
rect 26249 19737 26283 19771
rect 30297 19737 30331 19771
rect 32238 19737 32272 19771
rect 36277 19737 36311 19771
rect 37924 19737 37958 19771
rect 1777 19669 1811 19703
rect 2973 19669 3007 19703
rect 5549 19669 5583 19703
rect 6193 19669 6227 19703
rect 17141 19669 17175 19703
rect 19257 19669 19291 19703
rect 23857 19669 23891 19703
rect 26525 19669 26559 19703
rect 30665 19669 30699 19703
rect 39037 19669 39071 19703
rect 2145 19465 2179 19499
rect 2605 19465 2639 19499
rect 5825 19465 5859 19499
rect 13369 19465 13403 19499
rect 14565 19465 14599 19499
rect 18705 19465 18739 19499
rect 24593 19465 24627 19499
rect 25789 19465 25823 19499
rect 31217 19465 31251 19499
rect 35909 19465 35943 19499
rect 38117 19465 38151 19499
rect 1777 19397 1811 19431
rect 1961 19397 1995 19431
rect 3718 19397 3752 19431
rect 4712 19397 4746 19431
rect 6745 19397 6779 19431
rect 11713 19397 11747 19431
rect 14289 19397 14323 19431
rect 15577 19397 15611 19431
rect 20177 19397 20211 19431
rect 22937 19397 22971 19431
rect 24225 19397 24259 19431
rect 24317 19397 24351 19431
rect 37657 19397 37691 19431
rect 4445 19329 4479 19363
rect 8493 19329 8527 19363
rect 8953 19329 8987 19363
rect 9209 19329 9243 19363
rect 11529 19329 11563 19363
rect 12633 19329 12667 19363
rect 13921 19329 13955 19363
rect 14014 19329 14048 19363
rect 14197 19329 14231 19363
rect 14386 19329 14420 19363
rect 15393 19329 15427 19363
rect 17325 19329 17359 19363
rect 17581 19329 17615 19363
rect 19993 19329 20027 19363
rect 20913 19329 20947 19363
rect 21002 19329 21036 19363
rect 21097 19329 21131 19363
rect 21281 19329 21315 19363
rect 22063 19329 22097 19363
rect 22198 19329 22232 19363
rect 22293 19329 22327 19363
rect 22477 19329 22511 19363
rect 23121 19329 23155 19363
rect 23305 19329 23339 19363
rect 24041 19329 24075 19363
rect 24409 19329 24443 19363
rect 25927 19329 25961 19363
rect 26065 19329 26099 19363
rect 26157 19329 26191 19363
rect 26340 19329 26374 19363
rect 26433 19329 26467 19363
rect 29745 19329 29779 19363
rect 29929 19329 29963 19363
rect 30573 19329 30607 19363
rect 30757 19329 30791 19363
rect 30852 19329 30886 19363
rect 30941 19329 30975 19363
rect 34733 19329 34767 19363
rect 34989 19329 35023 19363
rect 36185 19329 36219 19363
rect 36274 19332 36308 19366
rect 36390 19329 36424 19363
rect 36553 19329 36587 19363
rect 37289 19329 37323 19363
rect 37473 19329 37507 19363
rect 38347 19329 38381 19363
rect 38485 19329 38519 19363
rect 38577 19329 38611 19363
rect 38761 19329 38795 19363
rect 3985 19261 4019 19295
rect 11897 19261 11931 19295
rect 15209 19261 15243 19295
rect 16865 19261 16899 19295
rect 19809 19261 19843 19295
rect 12817 19193 12851 19227
rect 20637 19193 20671 19227
rect 32229 19193 32263 19227
rect 10333 19125 10367 19159
rect 16037 19125 16071 19159
rect 19349 19125 19383 19159
rect 21833 19125 21867 19159
rect 30113 19125 30147 19159
rect 33609 19125 33643 19159
rect 6469 18921 6503 18955
rect 8953 18921 8987 18955
rect 17233 18921 17267 18955
rect 18705 18921 18739 18955
rect 20085 18921 20119 18955
rect 31585 18921 31619 18955
rect 34713 18921 34747 18955
rect 14105 18853 14139 18887
rect 19441 18853 19475 18887
rect 31033 18853 31067 18887
rect 2329 18785 2363 18819
rect 2605 18785 2639 18819
rect 7849 18785 7883 18819
rect 11253 18785 11287 18819
rect 15209 18785 15243 18819
rect 20913 18785 20947 18819
rect 29837 18785 29871 18819
rect 33793 18785 33827 18819
rect 6745 18717 6779 18751
rect 6837 18717 6871 18751
rect 6929 18717 6963 18751
rect 7113 18717 7147 18751
rect 7573 18717 7607 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 10425 18717 10459 18751
rect 10517 18717 10551 18751
rect 12357 18717 12391 18751
rect 12633 18717 12667 18751
rect 12725 18717 12759 18751
rect 15485 18717 15519 18751
rect 19257 18717 19291 18751
rect 20269 18717 20303 18751
rect 21180 18717 21214 18751
rect 23029 18717 23063 18751
rect 23305 18717 23339 18751
rect 24956 18717 24990 18751
rect 25053 18717 25087 18751
rect 25328 18717 25362 18751
rect 25421 18717 25455 18751
rect 26709 18717 26743 18751
rect 27537 18717 27571 18751
rect 29561 18717 29595 18751
rect 30849 18717 30883 18751
rect 32965 18717 32999 18751
rect 34943 18717 34977 18751
rect 35078 18717 35112 18751
rect 35178 18717 35212 18751
rect 35357 18717 35391 18751
rect 37298 18717 37332 18751
rect 37565 18717 37599 18751
rect 68109 18717 68143 18751
rect 12541 18649 12575 18683
rect 15945 18649 15979 18683
rect 25145 18649 25179 18683
rect 26893 18649 26927 18683
rect 27804 18649 27838 18683
rect 32698 18649 32732 18683
rect 33977 18649 34011 18683
rect 34161 18649 34195 18683
rect 3157 18581 3191 18615
rect 10793 18581 10827 18615
rect 12909 18581 12943 18615
rect 22293 18581 22327 18615
rect 24777 18581 24811 18615
rect 27077 18581 27111 18615
rect 28917 18581 28951 18615
rect 36185 18581 36219 18615
rect 38025 18581 38059 18615
rect 7297 18377 7331 18411
rect 10333 18377 10367 18411
rect 13185 18377 13219 18411
rect 15025 18377 15059 18411
rect 16129 18377 16163 18411
rect 19993 18377 20027 18411
rect 24317 18377 24351 18411
rect 27813 18377 27847 18411
rect 30757 18377 30791 18411
rect 34253 18377 34287 18411
rect 36461 18377 36495 18411
rect 2789 18309 2823 18343
rect 3862 18309 3896 18343
rect 7481 18309 7515 18343
rect 7665 18309 7699 18343
rect 10517 18309 10551 18343
rect 17233 18309 17267 18343
rect 18858 18309 18892 18343
rect 24041 18309 24075 18343
rect 25053 18309 25087 18343
rect 32229 18309 32263 18343
rect 32781 18309 32815 18343
rect 36093 18309 36127 18343
rect 2145 18241 2179 18275
rect 2329 18241 2363 18275
rect 2421 18241 2455 18275
rect 2513 18241 2547 18275
rect 6653 18241 6687 18275
rect 8125 18241 8159 18275
rect 10701 18241 10735 18275
rect 12357 18241 12391 18275
rect 12541 18241 12575 18275
rect 13093 18241 13127 18275
rect 13737 18241 13771 18275
rect 13830 18241 13864 18275
rect 14013 18241 14047 18275
rect 14105 18241 14139 18275
rect 14243 18241 14277 18275
rect 15485 18241 15519 18275
rect 15669 18241 15703 18275
rect 15761 18241 15795 18275
rect 15853 18241 15887 18275
rect 17049 18241 17083 18275
rect 18613 18241 18647 18275
rect 20453 18241 20487 18275
rect 23765 18241 23799 18275
rect 23949 18241 23983 18275
rect 24133 18241 24167 18275
rect 24777 18241 24811 18275
rect 24961 18241 24995 18275
rect 25145 18241 25179 18275
rect 27169 18241 27203 18275
rect 27353 18241 27387 18275
rect 27445 18241 27479 18275
rect 27583 18241 27617 18275
rect 28549 18241 28583 18275
rect 30119 18241 30153 18275
rect 30297 18241 30331 18275
rect 30389 18241 30423 18275
rect 30481 18241 30515 18275
rect 35081 18241 35115 18275
rect 36277 18241 36311 18275
rect 37749 18241 37783 18275
rect 38016 18241 38050 18275
rect 3617 18173 3651 18207
rect 6469 18173 6503 18207
rect 12449 18173 12483 18207
rect 20729 18173 20763 18207
rect 22477 18173 22511 18207
rect 22753 18173 22787 18207
rect 25789 18173 25823 18207
rect 28825 18173 28859 18207
rect 34805 18173 34839 18207
rect 25329 18105 25363 18139
rect 32965 18105 32999 18139
rect 4997 18037 5031 18071
rect 8309 18037 8343 18071
rect 9229 18037 9263 18071
rect 9873 18037 9907 18071
rect 14381 18037 14415 18071
rect 17417 18037 17451 18071
rect 18061 18037 18095 18071
rect 21925 18037 21959 18071
rect 31217 18037 31251 18071
rect 39129 18037 39163 18071
rect 1501 17833 1535 17867
rect 8953 17833 8987 17867
rect 11989 17833 12023 17867
rect 14933 17833 14967 17867
rect 15761 17833 15795 17867
rect 17693 17833 17727 17867
rect 21465 17833 21499 17867
rect 28825 17833 28859 17867
rect 34897 17833 34931 17867
rect 38209 17833 38243 17867
rect 21005 17765 21039 17799
rect 24501 17765 24535 17799
rect 35357 17765 35391 17799
rect 5365 17697 5399 17731
rect 9321 17697 9355 17731
rect 10609 17697 10643 17731
rect 22293 17697 22327 17731
rect 32229 17697 32263 17731
rect 36185 17697 36219 17731
rect 1961 17629 1995 17663
rect 2145 17629 2179 17663
rect 2237 17629 2271 17663
rect 2329 17629 2363 17663
rect 7205 17629 7239 17663
rect 7481 17629 7515 17663
rect 9137 17629 9171 17663
rect 9965 17629 9999 17663
rect 10876 17629 10910 17663
rect 12725 17629 12759 17663
rect 13001 17629 13035 17663
rect 14565 17629 14599 17663
rect 14749 17629 14783 17663
rect 15945 17629 15979 17663
rect 17049 17629 17083 17663
rect 17233 17629 17267 17663
rect 17325 17629 17359 17663
rect 17417 17629 17451 17663
rect 19809 17629 19843 17663
rect 20453 17629 20487 17663
rect 20637 17629 20671 17663
rect 20821 17629 20855 17663
rect 22017 17629 22051 17663
rect 25651 17629 25685 17663
rect 25881 17629 25915 17663
rect 26064 17629 26098 17663
rect 26157 17629 26191 17663
rect 26617 17629 26651 17663
rect 26801 17629 26835 17663
rect 29009 17629 29043 17663
rect 29745 17629 29779 17663
rect 29837 17629 29871 17663
rect 30113 17629 30147 17663
rect 32965 17629 32999 17663
rect 33701 17629 33735 17663
rect 33793 17629 33827 17663
rect 33885 17629 33919 17663
rect 34069 17629 34103 17663
rect 34713 17629 34747 17663
rect 35909 17629 35943 17663
rect 38485 17629 38519 17663
rect 38577 17629 38611 17663
rect 38669 17629 38703 17663
rect 38853 17629 38887 17663
rect 5610 17561 5644 17595
rect 16129 17561 16163 17595
rect 18705 17561 18739 17595
rect 19993 17561 20027 17595
rect 20729 17561 20763 17595
rect 23397 17561 23431 17595
rect 25789 17561 25823 17595
rect 29929 17561 29963 17595
rect 31984 17561 32018 17595
rect 33425 17561 33459 17595
rect 2605 17493 2639 17527
rect 6745 17493 6779 17527
rect 9781 17493 9815 17527
rect 23489 17493 23523 17527
rect 25053 17493 25087 17527
rect 25513 17493 25547 17527
rect 26985 17493 27019 17527
rect 27997 17493 28031 17527
rect 29561 17493 29595 17527
rect 30849 17493 30883 17527
rect 37657 17493 37691 17527
rect 2329 17289 2363 17323
rect 2789 17289 2823 17323
rect 6837 17289 6871 17323
rect 14565 17289 14599 17323
rect 16037 17289 16071 17323
rect 19165 17289 19199 17323
rect 26065 17289 26099 17323
rect 29653 17289 29687 17323
rect 32413 17289 32447 17323
rect 33241 17289 33275 17323
rect 38853 17289 38887 17323
rect 3862 17221 3896 17255
rect 9750 17221 9784 17255
rect 15209 17221 15243 17255
rect 15393 17221 15427 17255
rect 16865 17221 16899 17255
rect 17049 17221 17083 17255
rect 21005 17221 21039 17255
rect 29929 17221 29963 17255
rect 33057 17221 33091 17255
rect 1961 17153 1995 17187
rect 2145 17153 2179 17187
rect 2973 17153 3007 17187
rect 3157 17153 3191 17187
rect 3617 17153 3651 17187
rect 7297 17153 7331 17187
rect 7481 17153 7515 17187
rect 7573 17153 7607 17187
rect 7711 17153 7745 17187
rect 9505 17153 9539 17187
rect 13185 17153 13219 17187
rect 13441 17153 13475 17187
rect 15853 17153 15887 17187
rect 17785 17153 17819 17187
rect 18052 17153 18086 17187
rect 19993 17153 20027 17187
rect 20729 17153 20763 17187
rect 20913 17153 20947 17187
rect 21097 17153 21131 17187
rect 22201 17153 22235 17187
rect 25881 17153 25915 17187
rect 28374 17153 28408 17187
rect 28641 17153 28675 17187
rect 29837 17153 29871 17187
rect 30021 17153 30055 17187
rect 30205 17153 30239 17187
rect 32229 17153 32263 17187
rect 32404 17153 32438 17187
rect 32873 17153 32907 17187
rect 34345 17153 34379 17187
rect 34805 17153 34839 17187
rect 35081 17153 35115 17187
rect 36369 17153 36403 17187
rect 36461 17153 36495 17187
rect 36553 17153 36587 17187
rect 36737 17153 36771 17187
rect 38485 17153 38519 17187
rect 38669 17153 38703 17187
rect 24961 17085 24995 17119
rect 25237 17085 25271 17119
rect 25697 17085 25731 17119
rect 27261 17017 27295 17051
rect 37289 17017 37323 17051
rect 67649 17017 67683 17051
rect 4997 16949 5031 16983
rect 7941 16949 7975 16983
rect 8401 16949 8435 16983
rect 10885 16949 10919 16983
rect 15025 16949 15059 16983
rect 17233 16949 17267 16983
rect 20177 16949 20211 16983
rect 21281 16949 21315 16983
rect 23489 16949 23523 16983
rect 29193 16949 29227 16983
rect 31493 16949 31527 16983
rect 34161 16949 34195 16983
rect 36093 16949 36127 16983
rect 12817 16745 12851 16779
rect 15485 16745 15519 16779
rect 16635 16745 16669 16779
rect 17969 16745 18003 16779
rect 21741 16745 21775 16779
rect 27721 16745 27755 16779
rect 32689 16745 32723 16779
rect 35081 16745 35115 16779
rect 3065 16677 3099 16711
rect 7665 16677 7699 16711
rect 14381 16677 14415 16711
rect 18705 16677 18739 16711
rect 2329 16609 2363 16643
rect 2605 16609 2639 16643
rect 9505 16609 9539 16643
rect 10977 16609 11011 16643
rect 16865 16609 16899 16643
rect 19809 16609 19843 16643
rect 23121 16609 23155 16643
rect 25789 16609 25823 16643
rect 31033 16609 31067 16643
rect 35909 16609 35943 16643
rect 3801 16541 3835 16575
rect 3985 16541 4019 16575
rect 8125 16541 8159 16575
rect 9781 16541 9815 16575
rect 10333 16541 10367 16575
rect 13093 16541 13127 16575
rect 13185 16541 13219 16575
rect 13277 16541 13311 16575
rect 13461 16541 13495 16575
rect 17325 16541 17359 16575
rect 17509 16541 17543 16575
rect 17601 16541 17635 16575
rect 17693 16541 17727 16575
rect 19533 16541 19567 16575
rect 20821 16541 20855 16575
rect 21920 16541 21954 16575
rect 22292 16541 22326 16575
rect 22385 16541 22419 16575
rect 22845 16541 22879 16575
rect 26249 16541 26283 16575
rect 26433 16541 26467 16575
rect 29745 16541 29779 16575
rect 29929 16541 29963 16575
rect 30113 16541 30147 16575
rect 30757 16541 30791 16575
rect 32321 16541 32355 16575
rect 32505 16541 32539 16575
rect 34713 16541 34747 16575
rect 36176 16541 36210 16575
rect 39129 16541 39163 16575
rect 6929 16473 6963 16507
rect 7481 16473 7515 16507
rect 11222 16473 11256 16507
rect 22017 16473 22051 16507
rect 22109 16473 22143 16507
rect 25544 16473 25578 16507
rect 29009 16473 29043 16507
rect 29837 16473 29871 16507
rect 33149 16473 33183 16507
rect 34897 16473 34931 16507
rect 38862 16473 38896 16507
rect 4169 16405 4203 16439
rect 8309 16405 8343 16439
rect 12357 16405 12391 16439
rect 21005 16405 21039 16439
rect 24409 16405 24443 16439
rect 26433 16405 26467 16439
rect 29561 16405 29595 16439
rect 33977 16405 34011 16439
rect 37289 16405 37323 16439
rect 37749 16405 37783 16439
rect 3249 16201 3283 16235
rect 9781 16201 9815 16235
rect 10977 16201 11011 16235
rect 11897 16201 11931 16235
rect 18429 16201 18463 16235
rect 21097 16201 21131 16235
rect 24225 16201 24259 16235
rect 27629 16201 27663 16235
rect 28089 16201 28123 16235
rect 36553 16201 36587 16235
rect 3801 16133 3835 16167
rect 12449 16133 12483 16167
rect 15485 16133 15519 16167
rect 15853 16133 15887 16167
rect 19717 16133 19751 16167
rect 19809 16133 19843 16167
rect 22109 16133 22143 16167
rect 25973 16133 26007 16167
rect 31033 16133 31067 16167
rect 33456 16133 33490 16167
rect 34161 16133 34195 16167
rect 37289 16133 37323 16167
rect 37657 16133 37691 16167
rect 2605 16065 2639 16099
rect 2789 16065 2823 16099
rect 2881 16065 2915 16099
rect 2973 16065 3007 16099
rect 4537 16065 4571 16099
rect 4716 16065 4750 16099
rect 4816 16065 4850 16099
rect 4951 16065 4985 16099
rect 6653 16065 6687 16099
rect 6837 16065 6871 16099
rect 7757 16065 7791 16099
rect 8024 16065 8058 16099
rect 10333 16065 10367 16099
rect 10517 16065 10551 16099
rect 10609 16065 10643 16099
rect 10701 16065 10735 16099
rect 12633 16065 12667 16099
rect 13553 16065 13587 16099
rect 13716 16065 13750 16099
rect 13832 16065 13866 16099
rect 13921 16065 13955 16099
rect 14657 16065 14691 16099
rect 15669 16065 15703 16099
rect 19625 16065 19659 16099
rect 19993 16065 20027 16099
rect 21189 16065 21223 16099
rect 21971 16065 22005 16099
rect 22201 16065 22235 16099
rect 22384 16065 22418 16099
rect 22477 16065 22511 16099
rect 23029 16065 23063 16099
rect 23581 16065 23615 16099
rect 25789 16065 25823 16099
rect 26985 16065 27019 16099
rect 27169 16065 27203 16099
rect 27264 16065 27298 16099
rect 27353 16065 27387 16099
rect 28365 16065 28399 16099
rect 28457 16065 28491 16099
rect 28549 16065 28583 16099
rect 28733 16065 28767 16099
rect 29929 16065 29963 16099
rect 30941 16065 30975 16099
rect 31125 16065 31159 16099
rect 31309 16065 31343 16099
rect 33701 16065 33735 16099
rect 34437 16065 34471 16099
rect 34529 16065 34563 16099
rect 34621 16065 34655 16099
rect 34805 16065 34839 16099
rect 35909 16065 35943 16099
rect 36093 16065 36127 16099
rect 36185 16065 36219 16099
rect 36277 16065 36311 16099
rect 37473 16065 37507 16099
rect 6469 15997 6503 16031
rect 14197 15997 14231 16031
rect 16681 15997 16715 16031
rect 16957 15997 16991 16031
rect 26157 15997 26191 16031
rect 30205 15997 30239 16031
rect 21833 15929 21867 15963
rect 5181 15861 5215 15895
rect 9137 15861 9171 15895
rect 18981 15861 19015 15895
rect 19441 15861 19475 15895
rect 20545 15861 20579 15895
rect 23673 15861 23707 15895
rect 25237 15861 25271 15895
rect 30757 15861 30791 15895
rect 32321 15861 32355 15895
rect 35357 15861 35391 15895
rect 67649 15861 67683 15895
rect 2973 15657 3007 15691
rect 4537 15657 4571 15691
rect 6377 15657 6411 15691
rect 7665 15657 7699 15691
rect 8309 15657 8343 15691
rect 10885 15657 10919 15691
rect 14197 15657 14231 15691
rect 15393 15657 15427 15691
rect 21465 15657 21499 15691
rect 22385 15657 22419 15691
rect 23765 15657 23799 15691
rect 26341 15657 26375 15691
rect 33793 15657 33827 15691
rect 9505 15589 9539 15623
rect 15485 15521 15519 15555
rect 27169 15521 27203 15555
rect 32965 15521 32999 15555
rect 38945 15521 38979 15555
rect 2329 15453 2363 15487
rect 2513 15453 2547 15487
rect 2605 15453 2639 15487
rect 2743 15453 2777 15487
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 4997 15453 5031 15487
rect 5264 15453 5298 15487
rect 7113 15453 7147 15487
rect 7389 15453 7423 15487
rect 7481 15453 7515 15487
rect 8953 15453 8987 15487
rect 9229 15453 9263 15487
rect 9321 15453 9355 15487
rect 15577 15453 15611 15487
rect 16957 15453 16991 15487
rect 17141 15453 17175 15487
rect 17236 15453 17270 15487
rect 17345 15453 17379 15487
rect 18613 15453 18647 15487
rect 19855 15453 19889 15487
rect 19996 15453 20030 15487
rect 20268 15453 20302 15487
rect 20361 15453 20395 15487
rect 22293 15453 22327 15487
rect 22385 15453 22419 15487
rect 23121 15453 23155 15487
rect 24409 15453 24443 15487
rect 26801 15453 26835 15487
rect 26985 15453 27019 15487
rect 27629 15453 27663 15487
rect 27813 15453 27847 15487
rect 27905 15453 27939 15487
rect 27997 15453 28031 15487
rect 30021 15453 30055 15487
rect 30113 15453 30147 15487
rect 30389 15453 30423 15487
rect 31217 15453 31251 15487
rect 33977 15453 34011 15487
rect 34161 15453 34195 15487
rect 35265 15453 35299 15487
rect 35449 15453 35483 15487
rect 35541 15453 35575 15487
rect 35633 15453 35667 15487
rect 1501 15385 1535 15419
rect 1685 15385 1719 15419
rect 1869 15385 1903 15419
rect 7297 15385 7331 15419
rect 8217 15385 8251 15419
rect 9137 15385 9171 15419
rect 12173 15385 12207 15419
rect 13461 15385 13495 15419
rect 16405 15385 16439 15419
rect 18061 15385 18095 15419
rect 20085 15385 20119 15419
rect 21557 15385 21591 15419
rect 22109 15385 22143 15419
rect 23305 15385 23339 15419
rect 30205 15385 30239 15419
rect 35909 15385 35943 15419
rect 38678 15385 38712 15419
rect 3893 15317 3927 15351
rect 12817 15317 12851 15351
rect 14657 15317 14691 15351
rect 15209 15317 15243 15351
rect 17601 15317 17635 15351
rect 19717 15317 19751 15351
rect 20821 15317 20855 15351
rect 22569 15317 22603 15351
rect 28273 15317 28307 15351
rect 28733 15317 28767 15351
rect 29837 15317 29871 15351
rect 34713 15317 34747 15351
rect 37565 15317 37599 15351
rect 7849 15113 7883 15147
rect 9873 15113 9907 15147
rect 11713 15113 11747 15147
rect 19257 15113 19291 15147
rect 19901 15113 19935 15147
rect 29561 15113 29595 15147
rect 30389 15113 30423 15147
rect 36185 15113 36219 15147
rect 39681 15113 39715 15147
rect 4905 15045 4939 15079
rect 6837 15045 6871 15079
rect 8033 15045 8067 15079
rect 9045 15045 9079 15079
rect 12541 15045 12575 15079
rect 14197 15045 14231 15079
rect 18122 15045 18156 15079
rect 21281 15045 21315 15079
rect 21833 15045 21867 15079
rect 25912 15045 25946 15079
rect 26985 15045 27019 15079
rect 28426 15045 28460 15079
rect 31125 15045 31159 15079
rect 33517 15045 33551 15079
rect 33977 15045 34011 15079
rect 2421 14977 2455 15011
rect 3709 14977 3743 15011
rect 3893 14977 3927 15011
rect 3985 14977 4019 15011
rect 4077 14977 4111 15011
rect 6653 14977 6687 15011
rect 6929 14977 6963 15011
rect 7021 14977 7055 15011
rect 8217 14977 8251 15011
rect 8677 14977 8711 15011
rect 8861 14977 8895 15011
rect 9505 14977 9539 15011
rect 9689 14977 9723 15011
rect 10333 14977 10367 15011
rect 10496 14980 10530 15014
rect 10609 14977 10643 15011
rect 10721 14977 10755 15011
rect 11529 14977 11563 15011
rect 14749 14977 14783 15011
rect 15005 14977 15039 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 17877 14977 17911 15011
rect 20269 14977 20303 15011
rect 21005 14977 21039 15011
rect 22109 14977 22143 15011
rect 23020 14977 23054 15011
rect 27261 14977 27295 15011
rect 27353 14977 27387 15011
rect 27445 14977 27479 15011
rect 27629 14977 27663 15011
rect 31033 14977 31067 15011
rect 31217 14977 31251 15011
rect 31401 14977 31435 15011
rect 36369 14977 36403 15011
rect 36553 14977 36587 15011
rect 2697 14909 2731 14943
rect 20177 14909 20211 14943
rect 21189 14909 21223 14943
rect 21925 14909 21959 14943
rect 22753 14909 22787 14943
rect 26157 14909 26191 14943
rect 28181 14909 28215 14943
rect 7205 14841 7239 14875
rect 10977 14841 11011 14875
rect 16129 14841 16163 14875
rect 20821 14841 20855 14875
rect 24777 14841 24811 14875
rect 4353 14773 4387 14807
rect 20085 14773 20119 14807
rect 21281 14773 21315 14807
rect 21833 14773 21867 14807
rect 22293 14773 22327 14807
rect 24133 14773 24167 14807
rect 30849 14773 30883 14807
rect 35265 14773 35299 14807
rect 6009 14569 6043 14603
rect 7481 14569 7515 14603
rect 11069 14569 11103 14603
rect 14289 14569 14323 14603
rect 16589 14569 16623 14603
rect 17417 14569 17451 14603
rect 18613 14569 18647 14603
rect 21557 14569 21591 14603
rect 24685 14569 24719 14603
rect 26709 14569 26743 14603
rect 27537 14569 27571 14603
rect 37749 14569 37783 14603
rect 5365 14501 5399 14535
rect 7941 14501 7975 14535
rect 11529 14501 11563 14535
rect 13553 14501 13587 14535
rect 24869 14501 24903 14535
rect 9597 14433 9631 14467
rect 12909 14433 12943 14467
rect 16589 14433 16623 14467
rect 20913 14433 20947 14467
rect 24501 14433 24535 14467
rect 28825 14433 28859 14467
rect 30389 14433 30423 14467
rect 1869 14365 1903 14399
rect 2513 14365 2547 14399
rect 2697 14365 2731 14399
rect 3157 14365 3191 14399
rect 3985 14365 4019 14399
rect 4252 14365 4286 14399
rect 6193 14365 6227 14399
rect 6377 14365 6411 14399
rect 7113 14365 7147 14399
rect 7317 14365 7351 14399
rect 8953 14365 8987 14399
rect 9137 14365 9171 14399
rect 9873 14365 9907 14399
rect 14381 14365 14415 14399
rect 14473 14365 14507 14399
rect 14933 14365 14967 14399
rect 16681 14365 16715 14399
rect 17417 14365 17451 14399
rect 17601 14365 17635 14399
rect 24409 14365 24443 14399
rect 24685 14365 24719 14399
rect 28089 14365 28123 14399
rect 30113 14365 30147 14399
rect 31861 14365 31895 14399
rect 32045 14365 32079 14399
rect 32229 14365 32263 14399
rect 33149 14365 33183 14399
rect 33241 14365 33275 14399
rect 33517 14365 33551 14399
rect 37105 14365 37139 14399
rect 38873 14365 38907 14399
rect 39140 14365 39174 14399
rect 39865 14365 39899 14399
rect 40028 14365 40062 14399
rect 40141 14365 40175 14399
rect 40253 14365 40287 14399
rect 68109 14365 68143 14399
rect 8125 14297 8159 14331
rect 9045 14297 9079 14331
rect 12642 14297 12676 14331
rect 23121 14297 23155 14331
rect 23305 14297 23339 14331
rect 26341 14297 26375 14331
rect 26525 14297 26559 14331
rect 31953 14297 31987 14331
rect 33333 14297 33367 14331
rect 34897 14297 34931 14331
rect 35081 14297 35115 14331
rect 36838 14297 36872 14331
rect 40509 14297 40543 14331
rect 1685 14229 1719 14263
rect 2329 14229 2363 14263
rect 14105 14229 14139 14263
rect 15117 14229 15151 14263
rect 15853 14229 15887 14263
rect 16313 14229 16347 14263
rect 17785 14229 17819 14263
rect 19257 14229 19291 14263
rect 19901 14229 19935 14263
rect 22109 14229 22143 14263
rect 22937 14229 22971 14263
rect 28273 14229 28307 14263
rect 31677 14229 31711 14263
rect 32965 14229 32999 14263
rect 34713 14229 34747 14263
rect 35725 14229 35759 14263
rect 4077 14025 4111 14059
rect 5825 14025 5859 14059
rect 6561 14025 6595 14059
rect 7297 14025 7331 14059
rect 10885 14025 10919 14059
rect 12173 14025 12207 14059
rect 15577 14025 15611 14059
rect 19993 14025 20027 14059
rect 21281 14025 21315 14059
rect 32873 14025 32907 14059
rect 34069 14025 34103 14059
rect 35357 14025 35391 14059
rect 39313 14025 39347 14059
rect 40141 14025 40175 14059
rect 10517 13957 10551 13991
rect 11897 13957 11931 13991
rect 14657 13957 14691 13991
rect 18880 13957 18914 13991
rect 22937 13957 22971 13991
rect 24225 13957 24259 13991
rect 24961 13957 24995 13991
rect 26433 13957 26467 13991
rect 31309 13957 31343 13991
rect 33149 13957 33183 13991
rect 39957 13957 39991 13991
rect 1777 13889 1811 13923
rect 1961 13889 1995 13923
rect 2053 13889 2087 13923
rect 2145 13889 2179 13923
rect 2881 13889 2915 13923
rect 3065 13889 3099 13923
rect 3157 13889 3191 13923
rect 3249 13889 3283 13923
rect 5273 13889 5307 13923
rect 7113 13889 7147 13923
rect 7849 13889 7883 13923
rect 8033 13889 8067 13923
rect 8125 13889 8159 13923
rect 8217 13889 8251 13923
rect 8953 13889 8987 13923
rect 9229 13889 9263 13923
rect 10333 13889 10367 13923
rect 10609 13889 10643 13923
rect 10701 13889 10735 13923
rect 11621 13889 11655 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 13001 13889 13035 13923
rect 13921 13889 13955 13923
rect 14841 13889 14875 13923
rect 15393 13889 15427 13923
rect 20729 13889 20763 13923
rect 20913 13889 20947 13923
rect 21005 13889 21039 13923
rect 21143 13889 21177 13923
rect 22385 13889 22419 13923
rect 23167 13889 23201 13923
rect 23286 13889 23320 13923
rect 23397 13889 23431 13923
rect 23581 13889 23615 13923
rect 24409 13889 24443 13923
rect 26985 13889 27019 13923
rect 27169 13889 27203 13923
rect 28733 13889 28767 13923
rect 30573 13889 30607 13923
rect 31217 13889 31251 13923
rect 31401 13889 31435 13923
rect 31585 13889 31619 13923
rect 33057 13889 33091 13923
rect 33241 13889 33275 13923
rect 33425 13889 33459 13923
rect 34161 13889 34195 13923
rect 34713 13889 34747 13923
rect 34897 13889 34931 13923
rect 34989 13889 35023 13923
rect 35081 13889 35115 13923
rect 36185 13889 36219 13923
rect 36274 13892 36308 13926
rect 36369 13889 36403 13923
rect 36553 13889 36587 13923
rect 39773 13889 39807 13923
rect 2421 13821 2455 13855
rect 12909 13821 12943 13855
rect 17141 13821 17175 13855
rect 17601 13821 17635 13855
rect 18061 13821 18095 13855
rect 18613 13821 18647 13855
rect 28457 13821 28491 13855
rect 30297 13821 30331 13855
rect 35909 13821 35943 13855
rect 14105 13753 14139 13787
rect 17877 13753 17911 13787
rect 3525 13685 3559 13719
rect 8493 13685 8527 13719
rect 12633 13685 12667 13719
rect 12817 13685 12851 13719
rect 24041 13685 24075 13719
rect 27353 13685 27387 13719
rect 27905 13685 27939 13719
rect 31033 13685 31067 13719
rect 1961 13481 1995 13515
rect 8033 13481 8067 13515
rect 10885 13481 10919 13515
rect 17325 13481 17359 13515
rect 21373 13481 21407 13515
rect 22661 13481 22695 13515
rect 23213 13481 23247 13515
rect 28917 13481 28951 13515
rect 32873 13481 32907 13515
rect 34161 13481 34195 13515
rect 37565 13481 37599 13515
rect 6469 13413 6503 13447
rect 13461 13413 13495 13447
rect 14289 13413 14323 13447
rect 21833 13413 21867 13447
rect 32413 13413 32447 13447
rect 34713 13413 34747 13447
rect 36185 13413 36219 13447
rect 2421 13345 2455 13379
rect 5089 13345 5123 13379
rect 8953 13345 8987 13379
rect 11621 13345 11655 13379
rect 13553 13345 13587 13379
rect 14105 13345 14139 13379
rect 14565 13345 14599 13379
rect 15393 13345 15427 13379
rect 18705 13345 18739 13379
rect 26801 13345 26835 13379
rect 27537 13345 27571 13379
rect 31033 13345 31067 13379
rect 35633 13345 35667 13379
rect 38945 13345 38979 13379
rect 1593 13277 1627 13311
rect 2697 13277 2731 13311
rect 5345 13277 5379 13311
rect 7113 13277 7147 13311
rect 9229 13277 9263 13311
rect 10793 13277 10827 13311
rect 11897 13277 11931 13311
rect 18429 13277 18463 13311
rect 19625 13277 19659 13311
rect 20821 13277 20855 13311
rect 21189 13277 21223 13311
rect 21833 13277 21867 13311
rect 22017 13277 22051 13311
rect 23489 13277 23523 13311
rect 23581 13277 23615 13311
rect 23673 13277 23707 13311
rect 23857 13277 23891 13311
rect 29929 13277 29963 13311
rect 30297 13277 30331 13311
rect 30757 13277 30791 13311
rect 33057 13277 33091 13311
rect 33149 13277 33183 13311
rect 33425 13277 33459 13311
rect 35449 13277 35483 13311
rect 40141 13277 40175 13311
rect 40233 13277 40267 13311
rect 40325 13277 40359 13311
rect 40509 13277 40543 13311
rect 41153 13277 41187 13311
rect 68109 13277 68143 13311
rect 1777 13209 1811 13243
rect 7297 13209 7331 13243
rect 8217 13209 8251 13243
rect 8401 13209 8435 13243
rect 13093 13209 13127 13243
rect 15660 13209 15694 13243
rect 19441 13209 19475 13243
rect 21005 13209 21039 13243
rect 21097 13209 21131 13243
rect 24593 13209 24627 13243
rect 24777 13209 24811 13243
rect 26534 13209 26568 13243
rect 27782 13209 27816 13243
rect 30021 13209 30055 13243
rect 30113 13209 30147 13243
rect 33241 13209 33275 13243
rect 35265 13209 35299 13243
rect 38700 13209 38734 13243
rect 39865 13209 39899 13243
rect 40969 13209 41003 13243
rect 41337 13209 41371 13243
rect 6929 13141 6963 13175
rect 16773 13141 16807 13175
rect 19257 13141 19291 13175
rect 24961 13141 24995 13175
rect 25421 13141 25455 13175
rect 29745 13141 29779 13175
rect 3065 12937 3099 12971
rect 5733 12937 5767 12971
rect 8033 12937 8067 12971
rect 9873 12937 9907 12971
rect 10425 12937 10459 12971
rect 13277 12937 13311 12971
rect 15117 12937 15151 12971
rect 17141 12937 17175 12971
rect 17601 12937 17635 12971
rect 18981 12937 19015 12971
rect 21833 12937 21867 12971
rect 24317 12937 24351 12971
rect 25697 12937 25731 12971
rect 27629 12937 27663 12971
rect 10977 12869 11011 12903
rect 11989 12869 12023 12903
rect 12081 12869 12115 12903
rect 21281 12869 21315 12903
rect 24041 12869 24075 12903
rect 31401 12869 31435 12903
rect 32505 12869 32539 12903
rect 39037 12869 39071 12903
rect 1961 12801 1995 12835
rect 2697 12801 2731 12835
rect 2881 12801 2915 12835
rect 3801 12801 3835 12835
rect 4057 12801 4091 12835
rect 6745 12801 6779 12835
rect 6837 12801 6871 12835
rect 6929 12801 6963 12835
rect 7113 12801 7147 12835
rect 7849 12801 7883 12835
rect 8493 12801 8527 12835
rect 8760 12801 8794 12835
rect 11805 12801 11839 12835
rect 12173 12801 12207 12835
rect 13093 12801 13127 12835
rect 13277 12801 13311 12835
rect 14565 12801 14599 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 17877 12801 17911 12835
rect 17969 12801 18003 12835
rect 18061 12801 18095 12835
rect 18245 12801 18279 12835
rect 19533 12801 19567 12835
rect 23765 12801 23799 12835
rect 23949 12801 23983 12835
rect 24133 12801 24167 12835
rect 25053 12801 25087 12835
rect 25216 12801 25250 12835
rect 25329 12801 25363 12835
rect 25467 12801 25501 12835
rect 26985 12801 27019 12835
rect 27164 12801 27198 12835
rect 27261 12801 27295 12835
rect 27399 12801 27433 12835
rect 28457 12801 28491 12835
rect 29009 12801 29043 12835
rect 31217 12801 31251 12835
rect 31309 12801 31343 12835
rect 31585 12801 31619 12835
rect 32321 12801 32355 12835
rect 32413 12801 32447 12835
rect 32689 12801 32723 12835
rect 33977 12801 34011 12835
rect 35826 12801 35860 12835
rect 36093 12801 36127 12835
rect 39589 12801 39623 12835
rect 39865 12801 39899 12835
rect 14473 12733 14507 12767
rect 26433 12733 26467 12767
rect 29653 12733 29687 12767
rect 34253 12733 34287 12767
rect 5181 12665 5215 12699
rect 12357 12665 12391 12699
rect 15945 12665 15979 12699
rect 34713 12665 34747 12699
rect 38853 12665 38887 12699
rect 2145 12597 2179 12631
rect 6469 12597 6503 12631
rect 14197 12597 14231 12631
rect 14381 12597 14415 12631
rect 22661 12597 22695 12631
rect 29101 12597 29135 12631
rect 31033 12597 31067 12631
rect 32137 12597 32171 12631
rect 37473 12597 37507 12631
rect 10701 12393 10735 12427
rect 13001 12393 13035 12427
rect 15301 12393 15335 12427
rect 23673 12393 23707 12427
rect 26985 12393 27019 12427
rect 29837 12393 29871 12427
rect 30297 12393 30331 12427
rect 30941 12393 30975 12427
rect 39037 12393 39071 12427
rect 7941 12325 7975 12359
rect 10517 12325 10551 12359
rect 29009 12325 29043 12359
rect 32965 12325 32999 12359
rect 35725 12325 35759 12359
rect 3985 12257 4019 12291
rect 13093 12257 13127 12291
rect 20913 12257 20947 12291
rect 22845 12257 22879 12291
rect 25145 12257 25179 12291
rect 29929 12257 29963 12291
rect 32321 12257 32355 12291
rect 1685 12189 1719 12223
rect 1869 12189 1903 12223
rect 2605 12189 2639 12223
rect 2768 12189 2802 12223
rect 2881 12183 2915 12217
rect 2973 12189 3007 12223
rect 6561 12189 6595 12223
rect 6817 12189 6851 12223
rect 11161 12189 11195 12223
rect 11437 12189 11471 12223
rect 13185 12189 13219 12223
rect 14933 12189 14967 12223
rect 15117 12189 15151 12223
rect 17141 12189 17175 12223
rect 17969 12189 18003 12223
rect 18061 12189 18095 12223
rect 18153 12189 18187 12223
rect 18337 12189 18371 12223
rect 19809 12189 19843 12223
rect 19972 12183 20006 12217
rect 20104 12189 20138 12223
rect 20197 12189 20231 12223
rect 23029 12189 23063 12223
rect 23857 12189 23891 12223
rect 24869 12189 24903 12223
rect 26157 12189 26191 12223
rect 28457 12189 28491 12223
rect 28641 12189 28675 12223
rect 28733 12189 28767 12223
rect 28825 12189 28859 12223
rect 29837 12189 29871 12223
rect 30113 12189 30147 12223
rect 33747 12189 33781 12223
rect 33882 12189 33916 12223
rect 33977 12189 34011 12223
rect 34161 12189 34195 12223
rect 34713 12189 34747 12223
rect 34897 12189 34931 12223
rect 36838 12189 36872 12223
rect 37105 12189 37139 12223
rect 37565 12189 37599 12223
rect 40049 12189 40083 12223
rect 40233 12183 40267 12217
rect 40328 12183 40362 12217
rect 40417 12189 40451 12223
rect 41153 12189 41187 12223
rect 4230 12121 4264 12155
rect 10241 12121 10275 12155
rect 16896 12121 16930 12155
rect 17693 12121 17727 12155
rect 20453 12121 20487 12155
rect 21158 12121 21192 12155
rect 26341 12121 26375 12155
rect 32076 12121 32110 12155
rect 33517 12121 33551 12155
rect 40693 12121 40727 12155
rect 2053 12053 2087 12087
rect 3249 12053 3283 12087
rect 5365 12053 5399 12087
rect 12817 12053 12851 12087
rect 14473 12053 14507 12087
rect 15761 12053 15795 12087
rect 19349 12053 19383 12087
rect 22293 12053 22327 12087
rect 23213 12053 23247 12087
rect 26525 12053 26559 12087
rect 34805 12053 34839 12087
rect 3157 11849 3191 11883
rect 4077 11849 4111 11883
rect 7389 11849 7423 11883
rect 13093 11849 13127 11883
rect 14657 11849 14691 11883
rect 18061 11849 18095 11883
rect 19349 11849 19383 11883
rect 24593 11849 24627 11883
rect 25513 11849 25547 11883
rect 30021 11849 30055 11883
rect 30665 11849 30699 11883
rect 33793 11849 33827 11883
rect 35357 11849 35391 11883
rect 40233 11849 40267 11883
rect 3525 11781 3559 11815
rect 9321 11781 9355 11815
rect 10241 11781 10275 11815
rect 11989 11781 12023 11815
rect 12081 11781 12115 11815
rect 13921 11781 13955 11815
rect 17693 11781 17727 11815
rect 19165 11781 19199 11815
rect 22017 11781 22051 11815
rect 28733 11781 28767 11815
rect 32781 11781 32815 11815
rect 33609 11781 33643 11815
rect 39865 11781 39899 11815
rect 2053 11713 2087 11747
rect 2237 11713 2271 11747
rect 2329 11713 2363 11747
rect 2467 11713 2501 11747
rect 3341 11713 3375 11747
rect 9045 11713 9079 11747
rect 9229 11713 9263 11747
rect 9459 11713 9493 11747
rect 10057 11713 10091 11747
rect 10333 11713 10367 11747
rect 10425 11713 10459 11747
rect 11805 11713 11839 11747
rect 12173 11713 12207 11747
rect 12909 11713 12943 11747
rect 13737 11713 13771 11747
rect 17877 11713 17911 11747
rect 18981 11713 19015 11747
rect 19809 11713 19843 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 20223 11713 20257 11747
rect 21097 11713 21131 11747
rect 23305 11713 23339 11747
rect 23765 11713 23799 11747
rect 23949 11713 23983 11747
rect 24777 11713 24811 11747
rect 25053 11713 25087 11747
rect 25697 11713 25731 11747
rect 25973 11713 26007 11747
rect 26985 11713 27019 11747
rect 27148 11716 27182 11750
rect 27261 11713 27295 11747
rect 27399 11713 27433 11747
rect 28457 11713 28491 11747
rect 28641 11713 28675 11747
rect 28825 11713 28859 11747
rect 29561 11713 29595 11747
rect 29837 11713 29871 11747
rect 31401 11713 31435 11747
rect 32965 11713 32999 11747
rect 33425 11713 33459 11747
rect 34713 11713 34747 11747
rect 34876 11713 34910 11747
rect 34992 11713 35026 11747
rect 35081 11713 35115 11747
rect 35817 11713 35851 11747
rect 35980 11713 36014 11747
rect 36096 11713 36130 11747
rect 36231 11713 36265 11747
rect 38505 11713 38539 11747
rect 38761 11713 38795 11747
rect 40049 11713 40083 11747
rect 17141 11645 17175 11679
rect 23029 11645 23063 11679
rect 24869 11645 24903 11679
rect 25789 11645 25823 11679
rect 29653 11645 29687 11679
rect 31217 11645 31251 11679
rect 32597 11645 32631 11679
rect 2697 11577 2731 11611
rect 29009 11577 29043 11611
rect 37381 11577 37415 11611
rect 67649 11577 67683 11611
rect 6929 11509 6963 11543
rect 8401 11509 8435 11543
rect 9597 11509 9631 11543
rect 10609 11509 10643 11543
rect 12357 11509 12391 11543
rect 20453 11509 20487 11543
rect 20913 11509 20947 11543
rect 23857 11509 23891 11543
rect 25053 11509 25087 11543
rect 25973 11509 26007 11543
rect 27629 11509 27663 11543
rect 29837 11509 29871 11543
rect 31585 11509 31619 11543
rect 36461 11509 36495 11543
rect 6745 11305 6779 11339
rect 11529 11305 11563 11339
rect 12725 11305 12759 11339
rect 13277 11305 13311 11339
rect 16405 11305 16439 11339
rect 20085 11305 20119 11339
rect 22477 11305 22511 11339
rect 24409 11305 24443 11339
rect 28365 11305 28399 11339
rect 29009 11305 29043 11339
rect 29929 11305 29963 11339
rect 31125 11305 31159 11339
rect 32137 11305 32171 11339
rect 35265 11305 35299 11339
rect 16221 11237 16255 11271
rect 29653 11237 29687 11271
rect 35725 11237 35759 11271
rect 37565 11237 37599 11271
rect 2881 11169 2915 11203
rect 16497 11169 16531 11203
rect 17233 11169 17267 11203
rect 26985 11169 27019 11203
rect 38945 11169 38979 11203
rect 7941 11101 7975 11135
rect 8033 11101 8067 11135
rect 8125 11101 8159 11135
rect 8309 11101 8343 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 9689 11101 9723 11135
rect 10425 11101 10459 11135
rect 11069 11101 11103 11135
rect 11529 11101 11563 11135
rect 11713 11101 11747 11135
rect 14381 11101 14415 11135
rect 16589 11101 16623 11135
rect 17417 11101 17451 11135
rect 17601 11101 17635 11135
rect 18061 11101 18095 11135
rect 18245 11101 18279 11135
rect 18337 11101 18371 11135
rect 18475 11101 18509 11135
rect 19901 11101 19935 11135
rect 20637 11101 20671 11135
rect 21097 11101 21131 11135
rect 23489 11101 23523 11135
rect 23581 11101 23615 11135
rect 23673 11101 23707 11135
rect 23857 11101 23891 11135
rect 24961 11101 24995 11135
rect 25237 11101 25271 11135
rect 27252 11101 27286 11135
rect 29837 11101 29871 11135
rect 29929 11101 29963 11135
rect 31309 11101 31343 11135
rect 31401 11101 31435 11135
rect 31677 11101 31711 11135
rect 32321 11101 32355 11135
rect 32413 11101 32447 11135
rect 32689 11101 32723 11135
rect 33885 11101 33919 11135
rect 34161 11101 34195 11135
rect 34897 11101 34931 11135
rect 35081 11101 35115 11135
rect 37105 11101 37139 11135
rect 40141 11101 40175 11135
rect 40233 11101 40267 11135
rect 40325 11101 40359 11135
rect 40509 11101 40543 11135
rect 5457 11033 5491 11067
rect 13369 11033 13403 11067
rect 14648 11033 14682 11067
rect 18705 11033 18739 11067
rect 19717 11033 19751 11067
rect 21342 11033 21376 11067
rect 23213 11033 23247 11067
rect 30113 11033 30147 11067
rect 30573 11033 30607 11067
rect 31493 11033 31527 11067
rect 32505 11033 32539 11067
rect 36838 11033 36872 11067
rect 38700 11033 38734 11067
rect 39865 11033 39899 11067
rect 7665 10965 7699 10999
rect 9965 10965 9999 10999
rect 15761 10965 15795 10999
rect 2605 10761 2639 10795
rect 5825 10761 5859 10795
rect 6469 10761 6503 10795
rect 9321 10761 9355 10795
rect 13553 10761 13587 10795
rect 23305 10761 23339 10795
rect 30021 10761 30055 10795
rect 30573 10761 30607 10795
rect 31033 10761 31067 10795
rect 32137 10761 32171 10795
rect 39589 10761 39623 10795
rect 1409 10693 1443 10727
rect 1593 10693 1627 10727
rect 11713 10693 11747 10727
rect 31401 10693 31435 10727
rect 32505 10693 32539 10727
rect 35541 10693 35575 10727
rect 36277 10693 36311 10727
rect 39405 10693 39439 10727
rect 40141 10693 40175 10727
rect 3718 10625 3752 10659
rect 3985 10625 4019 10659
rect 4445 10625 4479 10659
rect 4712 10625 4746 10659
rect 6653 10625 6687 10659
rect 6837 10625 6871 10659
rect 7297 10625 7331 10659
rect 7564 10625 7598 10659
rect 9505 10625 9539 10659
rect 9689 10625 9723 10659
rect 11529 10625 11563 10659
rect 11805 10625 11839 10659
rect 11897 10625 11931 10659
rect 13369 10625 13403 10659
rect 14105 10625 14139 10659
rect 14289 10625 14323 10659
rect 14381 10625 14415 10659
rect 14657 10625 14691 10659
rect 17325 10625 17359 10659
rect 18153 10625 18187 10659
rect 18889 10625 18923 10659
rect 18981 10625 19015 10659
rect 19625 10625 19659 10659
rect 20545 10625 20579 10659
rect 21833 10625 21867 10659
rect 22017 10625 22051 10659
rect 22477 10625 22511 10659
rect 23765 10625 23799 10659
rect 24685 10625 24719 10659
rect 24961 10625 24995 10659
rect 27445 10625 27479 10659
rect 29561 10625 29595 10659
rect 29837 10625 29871 10659
rect 31217 10625 31251 10659
rect 31309 10625 31343 10659
rect 31585 10625 31619 10659
rect 32321 10625 32355 10659
rect 32413 10625 32447 10659
rect 32689 10625 32723 10659
rect 33333 10625 33367 10659
rect 34161 10625 34195 10659
rect 34437 10625 34471 10659
rect 39221 10625 39255 10659
rect 14473 10557 14507 10591
rect 17233 10557 17267 10591
rect 19441 10557 19475 10591
rect 20269 10557 20303 10591
rect 29653 10557 29687 10591
rect 33149 10557 33183 10591
rect 35725 10557 35759 10591
rect 12081 10489 12115 10523
rect 21925 10489 21959 10523
rect 27629 10489 27663 10523
rect 1777 10421 1811 10455
rect 8677 10421 8711 10455
rect 14841 10421 14875 10455
rect 16957 10421 16991 10455
rect 17141 10421 17175 10455
rect 18613 10421 18647 10455
rect 18797 10421 18831 10455
rect 19809 10421 19843 10455
rect 23949 10421 23983 10455
rect 26433 10421 26467 10455
rect 29837 10421 29871 10455
rect 33517 10421 33551 10455
rect 67649 10421 67683 10455
rect 3065 10217 3099 10251
rect 7481 10217 7515 10251
rect 11345 10217 11379 10251
rect 20637 10217 20671 10251
rect 22017 10217 22051 10251
rect 27537 10217 27571 10251
rect 29009 10217 29043 10251
rect 30113 10217 30147 10251
rect 35725 10217 35759 10251
rect 1961 10081 1995 10115
rect 9965 10081 9999 10115
rect 15577 10081 15611 10115
rect 17325 10081 17359 10115
rect 19257 10081 19291 10115
rect 23857 10081 23891 10115
rect 24685 10081 24719 10115
rect 27353 10081 27387 10115
rect 33241 10081 33275 10115
rect 1593 10013 1627 10047
rect 1777 10013 1811 10047
rect 2421 10013 2455 10047
rect 2605 10013 2639 10047
rect 2697 10013 2731 10047
rect 2789 10013 2823 10047
rect 3801 10013 3835 10047
rect 10221 10013 10255 10047
rect 13553 10013 13587 10047
rect 15301 10013 15335 10047
rect 15485 10013 15519 10047
rect 15669 10013 15703 10047
rect 15853 10013 15887 10047
rect 16957 10013 16991 10047
rect 17141 10013 17175 10047
rect 17233 10013 17267 10047
rect 17509 10013 17543 10047
rect 19513 10013 19547 10047
rect 21465 10013 21499 10047
rect 21833 10013 21867 10047
rect 23590 10013 23624 10047
rect 24961 10013 24995 10047
rect 25973 10013 26007 10047
rect 26249 10013 26283 10047
rect 27537 10013 27571 10047
rect 28457 10013 28491 10047
rect 28825 10013 28859 10047
rect 29561 10013 29595 10047
rect 29837 10013 29871 10047
rect 29929 10013 29963 10047
rect 31861 10013 31895 10047
rect 32137 10013 32171 10047
rect 32965 10013 32999 10047
rect 39129 10013 39163 10047
rect 40141 10013 40175 10047
rect 40233 10013 40267 10047
rect 40325 10013 40359 10047
rect 40509 10013 40543 10047
rect 13308 9945 13342 9979
rect 21649 9945 21683 9979
rect 21741 9945 21775 9979
rect 27261 9945 27295 9979
rect 28641 9945 28675 9979
rect 28733 9945 28767 9979
rect 29745 9945 29779 9979
rect 34713 9945 34747 9979
rect 34897 9945 34931 9979
rect 35633 9945 35667 9979
rect 38945 9945 38979 9979
rect 39313 9945 39347 9979
rect 12173 9877 12207 9911
rect 15117 9877 15151 9911
rect 17693 9877 17727 9911
rect 22477 9877 22511 9911
rect 27721 9877 27755 9911
rect 35081 9877 35115 9911
rect 39865 9877 39899 9911
rect 5273 9673 5307 9707
rect 13461 9673 13495 9707
rect 19349 9673 19383 9707
rect 21925 9673 21959 9707
rect 30297 9673 30331 9707
rect 37565 9673 37599 9707
rect 39773 9673 39807 9707
rect 2789 9605 2823 9639
rect 4138 9605 4172 9639
rect 8033 9605 8067 9639
rect 10333 9605 10367 9639
rect 10885 9605 10919 9639
rect 11713 9605 11747 9639
rect 21005 9605 21039 9639
rect 23489 9605 23523 9639
rect 23673 9605 23707 9639
rect 34897 9605 34931 9639
rect 36470 9605 36504 9639
rect 38700 9605 38734 9639
rect 2145 9537 2179 9571
rect 2308 9537 2342 9571
rect 2421 9537 2455 9571
rect 2513 9537 2547 9571
rect 3893 9537 3927 9571
rect 9137 9537 9171 9571
rect 9229 9537 9263 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 11529 9537 11563 9571
rect 11805 9537 11839 9571
rect 11897 9537 11931 9571
rect 12725 9537 12759 9571
rect 12909 9537 12943 9571
rect 13277 9537 13311 9571
rect 15016 9537 15050 9571
rect 18346 9537 18380 9571
rect 21189 9537 21223 9571
rect 21833 9537 21867 9571
rect 22017 9537 22051 9571
rect 22477 9537 22511 9571
rect 23305 9537 23339 9571
rect 25789 9537 25823 9571
rect 27629 9537 27663 9571
rect 27813 9537 27847 9571
rect 27905 9537 27939 9571
rect 27997 9537 28031 9571
rect 28733 9537 28767 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 33057 9537 33091 9571
rect 34253 9537 34287 9571
rect 34437 9537 34471 9571
rect 34529 9537 34563 9571
rect 34621 9537 34655 9571
rect 38945 9537 38979 9571
rect 3341 9469 3375 9503
rect 13001 9469 13035 9503
rect 13093 9469 13127 9503
rect 14749 9469 14783 9503
rect 18613 9469 18647 9503
rect 25513 9469 25547 9503
rect 31309 9469 31343 9503
rect 31585 9469 31619 9503
rect 32781 9469 32815 9503
rect 36737 9469 36771 9503
rect 32229 9401 32263 9435
rect 8861 9333 8895 9367
rect 12081 9333 12115 9367
rect 16129 9333 16163 9367
rect 17233 9333 17267 9367
rect 19993 9333 20027 9367
rect 20821 9333 20855 9367
rect 28273 9333 28307 9367
rect 35357 9333 35391 9367
rect 6837 9129 6871 9163
rect 10333 9129 10367 9163
rect 16313 9129 16347 9163
rect 24409 9129 24443 9163
rect 26157 9129 26191 9163
rect 27905 9129 27939 9163
rect 31401 9129 31435 9163
rect 34713 9129 34747 9163
rect 16865 9061 16899 9095
rect 33517 9061 33551 9095
rect 2329 8993 2363 9027
rect 2605 8993 2639 9027
rect 5457 8993 5491 9027
rect 8953 8993 8987 9027
rect 15393 8993 15427 9027
rect 15485 8993 15519 9027
rect 36645 8993 36679 9027
rect 3801 8925 3835 8959
rect 7573 8925 7607 8959
rect 7665 8925 7699 8959
rect 7757 8925 7791 8959
rect 7941 8925 7975 8959
rect 9209 8925 9243 8959
rect 15117 8925 15151 8959
rect 15301 8925 15335 8959
rect 15669 8925 15703 8959
rect 19441 8925 19475 8959
rect 19533 8925 19567 8959
rect 20177 8925 20211 8959
rect 20361 8925 20395 8959
rect 20453 8925 20487 8959
rect 20545 8925 20579 8959
rect 24593 8925 24627 8959
rect 24685 8925 24719 8959
rect 24961 8925 24995 8959
rect 25605 8925 25639 8959
rect 25789 8925 25823 8959
rect 25973 8925 26007 8959
rect 29561 8925 29595 8959
rect 29817 8925 29851 8959
rect 31585 8925 31619 8959
rect 31769 8925 31803 8959
rect 31953 8925 31987 8959
rect 32689 8925 32723 8959
rect 33057 8925 33091 8959
rect 33793 8925 33827 8959
rect 33885 8925 33919 8959
rect 33977 8925 34011 8959
rect 34161 8925 34195 8959
rect 68109 8925 68143 8959
rect 3985 8857 4019 8891
rect 5724 8857 5758 8891
rect 7297 8857 7331 8891
rect 12173 8857 12207 8891
rect 19717 8857 19751 8891
rect 24777 8857 24811 8891
rect 25881 8857 25915 8891
rect 27537 8857 27571 8891
rect 27721 8857 27755 8891
rect 31677 8857 31711 8891
rect 32781 8857 32815 8891
rect 32873 8857 32907 8891
rect 36378 8857 36412 8891
rect 3157 8789 3191 8823
rect 4169 8789 4203 8823
rect 11069 8789 11103 8823
rect 11713 8789 11747 8823
rect 12817 8789 12851 8823
rect 13461 8789 13495 8823
rect 14657 8789 14691 8823
rect 15853 8789 15887 8823
rect 18613 8789 18647 8823
rect 20821 8789 20855 8823
rect 30941 8789 30975 8823
rect 32505 8789 32539 8823
rect 35265 8789 35299 8823
rect 4813 8585 4847 8619
rect 7573 8585 7607 8619
rect 8125 8585 8159 8619
rect 21833 8585 21867 8619
rect 25697 8585 25731 8619
rect 29377 8585 29411 8619
rect 32137 8585 32171 8619
rect 33977 8585 34011 8619
rect 37381 8585 37415 8619
rect 7389 8517 7423 8551
rect 18806 8517 18840 8551
rect 22946 8517 22980 8551
rect 24409 8517 24443 8551
rect 25973 8517 26007 8551
rect 27445 8517 27479 8551
rect 27629 8517 27663 8551
rect 28733 8517 28767 8551
rect 30490 8517 30524 8551
rect 33793 8517 33827 8551
rect 35725 8517 35759 8551
rect 36369 8517 36403 8551
rect 2329 8449 2363 8483
rect 2513 8449 2547 8483
rect 2605 8449 2639 8483
rect 2697 8449 2731 8483
rect 3433 8449 3467 8483
rect 3689 8449 3723 8483
rect 7205 8449 7239 8483
rect 10721 8449 10755 8483
rect 10977 8449 11011 8483
rect 11713 8449 11747 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 14022 8449 14056 8483
rect 15117 8449 15151 8483
rect 20453 8449 20487 8483
rect 23213 8449 23247 8483
rect 24225 8449 24259 8483
rect 25881 8449 25915 8483
rect 26065 8449 26099 8483
rect 26249 8449 26283 8483
rect 27261 8449 27295 8483
rect 28089 8449 28123 8483
rect 28273 8449 28307 8483
rect 28365 8449 28399 8483
rect 28457 8449 28491 8483
rect 32321 8449 32355 8483
rect 32413 8449 32447 8483
rect 32505 8449 32539 8483
rect 32689 8449 32723 8483
rect 33609 8449 33643 8483
rect 35541 8449 35575 8483
rect 38494 8449 38528 8483
rect 38761 8449 38795 8483
rect 2973 8381 3007 8415
rect 11529 8381 11563 8415
rect 11897 8381 11931 8415
rect 11989 8381 12023 8415
rect 14289 8381 14323 8415
rect 14841 8381 14875 8415
rect 19073 8381 19107 8415
rect 20177 8381 20211 8415
rect 24593 8381 24627 8415
rect 30757 8381 30791 8415
rect 5825 8313 5859 8347
rect 6653 8313 6687 8347
rect 9045 8313 9079 8347
rect 9597 8313 9631 8347
rect 17049 8313 17083 8347
rect 17693 8313 17727 8347
rect 12909 8245 12943 8279
rect 25145 8245 25179 8279
rect 35909 8245 35943 8279
rect 3157 8041 3191 8075
rect 13277 8041 13311 8075
rect 26985 8041 27019 8075
rect 28917 8041 28951 8075
rect 31493 8041 31527 8075
rect 33425 8041 33459 8075
rect 34161 8041 34195 8075
rect 36829 8041 36863 8075
rect 14841 7973 14875 8007
rect 22293 7973 22327 8007
rect 5733 7905 5767 7939
rect 7941 7905 7975 7939
rect 9229 7905 9263 7939
rect 12817 7905 12851 7939
rect 17877 7905 17911 7939
rect 20361 7905 20395 7939
rect 35357 7905 35391 7939
rect 35633 7905 35667 7939
rect 5089 7837 5123 7871
rect 7757 7837 7791 7871
rect 8953 7837 8987 7871
rect 11253 7837 11287 7871
rect 11897 7837 11931 7871
rect 12541 7837 12575 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13093 7837 13127 7871
rect 15301 7837 15335 7871
rect 17601 7837 17635 7871
rect 17785 7831 17819 7865
rect 17969 7837 18003 7871
rect 18153 7837 18187 7871
rect 20085 7837 20119 7871
rect 21465 7837 21499 7871
rect 22017 7837 22051 7871
rect 22201 7837 22235 7871
rect 24961 7837 24995 7871
rect 25053 7837 25087 7871
rect 25145 7837 25179 7871
rect 25329 7837 25363 7871
rect 26065 7837 26099 7871
rect 26157 7837 26191 7871
rect 26249 7837 26283 7871
rect 26433 7837 26467 7871
rect 27813 7837 27847 7871
rect 27905 7837 27939 7871
rect 27997 7837 28031 7871
rect 28181 7837 28215 7871
rect 31677 7837 31711 7871
rect 32045 7837 32079 7871
rect 33977 7837 34011 7871
rect 36185 7837 36219 7871
rect 36369 7837 36403 7871
rect 36464 7831 36498 7865
rect 36553 7837 36587 7871
rect 68109 7837 68143 7871
rect 2513 7769 2547 7803
rect 5978 7769 6012 7803
rect 7573 7769 7607 7803
rect 10609 7769 10643 7803
rect 14657 7769 14691 7803
rect 31769 7769 31803 7803
rect 31861 7769 31895 7803
rect 1501 7701 1535 7735
rect 2053 7701 2087 7735
rect 3893 7701 3927 7735
rect 4629 7701 4663 7735
rect 5273 7701 5307 7735
rect 7113 7701 7147 7735
rect 11069 7701 11103 7735
rect 11989 7701 12023 7735
rect 16589 7701 16623 7735
rect 18337 7701 18371 7735
rect 24685 7701 24719 7735
rect 25789 7701 25823 7735
rect 27537 7701 27571 7735
rect 2421 7497 2455 7531
rect 7389 7497 7423 7531
rect 7849 7497 7883 7531
rect 20085 7497 20119 7531
rect 21189 7497 21223 7531
rect 26433 7497 26467 7531
rect 27813 7497 27847 7531
rect 37841 7497 37875 7531
rect 3402 7429 3436 7463
rect 5641 7429 5675 7463
rect 9904 7429 9938 7463
rect 11897 7429 11931 7463
rect 20729 7429 20763 7463
rect 23949 7429 23983 7463
rect 25605 7429 25639 7463
rect 27629 7429 27663 7463
rect 30941 7429 30975 7463
rect 32597 7429 32631 7463
rect 32781 7429 32815 7463
rect 2237 7361 2271 7395
rect 6929 7361 6963 7395
rect 7757 7361 7791 7395
rect 10149 7361 10183 7395
rect 10793 7361 10827 7395
rect 12173 7361 12207 7395
rect 12262 7361 12296 7395
rect 12378 7361 12412 7395
rect 12541 7361 12575 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 18254 7361 18288 7395
rect 20453 7361 20487 7395
rect 21833 7361 21867 7395
rect 22017 7361 22051 7395
rect 26065 7361 26099 7395
rect 26249 7361 26283 7395
rect 27445 7361 27479 7395
rect 31125 7361 31159 7395
rect 33793 7361 33827 7395
rect 35265 7361 35299 7395
rect 35909 7361 35943 7395
rect 36088 7361 36122 7395
rect 36188 7364 36222 7398
rect 36297 7361 36331 7395
rect 38669 7361 38703 7395
rect 38761 7361 38795 7395
rect 38853 7361 38887 7395
rect 39037 7361 39071 7395
rect 3157 7293 3191 7327
rect 4997 7293 5031 7327
rect 5365 7293 5399 7327
rect 5457 7293 5491 7327
rect 7941 7293 7975 7327
rect 13553 7293 13587 7327
rect 13829 7293 13863 7327
rect 18521 7293 18555 7327
rect 20545 7293 20579 7327
rect 34989 7293 35023 7327
rect 1777 7225 1811 7259
rect 22109 7225 22143 7259
rect 4537 7157 4571 7191
rect 8769 7157 8803 7191
rect 10977 7157 11011 7191
rect 16129 7157 16163 7191
rect 17141 7157 17175 7191
rect 18981 7157 19015 7191
rect 23305 7157 23339 7191
rect 28365 7157 28399 7191
rect 30297 7157 30331 7191
rect 30757 7157 30791 7191
rect 32413 7157 32447 7191
rect 33977 7157 34011 7191
rect 36553 7157 36587 7191
rect 38393 7157 38427 7191
rect 23857 6953 23891 6987
rect 26801 6953 26835 6987
rect 30941 6953 30975 6987
rect 32413 6953 32447 6987
rect 39129 6953 39163 6987
rect 36277 6885 36311 6919
rect 2329 6817 2363 6851
rect 5641 6817 5675 6851
rect 7205 6817 7239 6851
rect 9321 6817 9355 6851
rect 10149 6817 10183 6851
rect 10971 6817 11005 6851
rect 12725 6817 12759 6851
rect 14933 6817 14967 6851
rect 17233 6817 17267 6851
rect 19257 6817 19291 6851
rect 35725 6817 35759 6851
rect 2237 6749 2271 6783
rect 5365 6749 5399 6783
rect 5457 6749 5491 6783
rect 8217 6749 8251 6783
rect 9413 6749 9447 6783
rect 10057 6749 10091 6783
rect 10701 6749 10735 6783
rect 10885 6749 10919 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11897 6749 11931 6783
rect 13185 6749 13219 6783
rect 14565 6749 14599 6783
rect 14749 6749 14783 6783
rect 14841 6749 14875 6783
rect 15117 6749 15151 6783
rect 17969 6749 18003 6783
rect 18153 6749 18187 6783
rect 18245 6749 18279 6783
rect 18337 6749 18371 6783
rect 18521 6749 18555 6783
rect 21281 6749 21315 6783
rect 22477 6749 22511 6783
rect 25421 6749 25455 6783
rect 25688 6749 25722 6783
rect 28374 6749 28408 6783
rect 28641 6749 28675 6783
rect 29561 6749 29595 6783
rect 33793 6749 33827 6783
rect 35357 6749 35391 6783
rect 36921 6749 36955 6783
rect 38945 6749 38979 6783
rect 2145 6681 2179 6715
rect 2973 6681 3007 6715
rect 4537 6681 4571 6715
rect 9597 6681 9631 6715
rect 15301 6681 15335 6715
rect 16966 6681 17000 6715
rect 18705 6681 18739 6715
rect 19502 6681 19536 6715
rect 21465 6681 21499 6715
rect 22744 6681 22778 6715
rect 24777 6681 24811 6715
rect 24961 6681 24995 6715
rect 29828 6681 29862 6715
rect 31401 6681 31435 6715
rect 31585 6681 31619 6715
rect 33526 6681 33560 6715
rect 35541 6681 35575 6715
rect 37166 6681 37200 6715
rect 38761 6681 38795 6715
rect 1777 6613 1811 6647
rect 3985 6613 4019 6647
rect 4997 6613 5031 6647
rect 6653 6613 6687 6647
rect 7757 6613 7791 6647
rect 8401 6613 8435 6647
rect 8953 6613 8987 6647
rect 11437 6613 11471 6647
rect 12081 6613 12115 6647
rect 13369 6613 13403 6647
rect 15853 6613 15887 6647
rect 20637 6613 20671 6647
rect 21097 6613 21131 6647
rect 27261 6613 27295 6647
rect 31769 6613 31803 6647
rect 38301 6613 38335 6647
rect 2145 6409 2179 6443
rect 2789 6409 2823 6443
rect 7757 6409 7791 6443
rect 14749 6409 14783 6443
rect 17877 6409 17911 6443
rect 22017 6409 22051 6443
rect 25605 6409 25639 6443
rect 26249 6409 26283 6443
rect 30573 6409 30607 6443
rect 32965 6409 32999 6443
rect 15393 6341 15427 6375
rect 17233 6341 17267 6375
rect 21281 6341 21315 6375
rect 23130 6341 23164 6375
rect 33701 6341 33735 6375
rect 1961 6273 1995 6307
rect 3341 6273 3375 6307
rect 5825 6273 5859 6307
rect 6633 6273 6667 6307
rect 8401 6273 8435 6307
rect 9689 6273 9723 6307
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 10793 6273 10827 6307
rect 12642 6273 12676 6307
rect 12909 6273 12943 6307
rect 13737 6273 13771 6307
rect 14933 6273 14967 6307
rect 17601 6273 17635 6307
rect 20637 6273 20671 6307
rect 20816 6279 20850 6313
rect 20913 6273 20947 6307
rect 21005 6273 21039 6307
rect 23397 6273 23431 6307
rect 24492 6273 24526 6307
rect 26157 6273 26191 6307
rect 27997 6273 28031 6307
rect 30849 6273 30883 6307
rect 30941 6273 30975 6307
rect 31033 6273 31067 6307
rect 31217 6273 31251 6307
rect 32321 6273 32355 6307
rect 32500 6273 32534 6307
rect 32597 6273 32631 6307
rect 32689 6273 32723 6307
rect 33517 6273 33551 6307
rect 35495 6273 35529 6307
rect 35633 6273 35667 6307
rect 35746 6273 35780 6307
rect 35909 6273 35943 6307
rect 1777 6205 1811 6239
rect 3801 6205 3835 6239
rect 4169 6205 4203 6239
rect 4261 6205 4295 6239
rect 6377 6205 6411 6239
rect 9413 6205 9447 6239
rect 13461 6205 13495 6239
rect 15025 6205 15059 6239
rect 17693 6205 17727 6239
rect 20085 6205 20119 6239
rect 24225 6205 24259 6239
rect 26985 6205 27019 6239
rect 34713 6205 34747 6239
rect 10977 6137 11011 6171
rect 29285 6137 29319 6171
rect 67649 6137 67683 6171
rect 4445 6069 4479 6103
rect 5181 6069 5215 6103
rect 5641 6069 5675 6103
rect 8217 6069 8251 6103
rect 10333 6069 10367 6103
rect 11529 6069 11563 6103
rect 16129 6069 16163 6103
rect 16773 6069 16807 6103
rect 18705 6069 18739 6103
rect 19349 6069 19383 6103
rect 33885 6069 33919 6103
rect 35265 6069 35299 6103
rect 1593 5865 1627 5899
rect 6285 5865 6319 5899
rect 7389 5865 7423 5899
rect 12081 5865 12115 5899
rect 14749 5865 14783 5899
rect 18061 5865 18095 5899
rect 19257 5865 19291 5899
rect 22293 5865 22327 5899
rect 24409 5865 24443 5899
rect 26341 5865 26375 5899
rect 26893 5865 26927 5899
rect 27537 5865 27571 5899
rect 29561 5865 29595 5899
rect 32965 5865 32999 5899
rect 38761 5865 38795 5899
rect 10977 5797 11011 5831
rect 12725 5797 12759 5831
rect 2605 5729 2639 5763
rect 6745 5729 6779 5763
rect 7205 5729 7239 5763
rect 10425 5729 10459 5763
rect 14473 5729 14507 5763
rect 14565 5729 14599 5763
rect 15301 5729 15335 5763
rect 16497 5729 16531 5763
rect 18245 5729 18279 5763
rect 19441 5729 19475 5763
rect 19533 5729 19567 5763
rect 20361 5729 20395 5763
rect 22937 5729 22971 5763
rect 23213 5729 23247 5763
rect 30941 5729 30975 5763
rect 5181 5661 5215 5695
rect 6101 5661 6135 5695
rect 7113 5661 7147 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 12817 5661 12851 5695
rect 13553 5661 13587 5695
rect 14105 5661 14139 5695
rect 15209 5661 15243 5695
rect 15393 5661 15427 5695
rect 17601 5661 17635 5695
rect 18337 5661 18371 5695
rect 20637 5661 20671 5695
rect 21649 5661 21683 5695
rect 24639 5661 24673 5695
rect 24777 5661 24811 5695
rect 24869 5661 24903 5695
rect 25053 5661 25087 5695
rect 25697 5661 25731 5695
rect 27997 5661 28031 5695
rect 28176 5661 28210 5695
rect 28276 5655 28310 5689
rect 28365 5661 28399 5695
rect 31677 5661 31711 5695
rect 31766 5658 31800 5692
rect 31866 5661 31900 5695
rect 32045 5661 32079 5695
rect 33793 5661 33827 5695
rect 33885 5661 33919 5695
rect 33977 5661 34011 5695
rect 34161 5661 34195 5695
rect 37381 5661 37415 5695
rect 37648 5661 37682 5695
rect 2421 5593 2455 5627
rect 4914 5593 4948 5627
rect 7941 5593 7975 5627
rect 10241 5593 10275 5627
rect 10977 5593 11011 5627
rect 12541 5593 12575 5627
rect 16129 5593 16163 5627
rect 16589 5593 16623 5627
rect 18705 5593 18739 5627
rect 19901 5593 19935 5627
rect 25513 5593 25547 5627
rect 25881 5593 25915 5627
rect 28641 5593 28675 5627
rect 30674 5593 30708 5627
rect 35081 5593 35115 5627
rect 36829 5593 36863 5627
rect 2053 5525 2087 5559
rect 2513 5525 2547 5559
rect 3801 5525 3835 5559
rect 10517 5525 10551 5559
rect 12817 5525 12851 5559
rect 16405 5525 16439 5559
rect 16773 5525 16807 5559
rect 21833 5525 21867 5559
rect 31401 5525 31435 5559
rect 33517 5525 33551 5559
rect 2789 5321 2823 5355
rect 4445 5321 4479 5355
rect 5089 5321 5123 5355
rect 7481 5321 7515 5355
rect 8677 5321 8711 5355
rect 9045 5321 9079 5355
rect 9137 5321 9171 5355
rect 10977 5321 11011 5355
rect 15117 5321 15151 5355
rect 16957 5321 16991 5355
rect 20729 5321 20763 5355
rect 21833 5321 21867 5355
rect 24961 5321 24995 5355
rect 29653 5321 29687 5355
rect 37289 5321 37323 5355
rect 11529 5253 11563 5287
rect 17141 5253 17175 5287
rect 17417 5253 17451 5287
rect 26065 5253 26099 5287
rect 26249 5253 26283 5287
rect 28273 5253 28307 5287
rect 32229 5253 32263 5287
rect 33793 5253 33827 5287
rect 33977 5253 34011 5287
rect 34161 5253 34195 5287
rect 38117 5253 38151 5287
rect 38301 5253 38335 5287
rect 1777 5185 1811 5219
rect 1961 5185 1995 5219
rect 2145 5185 2179 5219
rect 2605 5185 2639 5219
rect 4905 5185 4939 5219
rect 5641 5185 5675 5219
rect 6653 5185 6687 5219
rect 7297 5185 7331 5219
rect 8125 5185 8159 5219
rect 10149 5185 10183 5219
rect 10793 5185 10827 5219
rect 11989 5185 12023 5219
rect 13277 5185 13311 5219
rect 13921 5185 13955 5219
rect 14657 5185 14691 5219
rect 14933 5185 14967 5219
rect 15301 5185 15335 5219
rect 17049 5185 17083 5219
rect 18981 5185 19015 5219
rect 19625 5185 19659 5219
rect 20637 5185 20671 5219
rect 22946 5185 22980 5219
rect 23213 5185 23247 5219
rect 23673 5185 23707 5219
rect 23949 5185 23983 5219
rect 26985 5185 27019 5219
rect 27148 5185 27182 5219
rect 27261 5185 27295 5219
rect 27353 5185 27387 5219
rect 28089 5185 28123 5219
rect 28457 5185 28491 5219
rect 31318 5185 31352 5219
rect 31585 5185 31619 5219
rect 34713 5185 34747 5219
rect 34897 5185 34931 5219
rect 34989 5185 35023 5219
rect 35081 5185 35115 5219
rect 36001 5185 36035 5219
rect 36185 5185 36219 5219
rect 36277 5185 36311 5219
rect 36369 5185 36403 5219
rect 37473 5185 37507 5219
rect 37657 5185 37691 5219
rect 38485 5185 38519 5219
rect 4813 5117 4847 5151
rect 9321 5117 9355 5151
rect 11897 5117 11931 5151
rect 13461 5117 13495 5151
rect 16681 5117 16715 5151
rect 18521 5117 18555 5151
rect 20821 5117 20855 5151
rect 26433 5117 26467 5151
rect 59461 5117 59495 5151
rect 3985 5049 4019 5083
rect 6837 5049 6871 5083
rect 10333 5049 10367 5083
rect 13093 5049 13127 5083
rect 16129 5049 16163 5083
rect 30205 5049 30239 5083
rect 60105 5049 60139 5083
rect 3433 4981 3467 5015
rect 5825 4981 5859 5015
rect 8033 4981 8067 5015
rect 11621 4981 11655 5015
rect 12173 4981 12207 5015
rect 14105 4981 14139 5015
rect 14841 4981 14875 5015
rect 19165 4981 19199 5015
rect 19809 4981 19843 5015
rect 20269 4981 20303 5015
rect 27629 4981 27663 5015
rect 35357 4981 35391 5015
rect 36645 4981 36679 5015
rect 58817 4981 58851 5015
rect 67649 4981 67683 5015
rect 5641 4777 5675 4811
rect 10425 4777 10459 4811
rect 14657 4777 14691 4811
rect 21189 4777 21223 4811
rect 23581 4777 23615 4811
rect 31217 4777 31251 4811
rect 32137 4777 32171 4811
rect 34897 4777 34931 4811
rect 38669 4777 38703 4811
rect 4261 4709 4295 4743
rect 9045 4709 9079 4743
rect 12173 4709 12207 4743
rect 18613 4709 18647 4743
rect 25789 4709 25823 4743
rect 57897 4709 57931 4743
rect 59185 4709 59219 4743
rect 1593 4641 1627 4675
rect 10425 4641 10459 4675
rect 12265 4641 12299 4675
rect 17969 4641 18003 4675
rect 21649 4641 21683 4675
rect 24409 4641 24443 4675
rect 60473 4641 60507 4675
rect 2605 4573 2639 4607
rect 4077 4573 4111 4607
rect 4721 4573 4755 4607
rect 7113 4573 7147 4607
rect 8125 4573 8159 4607
rect 9689 4573 9723 4607
rect 10701 4573 10735 4607
rect 11161 4573 11195 4607
rect 12044 4573 12078 4607
rect 13553 4573 13587 4607
rect 14473 4573 14507 4607
rect 14749 4573 14783 4607
rect 15117 4573 15151 4607
rect 15577 4573 15611 4607
rect 16865 4573 16899 4607
rect 17785 4573 17819 4607
rect 19717 4573 19751 4607
rect 20177 4573 20211 4607
rect 20361 4573 20395 4607
rect 20545 4573 20579 4607
rect 21005 4573 21039 4607
rect 26433 4573 26467 4607
rect 28457 4573 28491 4607
rect 33517 4573 33551 4607
rect 35449 4573 35483 4607
rect 35716 4573 35750 4607
rect 37289 4573 37323 4607
rect 37545 4573 37579 4607
rect 57253 4573 57287 4607
rect 58541 4573 58575 4607
rect 11897 4505 11931 4539
rect 12633 4505 12667 4539
rect 22845 4505 22879 4539
rect 24676 4505 24710 4539
rect 26617 4505 26651 4539
rect 28273 4505 28307 4539
rect 33272 4505 33306 4539
rect 2145 4437 2179 4471
rect 2789 4437 2823 4471
rect 4905 4437 4939 4471
rect 8033 4437 8067 4471
rect 10149 4437 10183 4471
rect 11345 4437 11379 4471
rect 13369 4437 13403 4471
rect 14933 4437 14967 4471
rect 15761 4437 15795 4471
rect 16681 4437 16715 4471
rect 17417 4437 17451 4471
rect 17877 4437 17911 4471
rect 22293 4437 22327 4471
rect 26249 4437 26283 4471
rect 28641 4437 28675 4471
rect 34069 4437 34103 4471
rect 36829 4437 36863 4471
rect 2053 4233 2087 4267
rect 8493 4233 8527 4267
rect 8861 4233 8895 4267
rect 8953 4233 8987 4267
rect 10717 4233 10751 4267
rect 10885 4233 10919 4267
rect 12173 4233 12207 4267
rect 14473 4233 14507 4267
rect 17325 4233 17359 4267
rect 26985 4233 27019 4267
rect 29469 4233 29503 4267
rect 33793 4233 33827 4267
rect 35909 4233 35943 4267
rect 3586 4165 3620 4199
rect 5641 4165 5675 4199
rect 7021 4165 7055 4199
rect 10517 4165 10551 4199
rect 11621 4165 11655 4199
rect 20821 4165 20855 4199
rect 20913 4165 20947 4199
rect 28098 4165 28132 4199
rect 3341 4097 3375 4131
rect 7205 4097 7239 4131
rect 7665 4097 7699 4131
rect 7849 4097 7883 4131
rect 7941 4097 7975 4131
rect 9873 4097 9907 4131
rect 13277 4097 13311 4131
rect 14013 4097 14047 4131
rect 14841 4097 14875 4131
rect 15577 4097 15611 4131
rect 17509 4097 17543 4131
rect 17693 4097 17727 4131
rect 18797 4097 18831 4131
rect 19441 4097 19475 4131
rect 19625 4097 19659 4131
rect 21833 4097 21867 4131
rect 23590 4097 23624 4131
rect 23857 4097 23891 4131
rect 25467 4097 25501 4131
rect 25605 4097 25639 4131
rect 25697 4100 25731 4134
rect 25881 4097 25915 4131
rect 28365 4097 28399 4131
rect 28825 4097 28859 4131
rect 30582 4097 30616 4131
rect 30849 4097 30883 4131
rect 34906 4097 34940 4131
rect 35173 4097 35207 4131
rect 59829 4097 59863 4131
rect 1869 4029 1903 4063
rect 1961 4029 1995 4063
rect 9045 4029 9079 4063
rect 10057 4029 10091 4063
rect 12081 4029 12115 4063
rect 14749 4029 14783 4063
rect 16037 4029 16071 4063
rect 20729 4029 20763 4063
rect 25237 4029 25271 4063
rect 61117 4029 61151 4063
rect 5825 3961 5859 3995
rect 11621 3961 11655 3995
rect 15393 3961 15427 3995
rect 18337 3961 18371 3995
rect 19625 3961 19659 3995
rect 22017 3961 22051 3995
rect 58541 3961 58575 3995
rect 60473 3961 60507 3995
rect 2421 3893 2455 3927
rect 4721 3893 4755 3927
rect 6469 3893 6503 3927
rect 9689 3893 9723 3927
rect 10701 3893 10735 3927
rect 12357 3893 12391 3927
rect 13093 3893 13127 3927
rect 13829 3893 13863 3927
rect 14841 3893 14875 3927
rect 16865 3893 16899 3927
rect 18981 3893 19015 3927
rect 21281 3893 21315 3927
rect 22477 3893 22511 3927
rect 24685 3893 24719 3927
rect 56241 3893 56275 3927
rect 56885 3893 56919 3927
rect 57897 3893 57931 3927
rect 59185 3893 59219 3927
rect 2329 3689 2363 3723
rect 6745 3689 6779 3723
rect 10609 3689 10643 3723
rect 13553 3689 13587 3723
rect 17049 3689 17083 3723
rect 20085 3689 20119 3723
rect 21189 3689 21223 3723
rect 29009 3689 29043 3723
rect 3249 3621 3283 3655
rect 9781 3621 9815 3655
rect 12817 3621 12851 3655
rect 18705 3621 18739 3655
rect 19349 3621 19383 3655
rect 41797 3621 41831 3655
rect 57897 3621 57931 3655
rect 61117 3621 61151 3655
rect 1961 3553 1995 3587
rect 4629 3553 4663 3587
rect 4721 3553 4755 3587
rect 7665 3553 7699 3587
rect 7849 3553 7883 3587
rect 13369 3553 13403 3587
rect 15669 3553 15703 3587
rect 19809 3553 19843 3587
rect 19901 3553 19935 3587
rect 20821 3553 20855 3587
rect 56609 3553 56643 3587
rect 58541 3553 58575 3587
rect 61761 3553 61795 3587
rect 2145 3485 2179 3519
rect 3065 3485 3099 3519
rect 5365 3485 5399 3519
rect 5632 3485 5666 3519
rect 7573 3485 7607 3519
rect 9229 3485 9263 3519
rect 9965 3485 9999 3519
rect 11253 3485 11287 3519
rect 11529 3485 11563 3519
rect 14473 3485 14507 3519
rect 15936 3485 15970 3519
rect 18061 3485 18095 3519
rect 18521 3485 18555 3519
rect 21005 3485 21039 3519
rect 21925 3485 21959 3519
rect 22753 3485 22787 3519
rect 23581 3485 23615 3519
rect 24409 3485 24443 3519
rect 25237 3485 25271 3519
rect 26065 3485 26099 3519
rect 26893 3485 26927 3519
rect 27721 3485 27755 3519
rect 28365 3485 28399 3519
rect 28549 3485 28583 3519
rect 28641 3485 28675 3519
rect 28733 3485 28767 3519
rect 29929 3485 29963 3519
rect 30757 3485 30791 3519
rect 31585 3485 31619 3519
rect 32413 3485 32447 3519
rect 33241 3485 33275 3519
rect 39865 3485 39899 3519
rect 40509 3485 40543 3519
rect 41153 3485 41187 3519
rect 42625 3485 42659 3519
rect 43269 3485 43303 3519
rect 45109 3485 45143 3519
rect 45753 3485 45787 3519
rect 46397 3485 46431 3519
rect 47041 3485 47075 3519
rect 47869 3485 47903 3519
rect 48973 3485 49007 3519
rect 50353 3485 50387 3519
rect 50997 3485 51031 3519
rect 51641 3485 51675 3519
rect 52837 3485 52871 3519
rect 53481 3485 53515 3519
rect 55321 3485 55355 3519
rect 55965 3485 55999 3519
rect 57253 3485 57287 3519
rect 59185 3485 59219 3519
rect 60473 3485 60507 3519
rect 68109 3485 68143 3519
rect 1501 3417 1535 3451
rect 4537 3417 4571 3451
rect 10593 3417 10627 3451
rect 10793 3417 10827 3451
rect 12817 3417 12851 3451
rect 19349 3417 19383 3451
rect 4169 3349 4203 3383
rect 7205 3349 7239 3383
rect 9045 3349 9079 3383
rect 10425 3349 10459 3383
rect 13277 3349 13311 3383
rect 14657 3349 14691 3383
rect 5457 3145 5491 3179
rect 7757 3145 7791 3179
rect 11897 3145 11931 3179
rect 16773 3145 16807 3179
rect 21833 3145 21867 3179
rect 10885 3077 10919 3111
rect 13369 3077 13403 3111
rect 1501 3009 1535 3043
rect 2145 3009 2179 3043
rect 2329 3009 2363 3043
rect 3433 3009 3467 3043
rect 3689 3009 3723 3043
rect 5641 3009 5675 3043
rect 6377 3009 6411 3043
rect 6633 3009 6667 3043
rect 8217 3009 8251 3043
rect 8484 3009 8518 3043
rect 12725 3009 12759 3043
rect 13826 3009 13860 3043
rect 14473 3009 14507 3043
rect 14749 3009 14783 3043
rect 15761 3009 15795 3043
rect 16957 3009 16991 3043
rect 17417 3009 17451 3043
rect 61117 3009 61151 3043
rect 2513 2941 2547 2975
rect 5825 2941 5859 2975
rect 10609 2941 10643 2975
rect 12173 2941 12207 2975
rect 13645 2941 13679 2975
rect 14565 2941 14599 2975
rect 18705 2941 18739 2975
rect 20637 2941 20671 2975
rect 37933 2941 37967 2975
rect 45661 2941 45695 2975
rect 49525 2941 49559 2975
rect 53389 2941 53423 2975
rect 61761 2941 61795 2975
rect 1685 2873 1719 2907
rect 4813 2873 4847 2907
rect 12265 2873 12299 2907
rect 15577 2873 15611 2907
rect 17601 2873 17635 2907
rect 19349 2873 19383 2907
rect 39221 2873 39255 2907
rect 40509 2873 40543 2907
rect 43085 2873 43119 2907
rect 44373 2873 44407 2907
rect 48237 2873 48271 2907
rect 50169 2873 50203 2907
rect 51457 2873 51491 2907
rect 54033 2873 54067 2907
rect 55321 2873 55355 2907
rect 56609 2873 56643 2907
rect 58541 2873 58575 2907
rect 63049 2873 63083 2907
rect 9597 2805 9631 2839
rect 12357 2805 12391 2839
rect 13737 2805 13771 2839
rect 14013 2805 14047 2839
rect 14473 2805 14507 2839
rect 14933 2805 14967 2839
rect 19993 2805 20027 2839
rect 21281 2805 21315 2839
rect 22569 2805 22603 2839
rect 23213 2805 23247 2839
rect 23857 2805 23891 2839
rect 24501 2805 24535 2839
rect 25145 2805 25179 2839
rect 25789 2805 25823 2839
rect 26433 2805 26467 2839
rect 27721 2805 27755 2839
rect 28365 2805 28399 2839
rect 29009 2805 29043 2839
rect 29653 2805 29687 2839
rect 30297 2805 30331 2839
rect 30941 2805 30975 2839
rect 31585 2805 31619 2839
rect 32873 2805 32907 2839
rect 33517 2805 33551 2839
rect 34161 2805 34195 2839
rect 34621 2805 34655 2839
rect 35449 2805 35483 2839
rect 36277 2805 36311 2839
rect 37289 2805 37323 2839
rect 38577 2805 38611 2839
rect 39865 2805 39899 2839
rect 41153 2805 41187 2839
rect 42441 2805 42475 2839
rect 43729 2805 43763 2839
rect 45017 2805 45051 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48881 2805 48915 2839
rect 50813 2805 50847 2839
rect 52745 2805 52779 2839
rect 54677 2805 54711 2839
rect 55965 2805 55999 2839
rect 57897 2805 57931 2839
rect 59185 2805 59219 2839
rect 59829 2805 59863 2839
rect 60473 2805 60507 2839
rect 4537 2601 4571 2635
rect 5825 2601 5859 2635
rect 6837 2601 6871 2635
rect 9505 2601 9539 2635
rect 11621 2601 11655 2635
rect 11989 2601 12023 2635
rect 14841 2601 14875 2635
rect 16773 2601 16807 2635
rect 19349 2601 19383 2635
rect 21833 2601 21867 2635
rect 26985 2601 27019 2635
rect 55321 2601 55355 2635
rect 61117 2601 61151 2635
rect 2605 2533 2639 2567
rect 8217 2533 8251 2567
rect 12081 2533 12115 2567
rect 15853 2533 15887 2567
rect 18245 2533 18279 2567
rect 20637 2533 20671 2567
rect 22569 2533 22603 2567
rect 25789 2533 25823 2567
rect 28365 2533 28399 2567
rect 30297 2533 30331 2567
rect 42441 2533 42475 2567
rect 46305 2533 46339 2567
rect 50169 2533 50203 2567
rect 54033 2533 54067 2567
rect 57897 2533 57931 2567
rect 58541 2533 58575 2567
rect 60473 2533 60507 2567
rect 10701 2465 10735 2499
rect 11897 2465 11931 2499
rect 24409 2465 24443 2499
rect 25145 2465 25179 2499
rect 37933 2465 37967 2499
rect 39865 2465 39899 2499
rect 43085 2465 43119 2499
rect 45017 2465 45051 2499
rect 48237 2465 48271 2499
rect 50813 2465 50847 2499
rect 52745 2465 52779 2499
rect 56609 2465 56643 2499
rect 63693 2465 63727 2499
rect 1777 2397 1811 2431
rect 2421 2397 2455 2431
rect 3065 2397 3099 2431
rect 4353 2397 4387 2431
rect 5181 2397 5215 2431
rect 5641 2397 5675 2431
rect 6653 2397 6687 2431
rect 7665 2397 7699 2431
rect 8401 2397 8435 2431
rect 9689 2397 9723 2431
rect 10977 2397 11011 2431
rect 12449 2397 12483 2431
rect 13001 2397 13035 2431
rect 13369 2397 13403 2431
rect 16037 2397 16071 2431
rect 16865 2397 16899 2431
rect 17693 2397 17727 2431
rect 18429 2397 18463 2431
rect 19993 2397 20027 2431
rect 21281 2397 21315 2431
rect 23213 2397 23247 2431
rect 23857 2397 23891 2431
rect 26433 2397 26467 2431
rect 27721 2397 27755 2431
rect 29009 2397 29043 2431
rect 30941 2397 30975 2431
rect 31585 2397 31619 2431
rect 32873 2397 32907 2431
rect 33517 2397 33551 2431
rect 34161 2397 34195 2431
rect 34897 2397 34931 2431
rect 35541 2397 35575 2431
rect 36001 2397 36035 2431
rect 37289 2397 37323 2431
rect 38577 2397 38611 2431
rect 40509 2397 40543 2431
rect 41153 2397 41187 2431
rect 43729 2397 43763 2431
rect 45661 2397 45695 2431
rect 47593 2397 47627 2431
rect 48881 2397 48915 2431
rect 51457 2397 51491 2431
rect 53389 2397 53423 2431
rect 55965 2397 55999 2431
rect 59185 2397 59219 2431
rect 61761 2397 61795 2431
rect 63049 2397 63083 2431
rect 67005 2397 67039 2431
rect 67649 2397 67683 2431
rect 14565 2329 14599 2363
rect 1961 2261 1995 2295
rect 3249 2261 3283 2295
rect 3893 2261 3927 2295
rect 7481 2261 7515 2295
rect 17509 2261 17543 2295
<< metal1 >>
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 5166 57400 5172 57452
rect 5224 57440 5230 57452
rect 5261 57443 5319 57449
rect 5261 57440 5273 57443
rect 5224 57412 5273 57440
rect 5224 57400 5230 57412
rect 5261 57409 5273 57412
rect 5307 57409 5319 57443
rect 15194 57440 15200 57452
rect 15155 57412 15200 57440
rect 5261 57403 5319 57409
rect 15194 57400 15200 57412
rect 15252 57400 15258 57452
rect 25038 57400 25044 57452
rect 25096 57440 25102 57452
rect 25133 57443 25191 57449
rect 25133 57440 25145 57443
rect 25096 57412 25145 57440
rect 25096 57400 25102 57412
rect 25133 57409 25145 57412
rect 25179 57409 25191 57443
rect 25133 57403 25191 57409
rect 34974 57400 34980 57452
rect 35032 57440 35038 57452
rect 35069 57443 35127 57449
rect 35069 57440 35081 57443
rect 35032 57412 35081 57440
rect 35032 57400 35038 57412
rect 35069 57409 35081 57412
rect 35115 57409 35127 57443
rect 35069 57403 35127 57409
rect 44910 57400 44916 57452
rect 44968 57440 44974 57452
rect 45005 57443 45063 57449
rect 45005 57440 45017 57443
rect 44968 57412 45017 57440
rect 44968 57400 44974 57412
rect 45005 57409 45017 57412
rect 45051 57409 45063 57443
rect 45005 57403 45063 57409
rect 54846 57400 54852 57452
rect 54904 57440 54910 57452
rect 55309 57443 55367 57449
rect 55309 57440 55321 57443
rect 54904 57412 55321 57440
rect 54904 57400 54910 57412
rect 55309 57409 55321 57412
rect 55355 57409 55367 57443
rect 55309 57403 55367 57409
rect 64782 57400 64788 57452
rect 64840 57440 64846 57452
rect 64877 57443 64935 57449
rect 64877 57440 64889 57443
rect 64840 57412 64889 57440
rect 64840 57400 64846 57412
rect 64877 57409 64889 57412
rect 64923 57409 64935 57443
rect 66990 57440 66996 57452
rect 66951 57412 66996 57440
rect 64877 57403 64935 57409
rect 66990 57400 66996 57412
rect 67048 57400 67054 57452
rect 67542 57400 67548 57452
rect 67600 57440 67606 57452
rect 67637 57443 67695 57449
rect 67637 57440 67649 57443
rect 67600 57412 67649 57440
rect 67600 57400 67606 57412
rect 67637 57409 67649 57412
rect 67683 57409 67695 57443
rect 67637 57403 67695 57409
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 68094 56828 68100 56840
rect 68055 56800 68100 56828
rect 68094 56788 68100 56800
rect 68152 56788 68158 56840
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 67634 55128 67640 55140
rect 67595 55100 67640 55128
rect 67634 55088 67640 55100
rect 67692 55088 67698 55140
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 67542 53932 67548 53984
rect 67600 53972 67606 53984
rect 67637 53975 67695 53981
rect 67637 53972 67649 53975
rect 67600 53944 67649 53972
rect 67600 53932 67606 53944
rect 67637 53941 67649 53944
rect 67683 53941 67695 53975
rect 67637 53935 67695 53941
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 68094 52476 68100 52488
rect 68055 52448 68100 52476
rect 68094 52436 68100 52448
rect 68152 52436 68158 52488
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 68094 51388 68100 51400
rect 68055 51360 68100 51388
rect 68094 51348 68100 51360
rect 68152 51348 68158 51400
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 67634 49756 67640 49768
rect 67595 49728 67640 49756
rect 67634 49716 67640 49728
rect 67692 49716 67698 49768
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 67634 48532 67640 48544
rect 67595 48504 67640 48532
rect 67634 48492 67640 48504
rect 67692 48492 67698 48544
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 68094 47036 68100 47048
rect 68055 47008 68100 47036
rect 68094 46996 68100 47008
rect 68152 46996 68158 47048
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 68094 45948 68100 45960
rect 68055 45920 68100 45948
rect 68094 45908 68100 45920
rect 68152 45908 68158 45960
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 67634 44248 67640 44260
rect 67595 44220 67640 44248
rect 67634 44208 67640 44220
rect 67692 44208 67698 44260
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 67634 43092 67640 43104
rect 67595 43064 67640 43092
rect 67634 43052 67640 43064
rect 67692 43052 67698 43104
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 68094 41596 68100 41608
rect 68055 41568 68100 41596
rect 68094 41556 68100 41568
rect 68152 41556 68158 41608
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 68094 40508 68100 40520
rect 68055 40480 68100 40508
rect 68094 40468 68100 40480
rect 68152 40468 68158 40520
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 67634 38808 67640 38820
rect 67595 38780 67640 38808
rect 67634 38768 67640 38780
rect 67692 38768 67698 38820
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 67634 37652 67640 37664
rect 67595 37624 67640 37652
rect 67634 37612 67640 37624
rect 67692 37612 67698 37664
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 68094 36156 68100 36168
rect 68055 36128 68100 36156
rect 68094 36116 68100 36128
rect 68152 36116 68158 36168
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 68094 35068 68100 35080
rect 68055 35040 68100 35068
rect 68094 35028 68100 35040
rect 68152 35028 68158 35080
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 67634 33368 67640 33380
rect 67595 33340 67640 33368
rect 67634 33328 67640 33340
rect 67692 33328 67698 33380
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 67634 32212 67640 32224
rect 67595 32184 67640 32212
rect 67634 32172 67640 32184
rect 67692 32172 67698 32224
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 15102 31696 15108 31748
rect 15160 31736 15166 31748
rect 15749 31739 15807 31745
rect 15749 31736 15761 31739
rect 15160 31708 15761 31736
rect 15160 31696 15166 31708
rect 15749 31705 15761 31708
rect 15795 31736 15807 31739
rect 20530 31736 20536 31748
rect 15795 31708 20536 31736
rect 15795 31705 15807 31708
rect 15749 31699 15807 31705
rect 20530 31696 20536 31708
rect 20588 31696 20594 31748
rect 17402 31628 17408 31680
rect 17460 31668 17466 31680
rect 17773 31671 17831 31677
rect 17773 31668 17785 31671
rect 17460 31640 17785 31668
rect 17460 31628 17466 31640
rect 17773 31637 17785 31640
rect 17819 31637 17831 31671
rect 17773 31631 17831 31637
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 7834 31356 7840 31408
rect 7892 31396 7898 31408
rect 8757 31399 8815 31405
rect 8757 31396 8769 31399
rect 7892 31368 8769 31396
rect 7892 31356 7898 31368
rect 8757 31365 8769 31368
rect 8803 31365 8815 31399
rect 8757 31359 8815 31365
rect 12437 31399 12495 31405
rect 12437 31365 12449 31399
rect 12483 31396 12495 31399
rect 15013 31399 15071 31405
rect 12483 31368 13032 31396
rect 12483 31365 12495 31368
rect 12437 31359 12495 31365
rect 8386 31288 8392 31340
rect 8444 31328 8450 31340
rect 8573 31331 8631 31337
rect 8573 31328 8585 31331
rect 8444 31300 8585 31328
rect 8444 31288 8450 31300
rect 8573 31297 8585 31300
rect 8619 31328 8631 31331
rect 12066 31328 12072 31340
rect 8619 31300 12072 31328
rect 8619 31297 8631 31300
rect 8573 31291 8631 31297
rect 12066 31288 12072 31300
rect 12124 31288 12130 31340
rect 12253 31331 12311 31337
rect 12253 31297 12265 31331
rect 12299 31328 12311 31331
rect 12618 31328 12624 31340
rect 12299 31300 12624 31328
rect 12299 31297 12311 31300
rect 12253 31291 12311 31297
rect 12618 31288 12624 31300
rect 12676 31288 12682 31340
rect 12894 31328 12900 31340
rect 12855 31300 12900 31328
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 13004 31331 13032 31368
rect 15013 31365 15025 31399
rect 15059 31396 15071 31399
rect 15286 31396 15292 31408
rect 15059 31368 15292 31396
rect 15059 31365 15071 31368
rect 15013 31359 15071 31365
rect 15286 31356 15292 31368
rect 15344 31356 15350 31408
rect 17770 31396 17776 31408
rect 17052 31368 17776 31396
rect 13060 31334 13118 31340
rect 13060 31331 13072 31334
rect 13004 31303 13072 31331
rect 13060 31300 13072 31303
rect 13106 31300 13118 31334
rect 13060 31294 13118 31300
rect 13170 31288 13176 31340
rect 13228 31328 13234 31340
rect 13311 31331 13369 31337
rect 13228 31300 13273 31328
rect 13228 31288 13234 31300
rect 13311 31297 13323 31331
rect 13357 31328 13369 31331
rect 15194 31328 15200 31340
rect 13357 31300 14136 31328
rect 15155 31300 15200 31328
rect 13357 31297 13369 31300
rect 13311 31291 13369 31297
rect 14108 31201 14136 31300
rect 15194 31288 15200 31300
rect 15252 31288 15258 31340
rect 15933 31331 15991 31337
rect 15933 31297 15945 31331
rect 15979 31328 15991 31331
rect 16666 31328 16672 31340
rect 15979 31300 16672 31328
rect 15979 31297 15991 31300
rect 15933 31291 15991 31297
rect 16666 31288 16672 31300
rect 16724 31328 16730 31340
rect 17052 31337 17080 31368
rect 17770 31356 17776 31368
rect 17828 31356 17834 31408
rect 21821 31399 21879 31405
rect 21821 31396 21833 31399
rect 20548 31368 21833 31396
rect 20548 31340 20576 31368
rect 21821 31365 21833 31368
rect 21867 31396 21879 31399
rect 22738 31396 22744 31408
rect 21867 31368 22744 31396
rect 21867 31365 21879 31368
rect 21821 31359 21879 31365
rect 22738 31356 22744 31368
rect 22796 31356 22802 31408
rect 23014 31356 23020 31408
rect 23072 31396 23078 31408
rect 23477 31399 23535 31405
rect 23477 31396 23489 31399
rect 23072 31368 23489 31396
rect 23072 31356 23078 31368
rect 23477 31365 23489 31368
rect 23523 31365 23535 31399
rect 23477 31359 23535 31365
rect 23661 31399 23719 31405
rect 23661 31365 23673 31399
rect 23707 31396 23719 31399
rect 23707 31368 24348 31396
rect 23707 31365 23719 31368
rect 23661 31359 23719 31365
rect 17037 31331 17095 31337
rect 17037 31328 17049 31331
rect 16724 31300 17049 31328
rect 16724 31288 16730 31300
rect 17037 31297 17049 31300
rect 17083 31297 17095 31331
rect 17218 31328 17224 31340
rect 17179 31300 17224 31328
rect 17037 31291 17095 31297
rect 17218 31288 17224 31300
rect 17276 31288 17282 31340
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31297 17371 31331
rect 17313 31291 17371 31297
rect 14093 31195 14151 31201
rect 14093 31161 14105 31195
rect 14139 31192 14151 31195
rect 15470 31192 15476 31204
rect 14139 31164 15476 31192
rect 14139 31161 14151 31164
rect 14093 31155 14151 31161
rect 15470 31152 15476 31164
rect 15528 31152 15534 31204
rect 16574 31152 16580 31204
rect 16632 31192 16638 31204
rect 17328 31192 17356 31291
rect 17402 31288 17408 31340
rect 17460 31328 17466 31340
rect 20530 31328 20536 31340
rect 17460 31300 17505 31328
rect 20491 31300 20536 31328
rect 17460 31288 17466 31300
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 20625 31331 20683 31337
rect 20625 31297 20637 31331
rect 20671 31297 20683 31331
rect 20625 31291 20683 31297
rect 20640 31260 20668 31291
rect 20714 31288 20720 31340
rect 20772 31328 20778 31340
rect 20772 31300 20817 31328
rect 20772 31288 20778 31300
rect 20898 31288 20904 31340
rect 20956 31328 20962 31340
rect 23290 31328 23296 31340
rect 20956 31300 21001 31328
rect 23251 31300 23296 31328
rect 20956 31288 20962 31300
rect 23290 31288 23296 31300
rect 23348 31288 23354 31340
rect 24026 31288 24032 31340
rect 24084 31328 24090 31340
rect 24320 31337 24348 31368
rect 24121 31331 24179 31337
rect 24121 31328 24133 31331
rect 24084 31300 24133 31328
rect 24084 31288 24090 31300
rect 24121 31297 24133 31300
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 24305 31331 24363 31337
rect 24305 31297 24317 31331
rect 24351 31297 24363 31331
rect 24305 31291 24363 31297
rect 24397 31331 24455 31337
rect 24397 31297 24409 31331
rect 24443 31297 24455 31331
rect 24397 31291 24455 31297
rect 22094 31260 22100 31272
rect 20640 31232 22100 31260
rect 22094 31220 22100 31232
rect 22152 31260 22158 31272
rect 23750 31260 23756 31272
rect 22152 31232 23756 31260
rect 22152 31220 22158 31232
rect 23750 31220 23756 31232
rect 23808 31260 23814 31272
rect 24412 31260 24440 31291
rect 24486 31288 24492 31340
rect 24544 31328 24550 31340
rect 24544 31300 24589 31328
rect 24544 31288 24550 31300
rect 23808 31232 24440 31260
rect 23808 31220 23814 31232
rect 16632 31164 17356 31192
rect 16632 31152 16638 31164
rect 17770 31152 17776 31204
rect 17828 31192 17834 31204
rect 18141 31195 18199 31201
rect 18141 31192 18153 31195
rect 17828 31164 18153 31192
rect 17828 31152 17834 31164
rect 18141 31161 18153 31164
rect 18187 31161 18199 31195
rect 18141 31155 18199 31161
rect 8941 31127 8999 31133
rect 8941 31093 8953 31127
rect 8987 31124 8999 31127
rect 9398 31124 9404 31136
rect 8987 31096 9404 31124
rect 8987 31093 8999 31096
rect 8941 31087 8999 31093
rect 9398 31084 9404 31096
rect 9456 31084 9462 31136
rect 13538 31124 13544 31136
rect 13499 31096 13544 31124
rect 13538 31084 13544 31096
rect 13596 31084 13602 31136
rect 15378 31124 15384 31136
rect 15339 31096 15384 31124
rect 15378 31084 15384 31096
rect 15436 31084 15442 31136
rect 17681 31127 17739 31133
rect 17681 31093 17693 31127
rect 17727 31124 17739 31127
rect 18046 31124 18052 31136
rect 17727 31096 18052 31124
rect 17727 31093 17739 31096
rect 17681 31087 17739 31093
rect 18046 31084 18052 31096
rect 18104 31084 18110 31136
rect 20254 31124 20260 31136
rect 20215 31096 20260 31124
rect 20254 31084 20260 31096
rect 20312 31084 20318 31136
rect 24765 31127 24823 31133
rect 24765 31093 24777 31127
rect 24811 31124 24823 31127
rect 26142 31124 26148 31136
rect 24811 31096 26148 31124
rect 24811 31093 24823 31096
rect 24765 31087 24823 31093
rect 26142 31084 26148 31096
rect 26200 31084 26206 31136
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 9306 30880 9312 30932
rect 9364 30920 9370 30932
rect 10321 30923 10379 30929
rect 10321 30920 10333 30923
rect 9364 30892 10333 30920
rect 9364 30880 9370 30892
rect 10321 30889 10333 30892
rect 10367 30920 10379 30923
rect 15102 30920 15108 30932
rect 10367 30892 15108 30920
rect 10367 30889 10379 30892
rect 10321 30883 10379 30889
rect 15102 30880 15108 30892
rect 15160 30880 15166 30932
rect 17218 30880 17224 30932
rect 17276 30920 17282 30932
rect 17497 30923 17555 30929
rect 17497 30920 17509 30923
rect 17276 30892 17509 30920
rect 17276 30880 17282 30892
rect 17497 30889 17509 30892
rect 17543 30889 17555 30923
rect 17497 30883 17555 30889
rect 20257 30923 20315 30929
rect 20257 30889 20269 30923
rect 20303 30920 20315 30923
rect 20714 30920 20720 30932
rect 20303 30892 20720 30920
rect 20303 30889 20315 30892
rect 20257 30883 20315 30889
rect 20714 30880 20720 30892
rect 20772 30880 20778 30932
rect 13262 30852 13268 30864
rect 8956 30824 9628 30852
rect 8386 30716 8392 30728
rect 8347 30688 8392 30716
rect 8386 30676 8392 30688
rect 8444 30676 8450 30728
rect 8202 30648 8208 30660
rect 8163 30620 8208 30648
rect 8202 30608 8208 30620
rect 8260 30608 8266 30660
rect 8021 30583 8079 30589
rect 8021 30549 8033 30583
rect 8067 30580 8079 30583
rect 8956 30580 8984 30824
rect 9306 30676 9312 30728
rect 9364 30725 9370 30728
rect 9364 30719 9413 30725
rect 9364 30685 9367 30719
rect 9401 30685 9413 30719
rect 9364 30679 9413 30685
rect 9493 30719 9551 30725
rect 9600 30722 9628 30824
rect 11717 30824 13268 30852
rect 9674 30744 9680 30796
rect 9732 30784 9738 30796
rect 11717 30784 11745 30824
rect 13262 30812 13268 30824
rect 13320 30812 13326 30864
rect 17402 30852 17408 30864
rect 15166 30824 17408 30852
rect 11882 30784 11888 30796
rect 9732 30756 11745 30784
rect 9732 30744 9738 30756
rect 9493 30685 9505 30719
rect 9539 30685 9551 30719
rect 9493 30679 9551 30685
rect 9590 30716 9648 30722
rect 9590 30682 9602 30716
rect 9636 30682 9648 30716
rect 9364 30676 9370 30679
rect 9508 30648 9536 30679
rect 9590 30676 9648 30682
rect 9766 30676 9772 30728
rect 9824 30716 9830 30728
rect 11717 30725 11745 30756
rect 11808 30756 11888 30784
rect 11808 30725 11836 30756
rect 11882 30744 11888 30756
rect 11940 30744 11946 30796
rect 15166 30784 15194 30824
rect 17402 30812 17408 30824
rect 17460 30812 17466 30864
rect 16574 30784 16580 30796
rect 12452 30756 15194 30784
rect 15304 30756 16580 30784
rect 11589 30719 11647 30725
rect 11589 30716 11601 30719
rect 9824 30688 9869 30716
rect 11532 30688 11601 30716
rect 9824 30676 9830 30688
rect 9674 30648 9680 30660
rect 9508 30620 9680 30648
rect 9674 30608 9680 30620
rect 9732 30608 9738 30660
rect 9122 30580 9128 30592
rect 8067 30552 8984 30580
rect 9083 30552 9128 30580
rect 8067 30549 8079 30552
rect 8021 30543 8079 30549
rect 9122 30540 9128 30552
rect 9180 30540 9186 30592
rect 11330 30580 11336 30592
rect 11291 30552 11336 30580
rect 11330 30540 11336 30552
rect 11388 30540 11394 30592
rect 11532 30580 11560 30688
rect 11589 30685 11601 30688
rect 11635 30685 11647 30719
rect 11589 30679 11647 30685
rect 11701 30719 11759 30725
rect 11701 30685 11713 30719
rect 11747 30685 11759 30719
rect 11701 30679 11759 30685
rect 11798 30719 11856 30725
rect 11798 30685 11810 30719
rect 11844 30685 11856 30719
rect 11974 30716 11980 30728
rect 11935 30688 11980 30716
rect 11798 30679 11856 30685
rect 11974 30676 11980 30688
rect 12032 30676 12038 30728
rect 12452 30589 12480 30756
rect 15102 30676 15108 30728
rect 15160 30716 15166 30728
rect 15304 30725 15332 30756
rect 15197 30719 15255 30725
rect 15197 30716 15209 30719
rect 15160 30688 15209 30716
rect 15160 30676 15166 30688
rect 15197 30685 15209 30688
rect 15243 30685 15255 30719
rect 15197 30679 15255 30685
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30685 15347 30719
rect 15289 30679 15347 30685
rect 15378 30676 15384 30728
rect 15436 30716 15442 30728
rect 15565 30719 15623 30725
rect 15436 30688 15481 30716
rect 15436 30676 15442 30688
rect 15565 30685 15577 30719
rect 15611 30716 15623 30719
rect 16025 30719 16083 30725
rect 16025 30716 16037 30719
rect 15611 30688 16037 30716
rect 15611 30685 15623 30688
rect 15565 30679 15623 30685
rect 16025 30685 16037 30688
rect 16071 30685 16083 30719
rect 16206 30716 16212 30728
rect 16167 30688 16212 30716
rect 16025 30679 16083 30685
rect 16040 30648 16068 30679
rect 16206 30676 16212 30688
rect 16264 30676 16270 30728
rect 16316 30725 16344 30756
rect 16574 30744 16580 30756
rect 16632 30744 16638 30796
rect 16669 30787 16727 30793
rect 16669 30753 16681 30787
rect 16715 30784 16727 30787
rect 18414 30784 18420 30796
rect 16715 30756 18420 30784
rect 16715 30753 16727 30756
rect 16669 30747 16727 30753
rect 18414 30744 18420 30756
rect 18472 30744 18478 30796
rect 16301 30719 16359 30725
rect 16301 30685 16313 30719
rect 16347 30685 16359 30719
rect 16301 30679 16359 30685
rect 16390 30676 16396 30728
rect 16448 30716 16454 30728
rect 20441 30719 20499 30725
rect 16448 30688 18092 30716
rect 16448 30676 16454 30688
rect 16666 30648 16672 30660
rect 16040 30620 16672 30648
rect 16666 30608 16672 30620
rect 16724 30608 16730 30660
rect 17129 30651 17187 30657
rect 17129 30617 17141 30651
rect 17175 30617 17187 30651
rect 17129 30611 17187 30617
rect 12437 30583 12495 30589
rect 12437 30580 12449 30583
rect 11532 30552 12449 30580
rect 12437 30549 12449 30552
rect 12483 30549 12495 30583
rect 14918 30580 14924 30592
rect 14879 30552 14924 30580
rect 12437 30543 12495 30549
rect 14918 30540 14924 30552
rect 14976 30540 14982 30592
rect 15286 30540 15292 30592
rect 15344 30580 15350 30592
rect 17144 30580 17172 30611
rect 17218 30608 17224 30660
rect 17276 30648 17282 30660
rect 17313 30651 17371 30657
rect 17313 30648 17325 30651
rect 17276 30620 17325 30648
rect 17276 30608 17282 30620
rect 17313 30617 17325 30620
rect 17359 30617 17371 30651
rect 17313 30611 17371 30617
rect 18064 30589 18092 30688
rect 20441 30685 20453 30719
rect 20487 30716 20499 30719
rect 20714 30716 20720 30728
rect 20487 30688 20720 30716
rect 20487 30685 20499 30688
rect 20441 30679 20499 30685
rect 20714 30676 20720 30688
rect 20772 30676 20778 30728
rect 68094 30716 68100 30728
rect 68055 30688 68100 30716
rect 68094 30676 68100 30688
rect 68152 30676 68158 30728
rect 20622 30648 20628 30660
rect 20583 30620 20628 30648
rect 20622 30608 20628 30620
rect 20680 30608 20686 30660
rect 15344 30552 17172 30580
rect 18049 30583 18107 30589
rect 15344 30540 15350 30552
rect 18049 30549 18061 30583
rect 18095 30580 18107 30583
rect 18322 30580 18328 30592
rect 18095 30552 18328 30580
rect 18095 30549 18107 30552
rect 18049 30543 18107 30549
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 24394 30580 24400 30592
rect 24355 30552 24400 30580
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 5813 30379 5871 30385
rect 5813 30345 5825 30379
rect 5859 30376 5871 30379
rect 7834 30376 7840 30388
rect 5859 30348 7840 30376
rect 5859 30345 5871 30348
rect 5813 30339 5871 30345
rect 7834 30336 7840 30348
rect 7892 30336 7898 30388
rect 11882 30376 11888 30388
rect 11843 30348 11888 30376
rect 11882 30336 11888 30348
rect 11940 30336 11946 30388
rect 15657 30379 15715 30385
rect 15657 30345 15669 30379
rect 15703 30376 15715 30379
rect 16206 30376 16212 30388
rect 15703 30348 16212 30376
rect 15703 30345 15715 30348
rect 15657 30339 15715 30345
rect 16206 30336 16212 30348
rect 16264 30336 16270 30388
rect 7092 30311 7150 30317
rect 4448 30280 6868 30308
rect 3786 30200 3792 30252
rect 3844 30240 3850 30252
rect 4448 30249 4476 30280
rect 4433 30243 4491 30249
rect 4433 30240 4445 30243
rect 3844 30212 4445 30240
rect 3844 30200 3850 30212
rect 4433 30209 4445 30212
rect 4479 30209 4491 30243
rect 4433 30203 4491 30209
rect 4700 30243 4758 30249
rect 4700 30209 4712 30243
rect 4746 30240 4758 30243
rect 4746 30212 6684 30240
rect 4746 30209 4758 30212
rect 4700 30203 4758 30209
rect 6656 30036 6684 30212
rect 6840 30184 6868 30280
rect 7092 30277 7104 30311
rect 7138 30308 7150 30311
rect 9122 30308 9128 30320
rect 7138 30280 9128 30308
rect 7138 30277 7150 30280
rect 7092 30271 7150 30277
rect 9122 30268 9128 30280
rect 9180 30268 9186 30320
rect 9674 30308 9680 30320
rect 9321 30280 9680 30308
rect 9321 30252 9349 30280
rect 9674 30268 9680 30280
rect 9732 30268 9738 30320
rect 10410 30268 10416 30320
rect 10468 30308 10474 30320
rect 11701 30311 11759 30317
rect 11701 30308 11713 30311
rect 10468 30280 11713 30308
rect 10468 30268 10474 30280
rect 11701 30277 11713 30280
rect 11747 30277 11759 30311
rect 11701 30271 11759 30277
rect 13538 30268 13544 30320
rect 13596 30308 13602 30320
rect 13734 30311 13792 30317
rect 13734 30308 13746 30311
rect 13596 30280 13746 30308
rect 13596 30268 13602 30280
rect 13734 30277 13746 30280
rect 13780 30277 13792 30311
rect 15473 30311 15531 30317
rect 15473 30308 15485 30311
rect 13734 30271 13792 30277
rect 15120 30280 15485 30308
rect 9217 30243 9275 30249
rect 9217 30209 9229 30243
rect 9263 30209 9275 30243
rect 9217 30203 9275 30209
rect 9306 30246 9364 30252
rect 9306 30212 9318 30246
rect 9352 30212 9364 30246
rect 9306 30206 9364 30212
rect 6822 30172 6828 30184
rect 6783 30144 6828 30172
rect 6822 30132 6828 30144
rect 6880 30132 6886 30184
rect 8941 30107 8999 30113
rect 8941 30104 8953 30107
rect 7760 30076 8953 30104
rect 7760 30036 7788 30076
rect 8941 30073 8953 30076
rect 8987 30073 8999 30107
rect 9232 30104 9260 30203
rect 9398 30200 9404 30252
rect 9456 30240 9462 30252
rect 9585 30243 9643 30249
rect 9456 30212 9501 30240
rect 9456 30200 9462 30212
rect 9585 30209 9597 30243
rect 9631 30209 9643 30243
rect 9585 30203 9643 30209
rect 11517 30243 11575 30249
rect 11517 30209 11529 30243
rect 11563 30240 11575 30243
rect 12066 30240 12072 30252
rect 11563 30212 12072 30240
rect 11563 30209 11575 30212
rect 11517 30203 11575 30209
rect 9600 30172 9628 30203
rect 12066 30200 12072 30212
rect 12124 30200 12130 30252
rect 12434 30200 12440 30252
rect 12492 30240 12498 30252
rect 15120 30240 15148 30280
rect 15473 30277 15485 30280
rect 15519 30308 15531 30311
rect 17310 30308 17316 30320
rect 15519 30280 17316 30308
rect 15519 30277 15531 30280
rect 15473 30271 15531 30277
rect 17310 30268 17316 30280
rect 17368 30268 17374 30320
rect 18046 30268 18052 30320
rect 18104 30308 18110 30320
rect 18610 30311 18668 30317
rect 18610 30308 18622 30311
rect 18104 30280 18622 30308
rect 18104 30268 18110 30280
rect 18610 30277 18622 30280
rect 18656 30277 18668 30311
rect 18610 30271 18668 30277
rect 19604 30311 19662 30317
rect 19604 30277 19616 30311
rect 19650 30308 19662 30311
rect 20254 30308 20260 30320
rect 19650 30280 20260 30308
rect 19650 30277 19662 30280
rect 19604 30271 19662 30277
rect 20254 30268 20260 30280
rect 20312 30268 20318 30320
rect 23290 30268 23296 30320
rect 23348 30308 23354 30320
rect 23661 30311 23719 30317
rect 23661 30308 23673 30311
rect 23348 30280 23673 30308
rect 23348 30268 23354 30280
rect 23661 30277 23673 30280
rect 23707 30277 23719 30311
rect 23661 30271 23719 30277
rect 24946 30268 24952 30320
rect 25004 30308 25010 30320
rect 25004 30280 26464 30308
rect 25004 30268 25010 30280
rect 15286 30240 15292 30252
rect 12492 30212 15148 30240
rect 15247 30212 15292 30240
rect 12492 30200 12498 30212
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 18874 30240 18880 30252
rect 18835 30212 18880 30240
rect 18874 30200 18880 30212
rect 18932 30240 18938 30252
rect 19337 30243 19395 30249
rect 19337 30240 19349 30243
rect 18932 30212 19349 30240
rect 18932 30200 18938 30212
rect 19337 30209 19349 30212
rect 19383 30209 19395 30243
rect 19337 30203 19395 30209
rect 21910 30200 21916 30252
rect 21968 30240 21974 30252
rect 22077 30243 22135 30249
rect 22077 30240 22089 30243
rect 21968 30212 22089 30240
rect 21968 30200 21974 30212
rect 22077 30209 22089 30212
rect 22123 30209 22135 30243
rect 22077 30203 22135 30209
rect 23845 30243 23903 30249
rect 23845 30209 23857 30243
rect 23891 30240 23903 30243
rect 24486 30240 24492 30252
rect 23891 30212 24492 30240
rect 23891 30209 23903 30212
rect 23845 30203 23903 30209
rect 24486 30200 24492 30212
rect 24544 30200 24550 30252
rect 26142 30200 26148 30252
rect 26200 30249 26206 30252
rect 26436 30249 26464 30280
rect 26200 30240 26212 30249
rect 26421 30243 26479 30249
rect 26200 30212 26245 30240
rect 26200 30203 26212 30212
rect 26421 30209 26433 30243
rect 26467 30240 26479 30243
rect 27614 30240 27620 30252
rect 26467 30212 27620 30240
rect 26467 30209 26479 30212
rect 26421 30203 26479 30209
rect 26200 30200 26206 30203
rect 27614 30200 27620 30212
rect 27672 30240 27678 30252
rect 28169 30243 28227 30249
rect 28169 30240 28181 30243
rect 27672 30212 28181 30240
rect 27672 30200 27678 30212
rect 28169 30209 28181 30212
rect 28215 30209 28227 30243
rect 28169 30203 28227 30209
rect 28258 30200 28264 30252
rect 28316 30240 28322 30252
rect 28425 30243 28483 30249
rect 28425 30240 28437 30243
rect 28316 30212 28437 30240
rect 28316 30200 28322 30212
rect 28425 30209 28437 30212
rect 28471 30209 28483 30243
rect 28425 30203 28483 30209
rect 12894 30172 12900 30184
rect 9600 30144 12900 30172
rect 12894 30132 12900 30144
rect 12952 30132 12958 30184
rect 13998 30172 14004 30184
rect 13959 30144 14004 30172
rect 13998 30132 14004 30144
rect 14056 30132 14062 30184
rect 21818 30172 21824 30184
rect 21779 30144 21824 30172
rect 21818 30132 21824 30144
rect 21876 30132 21882 30184
rect 10137 30107 10195 30113
rect 10137 30104 10149 30107
rect 9232 30076 10149 30104
rect 8941 30067 8999 30073
rect 10137 30073 10149 30076
rect 10183 30104 10195 30107
rect 17037 30107 17095 30113
rect 10183 30076 13124 30104
rect 10183 30073 10195 30076
rect 10137 30067 10195 30073
rect 8202 30036 8208 30048
rect 6656 30008 7788 30036
rect 8163 30008 8208 30036
rect 8202 29996 8208 30008
rect 8260 29996 8266 30048
rect 12618 30036 12624 30048
rect 12579 30008 12624 30036
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 13096 30036 13124 30076
rect 17037 30073 17049 30107
rect 17083 30104 17095 30107
rect 17770 30104 17776 30116
rect 17083 30076 17776 30104
rect 17083 30073 17095 30076
rect 17037 30067 17095 30073
rect 17770 30064 17776 30076
rect 17828 30064 17834 30116
rect 23014 30064 23020 30116
rect 23072 30104 23078 30116
rect 25041 30107 25099 30113
rect 25041 30104 25053 30107
rect 23072 30076 25053 30104
rect 23072 30064 23078 30076
rect 25041 30073 25053 30076
rect 25087 30073 25099 30107
rect 25041 30067 25099 30073
rect 16390 30036 16396 30048
rect 13096 30008 16396 30036
rect 16390 29996 16396 30008
rect 16448 29996 16454 30048
rect 17126 29996 17132 30048
rect 17184 30036 17190 30048
rect 17497 30039 17555 30045
rect 17497 30036 17509 30039
rect 17184 30008 17509 30036
rect 17184 29996 17190 30008
rect 17497 30005 17509 30008
rect 17543 30005 17555 30039
rect 20714 30036 20720 30048
rect 20675 30008 20720 30036
rect 17497 29999 17555 30005
rect 20714 29996 20720 30008
rect 20772 29996 20778 30048
rect 22462 29996 22468 30048
rect 22520 30036 22526 30048
rect 23106 30036 23112 30048
rect 22520 30008 23112 30036
rect 22520 29996 22526 30008
rect 23106 29996 23112 30008
rect 23164 30036 23170 30048
rect 23201 30039 23259 30045
rect 23201 30036 23213 30039
rect 23164 30008 23213 30036
rect 23164 29996 23170 30008
rect 23201 30005 23213 30008
rect 23247 30005 23259 30039
rect 23201 29999 23259 30005
rect 23934 29996 23940 30048
rect 23992 30036 23998 30048
rect 24029 30039 24087 30045
rect 24029 30036 24041 30039
rect 23992 30008 24041 30036
rect 23992 29996 23998 30008
rect 24029 30005 24041 30008
rect 24075 30005 24087 30039
rect 24029 29999 24087 30005
rect 29270 29996 29276 30048
rect 29328 30036 29334 30048
rect 29549 30039 29607 30045
rect 29549 30036 29561 30039
rect 29328 30008 29561 30036
rect 29328 29996 29334 30008
rect 29549 30005 29561 30008
rect 29595 30005 29607 30039
rect 29549 29999 29607 30005
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 10134 29792 10140 29844
rect 10192 29832 10198 29844
rect 10410 29832 10416 29844
rect 10192 29804 10416 29832
rect 10192 29792 10198 29804
rect 10410 29792 10416 29804
rect 10468 29792 10474 29844
rect 11974 29792 11980 29844
rect 12032 29832 12038 29844
rect 16758 29832 16764 29844
rect 12032 29804 16764 29832
rect 12032 29792 12038 29804
rect 16758 29792 16764 29804
rect 16816 29792 16822 29844
rect 17310 29832 17316 29844
rect 17271 29804 17316 29832
rect 17310 29792 17316 29804
rect 17368 29792 17374 29844
rect 18322 29792 18328 29844
rect 18380 29832 18386 29844
rect 20717 29835 20775 29841
rect 20717 29832 20729 29835
rect 18380 29804 20729 29832
rect 18380 29792 18386 29804
rect 20717 29801 20729 29804
rect 20763 29832 20775 29835
rect 21542 29832 21548 29844
rect 20763 29804 21548 29832
rect 20763 29801 20775 29804
rect 20717 29795 20775 29801
rect 21542 29792 21548 29804
rect 21600 29792 21606 29844
rect 21821 29835 21879 29841
rect 21821 29801 21833 29835
rect 21867 29832 21879 29835
rect 21910 29832 21916 29844
rect 21867 29804 21916 29832
rect 21867 29801 21879 29804
rect 21821 29795 21879 29801
rect 21910 29792 21916 29804
rect 21968 29792 21974 29844
rect 23750 29764 23756 29776
rect 21284 29736 21608 29764
rect 3786 29696 3792 29708
rect 3747 29668 3792 29696
rect 3786 29656 3792 29668
rect 3844 29656 3850 29708
rect 13998 29696 14004 29708
rect 12406 29668 14004 29696
rect 10502 29588 10508 29640
rect 10560 29628 10566 29640
rect 11793 29631 11851 29637
rect 11793 29628 11805 29631
rect 10560 29600 11805 29628
rect 10560 29588 10566 29600
rect 11793 29597 11805 29600
rect 11839 29628 11851 29631
rect 12406 29628 12434 29668
rect 13998 29656 14004 29668
rect 14056 29656 14062 29708
rect 11839 29600 12434 29628
rect 12529 29631 12587 29637
rect 11839 29597 11851 29600
rect 11793 29591 11851 29597
rect 12529 29597 12541 29631
rect 12575 29597 12587 29631
rect 12529 29591 12587 29597
rect 12621 29631 12679 29637
rect 12621 29597 12633 29631
rect 12667 29597 12679 29631
rect 12621 29591 12679 29597
rect 3326 29520 3332 29572
rect 3384 29560 3390 29572
rect 4034 29563 4092 29569
rect 4034 29560 4046 29563
rect 3384 29532 4046 29560
rect 3384 29520 3390 29532
rect 4034 29529 4046 29532
rect 4080 29529 4092 29563
rect 4034 29523 4092 29529
rect 11330 29520 11336 29572
rect 11388 29560 11394 29572
rect 11526 29563 11584 29569
rect 11526 29560 11538 29563
rect 11388 29532 11538 29560
rect 11388 29520 11394 29532
rect 11526 29529 11538 29532
rect 11572 29529 11584 29563
rect 11526 29523 11584 29529
rect 5166 29492 5172 29504
rect 5127 29464 5172 29492
rect 5166 29452 5172 29464
rect 5224 29452 5230 29504
rect 11054 29452 11060 29504
rect 11112 29492 11118 29504
rect 12253 29495 12311 29501
rect 12253 29492 12265 29495
rect 11112 29464 12265 29492
rect 11112 29452 11118 29464
rect 12253 29461 12265 29464
rect 12299 29461 12311 29495
rect 12544 29492 12572 29591
rect 12636 29560 12664 29591
rect 12710 29588 12716 29640
rect 12768 29628 12774 29640
rect 12768 29600 12813 29628
rect 12768 29588 12774 29600
rect 12894 29588 12900 29640
rect 12952 29628 12958 29640
rect 16577 29631 16635 29637
rect 12952 29600 12997 29628
rect 12952 29588 12958 29600
rect 16577 29597 16589 29631
rect 16623 29628 16635 29631
rect 18046 29628 18052 29640
rect 16623 29600 18052 29628
rect 16623 29597 16635 29600
rect 16577 29591 16635 29597
rect 18046 29588 18052 29600
rect 18104 29628 18110 29640
rect 18693 29631 18751 29637
rect 18693 29628 18705 29631
rect 18104 29600 18705 29628
rect 18104 29588 18110 29600
rect 18693 29597 18705 29600
rect 18739 29628 18751 29631
rect 18874 29628 18880 29640
rect 18739 29600 18880 29628
rect 18739 29597 18751 29600
rect 18693 29591 18751 29597
rect 18874 29588 18880 29600
rect 18932 29588 18938 29640
rect 20898 29588 20904 29640
rect 20956 29628 20962 29640
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 20956 29600 21189 29628
rect 20956 29588 20962 29600
rect 21177 29597 21189 29600
rect 21223 29597 21235 29631
rect 21284 29628 21312 29736
rect 21580 29696 21608 29736
rect 23676 29736 23756 29764
rect 22281 29699 22339 29705
rect 22281 29696 22293 29699
rect 21580 29668 22293 29696
rect 22281 29665 22293 29668
rect 22327 29665 22339 29699
rect 23676 29696 23704 29736
rect 23750 29724 23756 29736
rect 23808 29724 23814 29776
rect 22281 29659 22339 29665
rect 23584 29668 23704 29696
rect 21340 29631 21398 29637
rect 21340 29628 21352 29631
rect 21284 29600 21352 29628
rect 21177 29591 21235 29597
rect 21340 29597 21352 29600
rect 21386 29597 21398 29631
rect 21340 29591 21398 29597
rect 21440 29631 21498 29637
rect 21440 29597 21452 29631
rect 21486 29597 21498 29631
rect 21440 29591 21498 29597
rect 13262 29560 13268 29572
rect 12636 29532 13268 29560
rect 13262 29520 13268 29532
rect 13320 29520 13326 29572
rect 13449 29563 13507 29569
rect 13449 29529 13461 29563
rect 13495 29560 13507 29563
rect 13495 29532 16160 29560
rect 13495 29529 13507 29532
rect 13449 29523 13507 29529
rect 13464 29492 13492 29523
rect 12544 29464 13492 29492
rect 15197 29495 15255 29501
rect 12253 29455 12311 29461
rect 15197 29461 15209 29495
rect 15243 29492 15255 29495
rect 15562 29492 15568 29504
rect 15243 29464 15568 29492
rect 15243 29461 15255 29464
rect 15197 29455 15255 29461
rect 15562 29452 15568 29464
rect 15620 29452 15626 29504
rect 16132 29492 16160 29532
rect 16206 29520 16212 29572
rect 16264 29560 16270 29572
rect 16310 29563 16368 29569
rect 16310 29560 16322 29563
rect 16264 29532 16322 29560
rect 16264 29520 16270 29532
rect 16310 29529 16322 29532
rect 16356 29529 16368 29563
rect 16310 29523 16368 29529
rect 18414 29520 18420 29572
rect 18472 29569 18478 29572
rect 18472 29560 18484 29569
rect 21468 29560 21496 29591
rect 21542 29588 21548 29640
rect 21600 29628 21606 29640
rect 22462 29628 22468 29640
rect 21600 29600 21645 29628
rect 22423 29600 22468 29628
rect 21600 29588 21606 29600
rect 22462 29588 22468 29600
rect 22520 29588 22526 29640
rect 22646 29628 22652 29640
rect 22559 29600 22652 29628
rect 22646 29588 22652 29600
rect 22704 29628 22710 29640
rect 23290 29628 23296 29640
rect 22704 29600 23296 29628
rect 22704 29588 22710 29600
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 23477 29631 23535 29637
rect 23584 29631 23612 29668
rect 23682 29631 23740 29637
rect 23477 29597 23489 29631
rect 23523 29597 23535 29631
rect 23477 29591 23535 29597
rect 23582 29625 23640 29631
rect 23582 29591 23594 29625
rect 23628 29591 23640 29625
rect 23682 29597 23694 29631
rect 23728 29628 23740 29631
rect 23845 29631 23903 29637
rect 23728 29600 23796 29628
rect 23728 29597 23740 29600
rect 23682 29591 23740 29597
rect 22094 29560 22100 29572
rect 18472 29532 18517 29560
rect 21468 29532 22100 29560
rect 18472 29523 18484 29532
rect 18472 29520 18478 29523
rect 22094 29520 22100 29532
rect 22152 29520 22158 29572
rect 23492 29560 23520 29591
rect 23582 29585 23640 29591
rect 23124 29532 23520 29560
rect 23768 29560 23796 29600
rect 23845 29597 23857 29631
rect 23891 29628 23903 29631
rect 24026 29628 24032 29640
rect 23891 29600 24032 29628
rect 23891 29597 23903 29600
rect 23845 29591 23903 29597
rect 24026 29588 24032 29600
rect 24084 29588 24090 29640
rect 24946 29628 24952 29640
rect 24907 29600 24952 29628
rect 24946 29588 24952 29600
rect 25004 29588 25010 29640
rect 27614 29588 27620 29640
rect 27672 29628 27678 29640
rect 28169 29631 28227 29637
rect 28169 29628 28181 29631
rect 27672 29600 28181 29628
rect 27672 29588 27678 29600
rect 28169 29597 28181 29600
rect 28215 29597 28227 29631
rect 68094 29628 68100 29640
rect 68055 29600 68100 29628
rect 28169 29591 28227 29597
rect 68094 29588 68100 29600
rect 68152 29588 68158 29640
rect 23934 29560 23940 29572
rect 23768 29532 23940 29560
rect 16666 29492 16672 29504
rect 16132 29464 16672 29492
rect 16666 29452 16672 29464
rect 16724 29492 16730 29504
rect 17586 29492 17592 29504
rect 16724 29464 17592 29492
rect 16724 29452 16730 29464
rect 17586 29452 17592 29464
rect 17644 29492 17650 29504
rect 23124 29492 23152 29532
rect 17644 29464 23152 29492
rect 23201 29495 23259 29501
rect 17644 29452 17650 29464
rect 23201 29461 23213 29495
rect 23247 29492 23259 29495
rect 23290 29492 23296 29504
rect 23247 29464 23296 29492
rect 23247 29461 23259 29464
rect 23201 29455 23259 29461
rect 23290 29452 23296 29464
rect 23348 29452 23354 29504
rect 23492 29492 23520 29532
rect 23934 29520 23940 29532
rect 23992 29520 23998 29572
rect 25222 29569 25228 29572
rect 25216 29523 25228 29569
rect 25280 29560 25286 29572
rect 25280 29532 25316 29560
rect 25222 29520 25228 29523
rect 25280 29520 25286 29532
rect 25590 29520 25596 29572
rect 25648 29560 25654 29572
rect 25648 29532 26832 29560
rect 25648 29520 25654 29532
rect 24397 29495 24455 29501
rect 24397 29492 24409 29495
rect 23492 29464 24409 29492
rect 24397 29461 24409 29464
rect 24443 29492 24455 29495
rect 25130 29492 25136 29504
rect 24443 29464 25136 29492
rect 24443 29461 24455 29464
rect 24397 29455 24455 29461
rect 25130 29452 25136 29464
rect 25188 29452 25194 29504
rect 25866 29452 25872 29504
rect 25924 29492 25930 29504
rect 26804 29501 26832 29532
rect 27798 29520 27804 29572
rect 27856 29560 27862 29572
rect 27902 29563 27960 29569
rect 27902 29560 27914 29563
rect 27856 29532 27914 29560
rect 27856 29520 27862 29532
rect 27902 29529 27914 29532
rect 27948 29529 27960 29563
rect 27902 29523 27960 29529
rect 26329 29495 26387 29501
rect 26329 29492 26341 29495
rect 25924 29464 26341 29492
rect 25924 29452 25930 29464
rect 26329 29461 26341 29464
rect 26375 29461 26387 29495
rect 26329 29455 26387 29461
rect 26789 29495 26847 29501
rect 26789 29461 26801 29495
rect 26835 29461 26847 29495
rect 26789 29455 26847 29461
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 6730 29248 6736 29300
rect 6788 29288 6794 29300
rect 7745 29291 7803 29297
rect 7745 29288 7757 29291
rect 6788 29260 7757 29288
rect 6788 29248 6794 29260
rect 7745 29257 7757 29260
rect 7791 29288 7803 29291
rect 12158 29288 12164 29300
rect 7791 29260 11928 29288
rect 12119 29260 12164 29288
rect 7791 29257 7803 29260
rect 7745 29251 7803 29257
rect 6822 29220 6828 29232
rect 6380 29192 6828 29220
rect 6380 29161 6408 29192
rect 6822 29180 6828 29192
rect 6880 29220 6886 29232
rect 11790 29220 11796 29232
rect 6880 29192 9536 29220
rect 11751 29192 11796 29220
rect 6880 29180 6886 29192
rect 6638 29161 6644 29164
rect 6365 29155 6423 29161
rect 6365 29121 6377 29155
rect 6411 29121 6423 29155
rect 6365 29115 6423 29121
rect 6632 29115 6644 29161
rect 6696 29152 6702 29164
rect 6696 29124 6732 29152
rect 6638 29112 6644 29115
rect 6696 29112 6702 29124
rect 9508 29025 9536 29192
rect 11790 29180 11796 29192
rect 11848 29180 11854 29232
rect 10781 29155 10839 29161
rect 10781 29121 10793 29155
rect 10827 29152 10839 29155
rect 11330 29152 11336 29164
rect 10827 29124 11336 29152
rect 10827 29121 10839 29124
rect 10781 29115 10839 29121
rect 11330 29112 11336 29124
rect 11388 29112 11394 29164
rect 11900 29161 11928 29260
rect 12158 29248 12164 29260
rect 12216 29248 12222 29300
rect 12710 29248 12716 29300
rect 12768 29288 12774 29300
rect 12989 29291 13047 29297
rect 12989 29288 13001 29291
rect 12768 29260 13001 29288
rect 12768 29248 12774 29260
rect 12989 29257 13001 29260
rect 13035 29257 13047 29291
rect 15013 29291 15071 29297
rect 15013 29288 15025 29291
rect 12989 29251 13047 29257
rect 13556 29260 15025 29288
rect 12250 29180 12256 29232
rect 12308 29220 12314 29232
rect 12805 29223 12863 29229
rect 12805 29220 12817 29223
rect 12308 29192 12817 29220
rect 12308 29180 12314 29192
rect 12805 29189 12817 29192
rect 12851 29189 12863 29223
rect 12805 29183 12863 29189
rect 11517 29155 11575 29161
rect 11517 29121 11529 29155
rect 11563 29121 11575 29155
rect 11517 29115 11575 29121
rect 11665 29155 11723 29161
rect 11665 29121 11677 29155
rect 11711 29152 11723 29155
rect 11885 29155 11943 29161
rect 11711 29124 11836 29152
rect 11711 29121 11723 29124
rect 11665 29115 11723 29121
rect 9582 29044 9588 29096
rect 9640 29084 9646 29096
rect 11532 29084 11560 29115
rect 9640 29056 11560 29084
rect 11808 29084 11836 29124
rect 11885 29121 11897 29155
rect 11931 29121 11943 29155
rect 11885 29115 11943 29121
rect 11974 29112 11980 29164
rect 12032 29161 12038 29164
rect 12032 29152 12040 29161
rect 12032 29124 12077 29152
rect 12032 29115 12040 29124
rect 12032 29112 12038 29115
rect 12158 29112 12164 29164
rect 12216 29152 12222 29164
rect 12621 29155 12679 29161
rect 12621 29152 12633 29155
rect 12216 29124 12633 29152
rect 12216 29112 12222 29124
rect 12621 29121 12633 29124
rect 12667 29121 12679 29155
rect 12621 29115 12679 29121
rect 13556 29084 13584 29260
rect 15013 29257 15025 29260
rect 15059 29288 15071 29291
rect 15194 29288 15200 29300
rect 15059 29260 15200 29288
rect 15059 29257 15071 29260
rect 15013 29251 15071 29257
rect 15194 29248 15200 29260
rect 15252 29248 15258 29300
rect 17586 29288 17592 29300
rect 17547 29260 17592 29288
rect 17586 29248 17592 29260
rect 17644 29248 17650 29300
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 21266 29288 21272 29300
rect 20956 29260 21272 29288
rect 20956 29248 20962 29260
rect 21266 29248 21272 29260
rect 21324 29288 21330 29300
rect 24026 29288 24032 29300
rect 21324 29260 24032 29288
rect 21324 29248 21330 29260
rect 24026 29248 24032 29260
rect 24084 29248 24090 29300
rect 13998 29220 14004 29232
rect 13648 29192 14004 29220
rect 13648 29161 13676 29192
rect 13998 29180 14004 29192
rect 14056 29180 14062 29232
rect 15286 29180 15292 29232
rect 15344 29220 15350 29232
rect 16669 29223 16727 29229
rect 16669 29220 16681 29223
rect 15344 29192 16681 29220
rect 15344 29180 15350 29192
rect 16669 29189 16681 29192
rect 16715 29189 16727 29223
rect 20622 29220 20628 29232
rect 20583 29192 20628 29220
rect 16669 29183 16727 29189
rect 20622 29180 20628 29192
rect 20680 29220 20686 29232
rect 20680 29192 21036 29220
rect 20680 29180 20686 29192
rect 13633 29155 13691 29161
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13633 29115 13691 29121
rect 13900 29155 13958 29161
rect 13900 29121 13912 29155
rect 13946 29152 13958 29155
rect 14918 29152 14924 29164
rect 13946 29124 14924 29152
rect 13946 29121 13958 29124
rect 13900 29115 13958 29121
rect 14918 29112 14924 29124
rect 14976 29112 14982 29164
rect 16853 29155 16911 29161
rect 16853 29121 16865 29155
rect 16899 29152 16911 29155
rect 17310 29152 17316 29164
rect 16899 29124 17316 29152
rect 16899 29121 16911 29124
rect 16853 29115 16911 29121
rect 17310 29112 17316 29124
rect 17368 29112 17374 29164
rect 20070 29112 20076 29164
rect 20128 29152 20134 29164
rect 20809 29155 20867 29161
rect 20809 29152 20821 29155
rect 20128 29124 20821 29152
rect 20128 29112 20134 29124
rect 20809 29121 20821 29124
rect 20855 29121 20867 29155
rect 21008 29152 21036 29192
rect 21082 29180 21088 29232
rect 21140 29220 21146 29232
rect 21818 29220 21824 29232
rect 21140 29192 21824 29220
rect 21140 29180 21146 29192
rect 21818 29180 21824 29192
rect 21876 29220 21882 29232
rect 24946 29220 24952 29232
rect 21876 29192 24952 29220
rect 21876 29180 21882 29192
rect 22646 29152 22652 29164
rect 21008 29124 22652 29152
rect 20809 29115 20867 29121
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 23216 29161 23244 29192
rect 24946 29180 24952 29192
rect 25004 29180 25010 29232
rect 28905 29223 28963 29229
rect 28905 29189 28917 29223
rect 28951 29220 28963 29223
rect 29270 29220 29276 29232
rect 28951 29192 29276 29220
rect 28951 29189 28963 29192
rect 28905 29183 28963 29189
rect 29270 29180 29276 29192
rect 29328 29180 29334 29232
rect 31726 29192 33548 29220
rect 23201 29155 23259 29161
rect 23201 29121 23213 29155
rect 23247 29121 23259 29155
rect 23201 29115 23259 29121
rect 23290 29112 23296 29164
rect 23348 29152 23354 29164
rect 23457 29155 23515 29161
rect 23457 29152 23469 29155
rect 23348 29124 23469 29152
rect 23348 29112 23354 29124
rect 23457 29121 23469 29124
rect 23503 29121 23515 29155
rect 29086 29152 29092 29164
rect 29047 29124 29092 29152
rect 23457 29115 23515 29121
rect 29086 29112 29092 29124
rect 29144 29112 29150 29164
rect 30834 29152 30840 29164
rect 30892 29161 30898 29164
rect 30804 29124 30840 29152
rect 30834 29112 30840 29124
rect 30892 29115 30904 29161
rect 31113 29155 31171 29161
rect 31113 29121 31125 29155
rect 31159 29152 31171 29155
rect 31726 29152 31754 29192
rect 33520 29164 33548 29192
rect 31159 29124 31754 29152
rect 31159 29121 31171 29124
rect 31113 29115 31171 29121
rect 30892 29112 30898 29115
rect 32490 29112 32496 29164
rect 32548 29152 32554 29164
rect 33238 29155 33296 29161
rect 33238 29152 33250 29155
rect 32548 29124 33250 29152
rect 32548 29112 32554 29124
rect 33238 29121 33250 29124
rect 33284 29121 33296 29155
rect 33502 29152 33508 29164
rect 33415 29124 33508 29152
rect 33238 29115 33296 29121
rect 33502 29112 33508 29124
rect 33560 29112 33566 29164
rect 11808 29056 13584 29084
rect 9640 29044 9646 29056
rect 9493 29019 9551 29025
rect 9493 28985 9505 29019
rect 9539 29016 9551 29019
rect 10502 29016 10508 29028
rect 9539 28988 10508 29016
rect 9539 28985 9551 28988
rect 9493 28979 9551 28985
rect 10502 28976 10508 28988
rect 10560 28976 10566 29028
rect 12250 29016 12256 29028
rect 10612 28988 12256 29016
rect 7282 28908 7288 28960
rect 7340 28948 7346 28960
rect 8205 28951 8263 28957
rect 8205 28948 8217 28951
rect 7340 28920 8217 28948
rect 7340 28908 7346 28920
rect 8205 28917 8217 28920
rect 8251 28917 8263 28951
rect 8205 28911 8263 28917
rect 9674 28908 9680 28960
rect 9732 28948 9738 28960
rect 10612 28948 10640 28988
rect 12250 28976 12256 28988
rect 12308 28976 12314 29028
rect 20254 28976 20260 29028
rect 20312 29016 20318 29028
rect 21913 29019 21971 29025
rect 21913 29016 21925 29019
rect 20312 28988 21925 29016
rect 20312 28976 20318 28988
rect 21913 28985 21925 28988
rect 21959 29016 21971 29019
rect 22186 29016 22192 29028
rect 21959 28988 22192 29016
rect 21959 28985 21971 28988
rect 21913 28979 21971 28985
rect 22186 28976 22192 28988
rect 22244 28976 22250 29028
rect 24486 28976 24492 29028
rect 24544 29016 24550 29028
rect 24581 29019 24639 29025
rect 24581 29016 24593 29019
rect 24544 28988 24593 29016
rect 24544 28976 24550 28988
rect 24581 28985 24593 28988
rect 24627 28985 24639 29019
rect 24581 28979 24639 28985
rect 26234 28976 26240 29028
rect 26292 29016 26298 29028
rect 27893 29019 27951 29025
rect 27893 29016 27905 29019
rect 26292 28988 27905 29016
rect 26292 28976 26298 28988
rect 27893 28985 27905 28988
rect 27939 28985 27951 29019
rect 27893 28979 27951 28985
rect 29733 29019 29791 29025
rect 29733 28985 29745 29019
rect 29779 29016 29791 29019
rect 29914 29016 29920 29028
rect 29779 28988 29920 29016
rect 29779 28985 29791 28988
rect 29733 28979 29791 28985
rect 29914 28976 29920 28988
rect 29972 28976 29978 29028
rect 9732 28920 10640 28948
rect 9732 28908 9738 28920
rect 11882 28908 11888 28960
rect 11940 28948 11946 28960
rect 15010 28948 15016 28960
rect 11940 28920 15016 28948
rect 11940 28908 11946 28920
rect 15010 28908 15016 28920
rect 15068 28908 15074 28960
rect 17037 28951 17095 28957
rect 17037 28917 17049 28951
rect 17083 28948 17095 28951
rect 17402 28948 17408 28960
rect 17083 28920 17408 28948
rect 17083 28917 17095 28920
rect 17037 28911 17095 28917
rect 17402 28908 17408 28920
rect 17460 28908 17466 28960
rect 20990 28948 20996 28960
rect 20951 28920 20996 28948
rect 20990 28908 20996 28920
rect 21048 28908 21054 28960
rect 21542 28908 21548 28960
rect 21600 28948 21606 28960
rect 25774 28948 25780 28960
rect 21600 28920 25780 28948
rect 21600 28908 21606 28920
rect 25774 28908 25780 28920
rect 25832 28908 25838 28960
rect 28718 28948 28724 28960
rect 28679 28920 28724 28948
rect 28718 28908 28724 28920
rect 28776 28908 28782 28960
rect 32122 28948 32128 28960
rect 32083 28920 32128 28948
rect 32122 28908 32128 28920
rect 32180 28908 32186 28960
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 6549 28747 6607 28753
rect 6549 28713 6561 28747
rect 6595 28744 6607 28747
rect 6638 28744 6644 28756
rect 6595 28716 6644 28744
rect 6595 28713 6607 28716
rect 6549 28707 6607 28713
rect 6638 28704 6644 28716
rect 6696 28704 6702 28756
rect 8389 28747 8447 28753
rect 6748 28716 7512 28744
rect 5166 28636 5172 28688
rect 5224 28676 5230 28688
rect 6748 28676 6776 28716
rect 5224 28648 6776 28676
rect 5224 28636 5230 28648
rect 7484 28608 7512 28716
rect 8389 28713 8401 28747
rect 8435 28744 8447 28747
rect 16206 28744 16212 28756
rect 8435 28716 12204 28744
rect 16167 28716 16212 28744
rect 8435 28713 8447 28716
rect 8389 28707 8447 28713
rect 8110 28636 8116 28688
rect 8168 28676 8174 28688
rect 9493 28679 9551 28685
rect 8168 28648 8248 28676
rect 8168 28636 8174 28648
rect 7484 28580 8156 28608
rect 3418 28500 3424 28552
rect 3476 28540 3482 28552
rect 4065 28543 4123 28549
rect 4065 28540 4077 28543
rect 3476 28512 4077 28540
rect 3476 28500 3482 28512
rect 4065 28509 4077 28512
rect 4111 28509 4123 28543
rect 4065 28503 4123 28509
rect 5350 28500 5356 28552
rect 5408 28540 5414 28552
rect 6825 28543 6883 28549
rect 6825 28540 6837 28543
rect 5408 28512 6837 28540
rect 5408 28500 5414 28512
rect 6825 28509 6837 28512
rect 6871 28509 6883 28543
rect 6825 28503 6883 28509
rect 6917 28543 6975 28549
rect 6917 28509 6929 28543
rect 6963 28509 6975 28543
rect 6917 28503 6975 28509
rect 1762 28432 1768 28484
rect 1820 28472 1826 28484
rect 1949 28475 2007 28481
rect 1949 28472 1961 28475
rect 1820 28444 1961 28472
rect 1820 28432 1826 28444
rect 1949 28441 1961 28444
rect 1995 28441 2007 28475
rect 1949 28435 2007 28441
rect 2133 28475 2191 28481
rect 2133 28441 2145 28475
rect 2179 28472 2191 28475
rect 2179 28444 2774 28472
rect 2179 28441 2191 28444
rect 2133 28435 2191 28441
rect 2222 28364 2228 28416
rect 2280 28404 2286 28416
rect 2317 28407 2375 28413
rect 2317 28404 2329 28407
rect 2280 28376 2329 28404
rect 2280 28364 2286 28376
rect 2317 28373 2329 28376
rect 2363 28373 2375 28407
rect 2746 28404 2774 28444
rect 3234 28432 3240 28484
rect 3292 28472 3298 28484
rect 4310 28475 4368 28481
rect 4310 28472 4322 28475
rect 3292 28444 4322 28472
rect 3292 28432 3298 28444
rect 4310 28441 4322 28444
rect 4356 28441 4368 28475
rect 4310 28435 4368 28441
rect 5166 28404 5172 28416
rect 2746 28376 5172 28404
rect 2317 28367 2375 28373
rect 5166 28364 5172 28376
rect 5224 28364 5230 28416
rect 5442 28404 5448 28416
rect 5403 28376 5448 28404
rect 5442 28364 5448 28376
rect 5500 28364 5506 28416
rect 6840 28404 6868 28503
rect 6932 28472 6960 28503
rect 7006 28500 7012 28552
rect 7064 28540 7070 28552
rect 7193 28543 7251 28549
rect 7064 28512 7109 28540
rect 7064 28500 7070 28512
rect 7193 28509 7205 28543
rect 7239 28540 7251 28543
rect 7282 28540 7288 28552
rect 7239 28512 7288 28540
rect 7239 28509 7251 28512
rect 7193 28503 7251 28509
rect 7282 28500 7288 28512
rect 7340 28500 7346 28552
rect 7834 28540 7840 28552
rect 7795 28512 7840 28540
rect 7834 28500 7840 28512
rect 7892 28500 7898 28552
rect 8128 28549 8156 28580
rect 8220 28549 8248 28648
rect 9493 28645 9505 28679
rect 9539 28676 9551 28679
rect 9674 28676 9680 28688
rect 9539 28648 9680 28676
rect 9539 28645 9551 28648
rect 9493 28639 9551 28645
rect 9674 28636 9680 28648
rect 9732 28636 9738 28688
rect 12176 28549 12204 28716
rect 16206 28704 16212 28716
rect 16264 28704 16270 28756
rect 22189 28747 22247 28753
rect 22189 28713 22201 28747
rect 22235 28744 22247 28747
rect 22646 28744 22652 28756
rect 22235 28716 22652 28744
rect 22235 28713 22247 28716
rect 22189 28707 22247 28713
rect 22646 28704 22652 28716
rect 22704 28704 22710 28756
rect 27525 28747 27583 28753
rect 27525 28713 27537 28747
rect 27571 28744 27583 28747
rect 27614 28744 27620 28756
rect 27571 28716 27620 28744
rect 27571 28713 27583 28716
rect 27525 28707 27583 28713
rect 27614 28704 27620 28716
rect 27672 28704 27678 28756
rect 28258 28744 28264 28756
rect 28219 28716 28264 28744
rect 28258 28704 28264 28716
rect 28316 28704 28322 28756
rect 30929 28747 30987 28753
rect 30929 28713 30941 28747
rect 30975 28744 30987 28747
rect 32490 28744 32496 28756
rect 30975 28716 32496 28744
rect 30975 28713 30987 28716
rect 30929 28707 30987 28713
rect 32490 28704 32496 28716
rect 32548 28704 32554 28756
rect 12434 28676 12440 28688
rect 12268 28648 12440 28676
rect 12268 28549 12296 28648
rect 12434 28636 12440 28648
rect 12492 28636 12498 28688
rect 14642 28636 14648 28688
rect 14700 28676 14706 28688
rect 17310 28676 17316 28688
rect 14700 28648 17316 28676
rect 14700 28636 14706 28648
rect 17310 28636 17316 28648
rect 17368 28636 17374 28688
rect 30650 28676 30656 28688
rect 30484 28648 30656 28676
rect 15749 28611 15807 28617
rect 15749 28577 15761 28611
rect 15795 28608 15807 28611
rect 21082 28608 21088 28620
rect 15795 28580 16712 28608
rect 21043 28580 21088 28608
rect 15795 28577 15807 28580
rect 15749 28571 15807 28577
rect 8113 28543 8171 28549
rect 8113 28509 8125 28543
rect 8159 28509 8171 28543
rect 8113 28503 8171 28509
rect 8205 28543 8263 28549
rect 8205 28509 8217 28543
rect 8251 28509 8263 28543
rect 10873 28543 10931 28549
rect 10873 28540 10885 28543
rect 8205 28503 8263 28509
rect 10520 28512 10885 28540
rect 10520 28484 10548 28512
rect 10873 28509 10885 28512
rect 10919 28509 10931 28543
rect 10873 28503 10931 28509
rect 12161 28543 12219 28549
rect 12161 28509 12173 28543
rect 12207 28509 12219 28543
rect 12161 28503 12219 28509
rect 12254 28543 12312 28549
rect 12254 28509 12266 28543
rect 12300 28509 12312 28543
rect 12391 28543 12449 28549
rect 12391 28540 12403 28543
rect 12254 28503 12312 28509
rect 12365 28509 12403 28540
rect 12437 28509 12449 28543
rect 12526 28540 12532 28552
rect 12487 28512 12532 28540
rect 12365 28503 12449 28509
rect 7374 28472 7380 28484
rect 6932 28444 7380 28472
rect 7374 28432 7380 28444
rect 7432 28432 7438 28484
rect 8021 28475 8079 28481
rect 8021 28441 8033 28475
rect 8067 28472 8079 28475
rect 9122 28472 9128 28484
rect 8067 28444 9128 28472
rect 8067 28441 8079 28444
rect 8021 28435 8079 28441
rect 9122 28432 9128 28444
rect 9180 28432 9186 28484
rect 10502 28432 10508 28484
rect 10560 28432 10566 28484
rect 10628 28475 10686 28481
rect 10628 28441 10640 28475
rect 10674 28472 10686 28475
rect 11054 28472 11060 28484
rect 10674 28444 11060 28472
rect 10674 28441 10686 28444
rect 10628 28435 10686 28441
rect 11054 28432 11060 28444
rect 11112 28432 11118 28484
rect 11790 28432 11796 28484
rect 11848 28472 11854 28484
rect 12365 28472 12393 28503
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 12710 28549 12716 28552
rect 12667 28543 12716 28549
rect 12667 28509 12679 28543
rect 12713 28509 12716 28543
rect 12667 28503 12716 28509
rect 12710 28500 12716 28503
rect 12768 28500 12774 28552
rect 15286 28500 15292 28552
rect 15344 28540 15350 28552
rect 15381 28543 15439 28549
rect 15381 28540 15393 28543
rect 15344 28512 15393 28540
rect 15344 28500 15350 28512
rect 15381 28509 15393 28512
rect 15427 28509 15439 28543
rect 15381 28503 15439 28509
rect 16439 28543 16497 28549
rect 16439 28509 16451 28543
rect 16485 28509 16497 28543
rect 16574 28540 16580 28552
rect 16535 28512 16580 28540
rect 16439 28503 16497 28509
rect 15562 28472 15568 28484
rect 11848 28444 12393 28472
rect 15523 28444 15568 28472
rect 11848 28432 11854 28444
rect 15562 28432 15568 28444
rect 15620 28432 15626 28484
rect 16454 28472 16482 28503
rect 16574 28500 16580 28512
rect 16632 28500 16638 28552
rect 16684 28549 16712 28580
rect 21082 28568 21088 28580
rect 21140 28568 21146 28620
rect 22370 28568 22376 28620
rect 22428 28608 22434 28620
rect 22738 28608 22744 28620
rect 22428 28580 22744 28608
rect 22428 28568 22434 28580
rect 22738 28568 22744 28580
rect 22796 28608 22802 28620
rect 22796 28580 28212 28608
rect 22796 28568 22802 28580
rect 16669 28543 16727 28549
rect 16669 28509 16681 28543
rect 16715 28509 16727 28543
rect 16669 28503 16727 28509
rect 16853 28543 16911 28549
rect 16853 28509 16865 28543
rect 16899 28540 16911 28543
rect 17954 28540 17960 28552
rect 16899 28512 17960 28540
rect 16899 28509 16911 28512
rect 16853 28503 16911 28509
rect 17954 28500 17960 28512
rect 18012 28500 18018 28552
rect 18046 28500 18052 28552
rect 18104 28540 18110 28552
rect 18693 28543 18751 28549
rect 18693 28540 18705 28543
rect 18104 28512 18705 28540
rect 18104 28500 18110 28512
rect 18693 28509 18705 28512
rect 18739 28509 18751 28543
rect 18693 28503 18751 28509
rect 21818 28500 21824 28552
rect 21876 28540 21882 28552
rect 23492 28549 23520 28580
rect 28184 28552 28212 28580
rect 22005 28543 22063 28549
rect 22005 28540 22017 28543
rect 21876 28512 22017 28540
rect 21876 28500 21882 28512
rect 22005 28509 22017 28512
rect 22051 28509 22063 28543
rect 22005 28503 22063 28509
rect 23477 28543 23535 28549
rect 23477 28509 23489 28543
rect 23523 28509 23535 28543
rect 23477 28503 23535 28509
rect 23582 28540 23640 28546
rect 23582 28506 23594 28540
rect 23628 28506 23640 28540
rect 23582 28500 23640 28506
rect 23682 28540 23740 28546
rect 23682 28506 23694 28540
rect 23728 28512 23796 28540
rect 23728 28506 23740 28512
rect 23682 28500 23740 28506
rect 16454 28444 16574 28472
rect 8938 28404 8944 28416
rect 6840 28376 8944 28404
rect 8938 28364 8944 28376
rect 8996 28364 9002 28416
rect 11330 28404 11336 28416
rect 11291 28376 11336 28404
rect 11330 28364 11336 28376
rect 11388 28364 11394 28416
rect 12802 28404 12808 28416
rect 12763 28376 12808 28404
rect 12802 28364 12808 28376
rect 12860 28364 12866 28416
rect 16546 28404 16574 28444
rect 17862 28432 17868 28484
rect 17920 28472 17926 28484
rect 18426 28475 18484 28481
rect 18426 28472 18438 28475
rect 17920 28444 18438 28472
rect 17920 28432 17926 28444
rect 18426 28441 18438 28444
rect 18472 28441 18484 28475
rect 18426 28435 18484 28441
rect 20622 28432 20628 28484
rect 20680 28472 20686 28484
rect 20818 28475 20876 28481
rect 20818 28472 20830 28475
rect 20680 28444 20830 28472
rect 20680 28432 20686 28444
rect 20818 28441 20830 28444
rect 20864 28441 20876 28475
rect 20818 28435 20876 28441
rect 16666 28404 16672 28416
rect 16546 28376 16672 28404
rect 16666 28364 16672 28376
rect 16724 28404 16730 28416
rect 16942 28404 16948 28416
rect 16724 28376 16948 28404
rect 16724 28364 16730 28376
rect 16942 28364 16948 28376
rect 17000 28364 17006 28416
rect 19705 28407 19763 28413
rect 19705 28373 19717 28407
rect 19751 28404 19763 28407
rect 20070 28404 20076 28416
rect 19751 28376 20076 28404
rect 19751 28373 19763 28376
rect 19705 28367 19763 28373
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 23198 28404 23204 28416
rect 23159 28376 23204 28404
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 23584 28404 23612 28500
rect 23768 28472 23796 28512
rect 23842 28500 23848 28552
rect 23900 28540 23906 28552
rect 23900 28512 23945 28540
rect 23900 28500 23906 28512
rect 28166 28500 28172 28552
rect 28224 28540 28230 28552
rect 28537 28543 28595 28549
rect 28537 28540 28549 28543
rect 28224 28512 28549 28540
rect 28224 28500 28230 28512
rect 28537 28509 28549 28512
rect 28583 28509 28595 28543
rect 28537 28503 28595 28509
rect 28629 28543 28687 28549
rect 28629 28509 28641 28543
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 24302 28472 24308 28484
rect 23768 28444 24308 28472
rect 24302 28432 24308 28444
rect 24360 28432 24366 28484
rect 24854 28432 24860 28484
rect 24912 28472 24918 28484
rect 25225 28475 25283 28481
rect 25225 28472 25237 28475
rect 24912 28444 25237 28472
rect 24912 28432 24918 28444
rect 25225 28441 25237 28444
rect 25271 28441 25283 28475
rect 25225 28435 25283 28441
rect 25409 28475 25467 28481
rect 25409 28441 25421 28475
rect 25455 28472 25467 28475
rect 25866 28472 25872 28484
rect 25455 28444 25872 28472
rect 25455 28441 25467 28444
rect 25409 28435 25467 28441
rect 25866 28432 25872 28444
rect 25924 28432 25930 28484
rect 26053 28475 26111 28481
rect 26053 28441 26065 28475
rect 26099 28472 26111 28475
rect 26234 28472 26240 28484
rect 26099 28444 26240 28472
rect 26099 28441 26111 28444
rect 26053 28435 26111 28441
rect 26234 28432 26240 28444
rect 26292 28432 26298 28484
rect 28644 28472 28672 28503
rect 28718 28500 28724 28552
rect 28776 28540 28782 28552
rect 28776 28512 28821 28540
rect 28776 28500 28782 28512
rect 28902 28500 28908 28552
rect 28960 28540 28966 28552
rect 30285 28543 30343 28549
rect 30285 28540 30297 28543
rect 28960 28512 30297 28540
rect 28960 28500 28966 28512
rect 30285 28509 30297 28512
rect 30331 28509 30343 28543
rect 30285 28503 30343 28509
rect 30374 28500 30380 28552
rect 30432 28500 30438 28552
rect 30484 28549 30512 28648
rect 30650 28636 30656 28648
rect 30708 28636 30714 28688
rect 30469 28543 30527 28549
rect 30469 28509 30481 28543
rect 30515 28509 30527 28543
rect 30469 28503 30527 28509
rect 30558 28500 30564 28552
rect 30616 28540 30622 28552
rect 30742 28549 30748 28552
rect 30699 28543 30748 28549
rect 30616 28512 30661 28540
rect 30616 28500 30622 28512
rect 30699 28509 30711 28543
rect 30745 28509 30748 28543
rect 30699 28503 30748 28509
rect 30742 28500 30748 28503
rect 30800 28500 30806 28552
rect 28994 28472 29000 28484
rect 28644 28444 29000 28472
rect 28994 28432 29000 28444
rect 29052 28472 29058 28484
rect 30392 28472 30420 28500
rect 29052 28444 30420 28472
rect 29052 28432 29058 28444
rect 23750 28404 23756 28416
rect 23584 28376 23756 28404
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 25593 28407 25651 28413
rect 25593 28373 25605 28407
rect 25639 28404 25651 28407
rect 25682 28404 25688 28416
rect 25639 28376 25688 28404
rect 25639 28373 25651 28376
rect 25593 28367 25651 28373
rect 25682 28364 25688 28376
rect 25740 28364 25746 28416
rect 27338 28364 27344 28416
rect 27396 28404 27402 28416
rect 29733 28407 29791 28413
rect 29733 28404 29745 28407
rect 27396 28376 29745 28404
rect 27396 28364 27402 28376
rect 29733 28373 29745 28376
rect 29779 28404 29791 28407
rect 30466 28404 30472 28416
rect 29779 28376 30472 28404
rect 29779 28373 29791 28376
rect 29733 28367 29791 28373
rect 30466 28364 30472 28376
rect 30524 28364 30530 28416
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 3234 28200 3240 28212
rect 3195 28172 3240 28200
rect 3234 28160 3240 28172
rect 3292 28160 3298 28212
rect 6825 28203 6883 28209
rect 6825 28169 6837 28203
rect 6871 28200 6883 28203
rect 7006 28200 7012 28212
rect 6871 28172 7012 28200
rect 6871 28169 6883 28172
rect 6825 28163 6883 28169
rect 7006 28160 7012 28172
rect 7064 28160 7070 28212
rect 8110 28160 8116 28212
rect 8168 28200 8174 28212
rect 9493 28203 9551 28209
rect 8168 28172 9352 28200
rect 8168 28160 8174 28172
rect 1949 28135 2007 28141
rect 1949 28101 1961 28135
rect 1995 28132 2007 28135
rect 5442 28132 5448 28144
rect 1995 28104 5448 28132
rect 1995 28101 2007 28104
rect 1949 28095 2007 28101
rect 5442 28092 5448 28104
rect 5500 28132 5506 28144
rect 9217 28135 9275 28141
rect 9217 28132 9229 28135
rect 5500 28104 9229 28132
rect 5500 28092 5506 28104
rect 9217 28101 9229 28104
rect 9263 28101 9275 28135
rect 9217 28095 9275 28101
rect 9324 28132 9352 28172
rect 9493 28169 9505 28203
rect 9539 28200 9551 28203
rect 9582 28200 9588 28212
rect 9539 28172 9588 28200
rect 9539 28169 9551 28172
rect 9493 28163 9551 28169
rect 9582 28160 9588 28172
rect 9640 28160 9646 28212
rect 10689 28203 10747 28209
rect 10060 28172 10548 28200
rect 10060 28132 10088 28172
rect 10318 28132 10324 28144
rect 9324 28104 10088 28132
rect 10279 28104 10324 28132
rect 1762 28064 1768 28076
rect 1723 28036 1768 28064
rect 1762 28024 1768 28036
rect 1820 28024 1826 28076
rect 2314 28024 2320 28076
rect 2372 28064 2378 28076
rect 2593 28067 2651 28073
rect 2593 28064 2605 28067
rect 2372 28036 2605 28064
rect 2372 28024 2378 28036
rect 2593 28033 2605 28036
rect 2639 28033 2651 28067
rect 2593 28027 2651 28033
rect 2777 28067 2835 28073
rect 2777 28033 2789 28067
rect 2823 28033 2835 28067
rect 2777 28027 2835 28033
rect 2133 27999 2191 28005
rect 2133 27965 2145 27999
rect 2179 27996 2191 27999
rect 2792 27996 2820 28027
rect 2866 28024 2872 28076
rect 2924 28064 2930 28076
rect 3007 28067 3065 28073
rect 2924 28036 2969 28064
rect 2924 28024 2930 28036
rect 3007 28033 3019 28067
rect 3053 28064 3065 28067
rect 3697 28067 3755 28073
rect 3697 28064 3709 28067
rect 3053 28036 3709 28064
rect 3053 28033 3065 28036
rect 3007 28027 3065 28033
rect 3697 28033 3709 28036
rect 3743 28064 3755 28067
rect 5350 28064 5356 28076
rect 3743 28036 5356 28064
rect 3743 28033 3755 28036
rect 3697 28027 3755 28033
rect 5350 28024 5356 28036
rect 5408 28024 5414 28076
rect 5626 28064 5632 28076
rect 5587 28036 5632 28064
rect 5626 28024 5632 28036
rect 5684 28024 5690 28076
rect 5813 28067 5871 28073
rect 5813 28033 5825 28067
rect 5859 28064 5871 28067
rect 6457 28067 6515 28073
rect 6457 28064 6469 28067
rect 5859 28036 6469 28064
rect 5859 28033 5871 28036
rect 5813 28027 5871 28033
rect 6457 28033 6469 28036
rect 6503 28033 6515 28067
rect 6457 28027 6515 28033
rect 6641 28067 6699 28073
rect 6641 28033 6653 28067
rect 6687 28064 6699 28067
rect 6730 28064 6736 28076
rect 6687 28036 6736 28064
rect 6687 28033 6699 28036
rect 6641 28027 6699 28033
rect 2179 27968 2820 27996
rect 6472 27996 6500 28027
rect 6730 28024 6736 28036
rect 6788 28024 6794 28076
rect 7745 28067 7803 28073
rect 7745 28033 7757 28067
rect 7791 28033 7803 28067
rect 7745 28027 7803 28033
rect 7929 28067 7987 28073
rect 7929 28033 7941 28067
rect 7975 28033 7987 28067
rect 7929 28027 7987 28033
rect 7098 27996 7104 28008
rect 6472 27968 7104 27996
rect 2179 27965 2191 27968
rect 2133 27959 2191 27965
rect 7098 27956 7104 27968
rect 7156 27996 7162 28008
rect 7760 27996 7788 28027
rect 7156 27968 7788 27996
rect 7944 27996 7972 28027
rect 8202 28024 8208 28076
rect 8260 28064 8266 28076
rect 8941 28067 8999 28073
rect 8941 28064 8953 28067
rect 8260 28036 8953 28064
rect 8260 28024 8266 28036
rect 8941 28033 8953 28036
rect 8987 28033 8999 28067
rect 8941 28027 8999 28033
rect 9122 28024 9128 28076
rect 9180 28064 9186 28076
rect 9324 28073 9352 28104
rect 10318 28092 10324 28104
rect 10376 28092 10382 28144
rect 9309 28067 9367 28073
rect 9180 28036 9273 28064
rect 9180 28024 9186 28036
rect 9309 28033 9321 28067
rect 9355 28033 9367 28067
rect 10134 28064 10140 28076
rect 10095 28036 10140 28064
rect 9309 28027 9367 28033
rect 10134 28024 10140 28036
rect 10192 28024 10198 28076
rect 10410 28064 10416 28076
rect 10371 28036 10416 28064
rect 10410 28024 10416 28036
rect 10468 28024 10474 28076
rect 10520 28073 10548 28172
rect 10689 28169 10701 28203
rect 10735 28169 10747 28203
rect 10689 28163 10747 28169
rect 10505 28067 10563 28073
rect 10505 28033 10517 28067
rect 10551 28033 10563 28067
rect 10704 28064 10732 28163
rect 15286 28160 15292 28212
rect 15344 28200 15350 28212
rect 16025 28203 16083 28209
rect 16025 28200 16037 28203
rect 15344 28172 16037 28200
rect 15344 28160 15350 28172
rect 16025 28169 16037 28172
rect 16071 28169 16083 28203
rect 17862 28200 17868 28212
rect 17823 28172 17868 28200
rect 16025 28163 16083 28169
rect 17862 28160 17868 28172
rect 17920 28160 17926 28212
rect 20622 28200 20628 28212
rect 20583 28172 20628 28200
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 22094 28200 22100 28212
rect 21008 28172 22100 28200
rect 11146 28092 11152 28144
rect 11204 28132 11210 28144
rect 11790 28132 11796 28144
rect 11204 28104 11796 28132
rect 11204 28092 11210 28104
rect 11790 28092 11796 28104
rect 11848 28132 11854 28144
rect 11885 28135 11943 28141
rect 11885 28132 11897 28135
rect 11848 28104 11897 28132
rect 11848 28092 11854 28104
rect 11885 28101 11897 28104
rect 11931 28101 11943 28135
rect 11885 28095 11943 28101
rect 11977 28135 12035 28141
rect 11977 28101 11989 28135
rect 12023 28132 12035 28135
rect 12158 28132 12164 28144
rect 12023 28104 12164 28132
rect 12023 28101 12035 28104
rect 11977 28095 12035 28101
rect 12158 28092 12164 28104
rect 12216 28092 12222 28144
rect 17126 28132 17132 28144
rect 14389 28104 17132 28132
rect 11609 28067 11667 28073
rect 11609 28064 11621 28067
rect 10704 28036 11621 28064
rect 10505 28027 10563 28033
rect 11609 28033 11621 28036
rect 11655 28033 11667 28067
rect 11609 28027 11667 28033
rect 11702 28067 11760 28073
rect 11702 28033 11714 28067
rect 11748 28033 11760 28067
rect 11702 28027 11760 28033
rect 12074 28067 12132 28073
rect 12074 28033 12086 28067
rect 12120 28064 12132 28067
rect 12710 28064 12716 28076
rect 12120 28036 12716 28064
rect 12120 28033 12132 28036
rect 12074 28027 12132 28033
rect 9140 27996 9168 28024
rect 10226 27996 10232 28008
rect 7944 27968 8432 27996
rect 9140 27968 10232 27996
rect 7156 27956 7162 27968
rect 8404 27928 8432 27968
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 10318 27928 10324 27940
rect 8404 27900 10324 27928
rect 10318 27888 10324 27900
rect 10376 27888 10382 27940
rect 11717 27928 11745 28027
rect 11882 27956 11888 28008
rect 11940 27996 11946 28008
rect 12089 27996 12117 28027
rect 12710 28024 12716 28036
rect 12768 28024 12774 28076
rect 13262 28064 13268 28076
rect 13223 28036 13268 28064
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 11940 27968 12117 27996
rect 13541 27999 13599 28005
rect 11940 27956 11946 27968
rect 13541 27965 13553 27999
rect 13587 27996 13599 27999
rect 14090 27996 14096 28008
rect 13587 27968 14096 27996
rect 13587 27965 13599 27968
rect 13541 27959 13599 27965
rect 14090 27956 14096 27968
rect 14148 27956 14154 28008
rect 14389 27928 14417 28104
rect 17126 28092 17132 28104
rect 17184 28092 17190 28144
rect 17954 28132 17960 28144
rect 17236 28104 17960 28132
rect 14734 28024 14740 28076
rect 14792 28064 14798 28076
rect 15114 28067 15172 28073
rect 15114 28064 15126 28067
rect 14792 28036 15126 28064
rect 14792 28024 14798 28036
rect 15114 28033 15126 28036
rect 15160 28033 15172 28067
rect 15114 28027 15172 28033
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28064 15899 28067
rect 15930 28064 15936 28076
rect 15887 28036 15936 28064
rect 15887 28033 15899 28036
rect 15841 28027 15899 28033
rect 15930 28024 15936 28036
rect 15988 28024 15994 28076
rect 17236 28073 17264 28104
rect 17954 28092 17960 28104
rect 18012 28092 18018 28144
rect 17221 28067 17279 28073
rect 17221 28033 17233 28067
rect 17267 28033 17279 28067
rect 17402 28064 17408 28076
rect 17363 28036 17408 28064
rect 17221 28027 17279 28033
rect 17402 28024 17408 28036
rect 17460 28024 17466 28076
rect 17497 28067 17555 28073
rect 17497 28033 17509 28067
rect 17543 28033 17555 28067
rect 17497 28027 17555 28033
rect 17589 28067 17647 28073
rect 17589 28033 17601 28067
rect 17635 28064 17647 28067
rect 18325 28067 18383 28073
rect 18325 28064 18337 28067
rect 17635 28036 18337 28064
rect 17635 28033 17647 28036
rect 17589 28027 17647 28033
rect 18325 28033 18337 28036
rect 18371 28033 18383 28067
rect 18325 28027 18383 28033
rect 15381 27999 15439 28005
rect 15381 27965 15393 27999
rect 15427 27965 15439 27999
rect 15381 27959 15439 27965
rect 11717 27900 14417 27928
rect 5445 27863 5503 27869
rect 5445 27829 5457 27863
rect 5491 27860 5503 27863
rect 6822 27860 6828 27872
rect 5491 27832 6828 27860
rect 5491 27829 5503 27832
rect 5445 27823 5503 27829
rect 6822 27820 6828 27832
rect 6880 27820 6886 27872
rect 7926 27820 7932 27872
rect 7984 27860 7990 27872
rect 8113 27863 8171 27869
rect 8113 27860 8125 27863
rect 7984 27832 8125 27860
rect 7984 27820 7990 27832
rect 8113 27829 8125 27832
rect 8159 27829 8171 27863
rect 12250 27860 12256 27872
rect 12211 27832 12256 27860
rect 8113 27823 8171 27829
rect 12250 27820 12256 27832
rect 12308 27820 12314 27872
rect 12986 27820 12992 27872
rect 13044 27860 13050 27872
rect 14001 27863 14059 27869
rect 14001 27860 14013 27863
rect 13044 27832 14013 27860
rect 13044 27820 13050 27832
rect 14001 27829 14013 27832
rect 14047 27829 14059 27863
rect 15396 27860 15424 27959
rect 16574 27956 16580 28008
rect 16632 27996 16638 28008
rect 17512 27996 17540 28027
rect 16632 27968 17540 27996
rect 16632 27956 16638 27968
rect 15470 27888 15476 27940
rect 15528 27928 15534 27940
rect 17604 27928 17632 28027
rect 15528 27900 17632 27928
rect 15528 27888 15534 27900
rect 18046 27860 18052 27872
rect 15396 27832 18052 27860
rect 14001 27823 14059 27829
rect 18046 27820 18052 27832
rect 18104 27820 18110 27872
rect 18340 27860 18368 28027
rect 18874 28024 18880 28076
rect 18932 28064 18938 28076
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 18932 28036 19073 28064
rect 18932 28024 18938 28036
rect 19061 28033 19073 28036
rect 19107 28064 19119 28067
rect 19797 28067 19855 28073
rect 19797 28064 19809 28067
rect 19107 28036 19809 28064
rect 19107 28033 19119 28036
rect 19061 28027 19119 28033
rect 19797 28033 19809 28036
rect 19843 28033 19855 28067
rect 20898 28064 20904 28076
rect 20859 28036 20904 28064
rect 19797 28027 19855 28033
rect 20898 28024 20904 28036
rect 20956 28024 20962 28076
rect 21008 28073 21036 28172
rect 22094 28160 22100 28172
rect 22152 28160 22158 28212
rect 25222 28200 25228 28212
rect 25183 28172 25228 28200
rect 25222 28160 25228 28172
rect 25280 28160 25286 28212
rect 25774 28160 25780 28212
rect 25832 28200 25838 28212
rect 26329 28203 26387 28209
rect 26329 28200 26341 28203
rect 25832 28172 26341 28200
rect 25832 28160 25838 28172
rect 26329 28169 26341 28172
rect 26375 28200 26387 28203
rect 27338 28200 27344 28212
rect 26375 28172 27344 28200
rect 26375 28169 26387 28172
rect 26329 28163 26387 28169
rect 27338 28160 27344 28172
rect 27396 28160 27402 28212
rect 27617 28203 27675 28209
rect 27617 28169 27629 28203
rect 27663 28200 27675 28203
rect 27798 28200 27804 28212
rect 27663 28172 27804 28200
rect 27663 28169 27675 28172
rect 27617 28163 27675 28169
rect 27798 28160 27804 28172
rect 27856 28160 27862 28212
rect 28166 28200 28172 28212
rect 28127 28172 28172 28200
rect 28166 28160 28172 28172
rect 28224 28160 28230 28212
rect 28902 28200 28908 28212
rect 28736 28172 28908 28200
rect 22186 28132 22192 28144
rect 22147 28104 22192 28132
rect 22186 28092 22192 28104
rect 22244 28092 22250 28144
rect 22370 28132 22376 28144
rect 22331 28104 22376 28132
rect 22370 28092 22376 28104
rect 22428 28092 22434 28144
rect 23100 28135 23158 28141
rect 23100 28101 23112 28135
rect 23146 28132 23158 28135
rect 23198 28132 23204 28144
rect 23146 28104 23204 28132
rect 23146 28101 23158 28104
rect 23100 28095 23158 28101
rect 23198 28092 23204 28104
rect 23256 28092 23262 28144
rect 23750 28092 23756 28144
rect 23808 28132 23814 28144
rect 26418 28132 26424 28144
rect 23808 28104 26424 28132
rect 23808 28092 23814 28104
rect 20993 28067 21051 28073
rect 20993 28033 21005 28067
rect 21039 28033 21051 28067
rect 20993 28027 21051 28033
rect 21082 28024 21088 28076
rect 21140 28064 21146 28076
rect 21140 28036 21185 28064
rect 21140 28024 21146 28036
rect 21266 28024 21272 28076
rect 21324 28064 21330 28076
rect 25608 28073 25636 28104
rect 26418 28092 26424 28104
rect 26476 28132 26482 28144
rect 26476 28104 27292 28132
rect 26476 28092 26482 28104
rect 25501 28067 25559 28073
rect 21324 28036 21369 28064
rect 21324 28024 21330 28036
rect 25501 28033 25513 28067
rect 25547 28033 25559 28067
rect 25501 28027 25559 28033
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27996 19671 27999
rect 21542 27996 21548 28008
rect 19659 27968 21548 27996
rect 19659 27965 19671 27968
rect 19613 27959 19671 27965
rect 21542 27956 21548 27968
rect 21600 27956 21606 28008
rect 22830 27996 22836 28008
rect 22791 27968 22836 27996
rect 22830 27956 22836 27968
rect 22888 27956 22894 28008
rect 25516 27996 25544 28027
rect 25682 28024 25688 28076
rect 25740 28064 25746 28076
rect 27264 28073 27292 28104
rect 27356 28073 27384 28160
rect 25869 28067 25927 28073
rect 25740 28036 25785 28064
rect 25740 28024 25746 28036
rect 25869 28033 25881 28067
rect 25915 28064 25927 28067
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 25915 28036 26985 28064
rect 25915 28033 25927 28036
rect 25869 28027 25927 28033
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27157 28067 27215 28073
rect 27157 28033 27169 28067
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 27249 28067 27307 28073
rect 27249 28033 27261 28067
rect 27295 28033 27307 28067
rect 27249 28027 27307 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28033 27399 28067
rect 27341 28027 27399 28033
rect 25516 27968 25636 27996
rect 24394 27928 24400 27940
rect 24136 27900 24400 27928
rect 19978 27860 19984 27872
rect 18340 27832 19984 27860
rect 19978 27820 19984 27832
rect 20036 27860 20042 27872
rect 24136 27860 24164 27900
rect 24394 27888 24400 27900
rect 24452 27928 24458 27940
rect 24452 27900 24808 27928
rect 24452 27888 24458 27900
rect 20036 27832 24164 27860
rect 24213 27863 24271 27869
rect 20036 27820 20042 27832
rect 24213 27829 24225 27863
rect 24259 27860 24271 27863
rect 24578 27860 24584 27872
rect 24259 27832 24584 27860
rect 24259 27829 24271 27832
rect 24213 27823 24271 27829
rect 24578 27820 24584 27832
rect 24636 27820 24642 27872
rect 24780 27869 24808 27900
rect 24765 27863 24823 27869
rect 24765 27829 24777 27863
rect 24811 27860 24823 27863
rect 25608 27860 25636 27968
rect 25774 27956 25780 28008
rect 25832 27996 25838 28008
rect 25884 27996 25912 28027
rect 25832 27968 25912 27996
rect 25832 27956 25838 27968
rect 26142 27956 26148 28008
rect 26200 27996 26206 28008
rect 27172 27996 27200 28027
rect 28074 28024 28080 28076
rect 28132 28064 28138 28076
rect 28736 28073 28764 28172
rect 28902 28160 28908 28172
rect 28960 28160 28966 28212
rect 28994 28160 29000 28212
rect 29052 28160 29058 28212
rect 30469 28203 30527 28209
rect 30469 28169 30481 28203
rect 30515 28200 30527 28203
rect 30650 28200 30656 28212
rect 30515 28172 30656 28200
rect 30515 28169 30527 28172
rect 30469 28163 30527 28169
rect 30650 28160 30656 28172
rect 30708 28160 30714 28212
rect 29012 28079 29040 28160
rect 29365 28135 29423 28141
rect 29365 28101 29377 28135
rect 29411 28132 29423 28135
rect 30374 28132 30380 28144
rect 29411 28104 30380 28132
rect 29411 28101 29423 28104
rect 29365 28095 29423 28101
rect 30374 28092 30380 28104
rect 30432 28092 30438 28144
rect 32122 28132 32128 28144
rect 30668 28104 32128 28132
rect 28984 28073 29042 28079
rect 29178 28073 29184 28076
rect 28721 28067 28779 28073
rect 28721 28064 28733 28067
rect 28132 28036 28733 28064
rect 28132 28024 28138 28036
rect 28721 28033 28733 28036
rect 28767 28033 28779 28067
rect 28721 28027 28779 28033
rect 28884 28067 28942 28073
rect 28884 28033 28896 28067
rect 28930 28064 28942 28067
rect 28930 28033 28948 28064
rect 28984 28039 28996 28073
rect 29030 28039 29042 28073
rect 28984 28033 29042 28039
rect 29135 28067 29184 28073
rect 29135 28033 29147 28067
rect 29181 28033 29184 28067
rect 28884 28027 28948 28033
rect 29135 28027 29184 28033
rect 26200 27968 27200 27996
rect 28920 27996 28948 28027
rect 29178 28024 29184 28027
rect 29236 28064 29242 28076
rect 30668 28073 30696 28104
rect 32122 28092 32128 28104
rect 32180 28092 32186 28144
rect 29825 28067 29883 28073
rect 29825 28064 29837 28067
rect 29236 28036 29837 28064
rect 29236 28024 29242 28036
rect 29825 28033 29837 28036
rect 29871 28033 29883 28067
rect 30653 28067 30711 28073
rect 30653 28064 30665 28067
rect 29825 28027 29883 28033
rect 30392 28036 30665 28064
rect 30392 28008 30420 28036
rect 30653 28033 30665 28036
rect 30699 28033 30711 28067
rect 30834 28064 30840 28076
rect 30795 28036 30840 28064
rect 30653 28027 30711 28033
rect 30834 28024 30840 28036
rect 30892 28024 30898 28076
rect 32490 28024 32496 28076
rect 32548 28064 32554 28076
rect 33238 28067 33296 28073
rect 33238 28064 33250 28067
rect 32548 28036 33250 28064
rect 32548 28024 32554 28036
rect 33238 28033 33250 28036
rect 33284 28033 33296 28067
rect 33502 28064 33508 28076
rect 33463 28036 33508 28064
rect 33238 28027 33296 28033
rect 33502 28024 33508 28036
rect 33560 28024 33566 28076
rect 29362 27996 29368 28008
rect 28920 27968 29368 27996
rect 26200 27956 26206 27968
rect 29362 27956 29368 27968
rect 29420 27956 29426 28008
rect 30374 27956 30380 28008
rect 30432 27956 30438 28008
rect 67634 27928 67640 27940
rect 67595 27900 67640 27928
rect 67634 27888 67640 27900
rect 67692 27888 67698 27940
rect 31018 27860 31024 27872
rect 24811 27832 31024 27860
rect 24811 27829 24823 27832
rect 24765 27823 24823 27829
rect 31018 27820 31024 27832
rect 31076 27820 31082 27872
rect 32122 27860 32128 27872
rect 32083 27832 32128 27860
rect 32122 27820 32128 27832
rect 32180 27820 32186 27872
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 5626 27616 5632 27668
rect 5684 27656 5690 27668
rect 10778 27656 10784 27668
rect 5684 27628 10784 27656
rect 5684 27616 5690 27628
rect 10778 27616 10784 27628
rect 10836 27616 10842 27668
rect 11330 27616 11336 27668
rect 11388 27656 11394 27668
rect 14734 27656 14740 27668
rect 11388 27628 12296 27656
rect 14695 27628 14740 27656
rect 11388 27616 11394 27628
rect 1581 27591 1639 27597
rect 1581 27557 1593 27591
rect 1627 27588 1639 27591
rect 2590 27588 2596 27600
rect 1627 27560 2596 27588
rect 1627 27557 1639 27560
rect 1581 27551 1639 27557
rect 2590 27548 2596 27560
rect 2648 27548 2654 27600
rect 2685 27591 2743 27597
rect 2685 27557 2697 27591
rect 2731 27588 2743 27591
rect 3326 27588 3332 27600
rect 2731 27560 3332 27588
rect 2731 27557 2743 27560
rect 2685 27551 2743 27557
rect 3326 27548 3332 27560
rect 3384 27548 3390 27600
rect 5261 27591 5319 27597
rect 5261 27557 5273 27591
rect 5307 27588 5319 27591
rect 5644 27588 5672 27616
rect 10318 27588 10324 27600
rect 5307 27560 5672 27588
rect 10279 27560 10324 27588
rect 5307 27557 5319 27560
rect 5261 27551 5319 27557
rect 10318 27548 10324 27560
rect 10376 27548 10382 27600
rect 11238 27548 11244 27600
rect 11296 27588 11302 27600
rect 11517 27591 11575 27597
rect 11517 27588 11529 27591
rect 11296 27560 11529 27588
rect 11296 27548 11302 27560
rect 11517 27557 11529 27560
rect 11563 27557 11575 27591
rect 12268 27588 12296 27628
rect 14734 27616 14740 27628
rect 14792 27616 14798 27668
rect 17494 27616 17500 27668
rect 17552 27656 17558 27668
rect 20438 27656 20444 27668
rect 17552 27628 20444 27656
rect 17552 27616 17558 27628
rect 20438 27616 20444 27628
rect 20496 27656 20502 27668
rect 20898 27656 20904 27668
rect 20496 27628 20904 27656
rect 20496 27616 20502 27628
rect 20898 27616 20904 27628
rect 20956 27616 20962 27668
rect 24302 27616 24308 27668
rect 24360 27656 24366 27668
rect 24397 27659 24455 27665
rect 24397 27656 24409 27659
rect 24360 27628 24409 27656
rect 24360 27616 24366 27628
rect 24397 27625 24409 27628
rect 24443 27625 24455 27659
rect 24397 27619 24455 27625
rect 24877 27628 25360 27656
rect 17129 27591 17187 27597
rect 17129 27588 17141 27591
rect 12268 27560 17141 27588
rect 11517 27551 11575 27557
rect 17129 27557 17141 27560
rect 17175 27588 17187 27591
rect 18138 27588 18144 27600
rect 17175 27560 18144 27588
rect 17175 27557 17187 27560
rect 17129 27551 17187 27557
rect 18138 27548 18144 27560
rect 18196 27548 18202 27600
rect 21453 27591 21511 27597
rect 21453 27557 21465 27591
rect 21499 27588 21511 27591
rect 24877 27588 24905 27628
rect 21499 27560 24905 27588
rect 21499 27557 21511 27560
rect 21453 27551 21511 27557
rect 2866 27520 2872 27532
rect 2332 27492 2872 27520
rect 2041 27455 2099 27461
rect 2041 27421 2053 27455
rect 2087 27421 2099 27455
rect 2222 27452 2228 27464
rect 2183 27424 2228 27452
rect 2041 27415 2099 27421
rect 2056 27384 2084 27415
rect 2222 27412 2228 27424
rect 2280 27412 2286 27464
rect 2332 27461 2360 27492
rect 2866 27480 2872 27492
rect 2924 27480 2930 27532
rect 6641 27523 6699 27529
rect 6641 27489 6653 27523
rect 6687 27520 6699 27523
rect 15562 27520 15568 27532
rect 6687 27492 8984 27520
rect 6687 27489 6699 27492
rect 6641 27483 6699 27489
rect 2317 27455 2375 27461
rect 2317 27421 2329 27455
rect 2363 27421 2375 27455
rect 2317 27415 2375 27421
rect 2409 27455 2467 27461
rect 2409 27421 2421 27455
rect 2455 27452 2467 27455
rect 2590 27452 2596 27464
rect 2455 27424 2596 27452
rect 2455 27421 2467 27424
rect 2409 27415 2467 27421
rect 2590 27412 2596 27424
rect 2648 27452 2654 27464
rect 7193 27455 7251 27461
rect 7193 27452 7205 27455
rect 2648 27424 7205 27452
rect 2648 27412 2654 27424
rect 7193 27421 7205 27424
rect 7239 27421 7251 27455
rect 7742 27452 7748 27464
rect 7703 27424 7748 27452
rect 7193 27415 7251 27421
rect 6396 27387 6454 27393
rect 2056 27356 2360 27384
rect 2332 27328 2360 27356
rect 6396 27353 6408 27387
rect 6442 27384 6454 27387
rect 6546 27384 6552 27396
rect 6442 27356 6552 27384
rect 6442 27353 6454 27356
rect 6396 27347 6454 27353
rect 6546 27344 6552 27356
rect 6604 27344 6610 27396
rect 7208 27384 7236 27415
rect 7742 27412 7748 27424
rect 7800 27412 7806 27464
rect 7926 27452 7932 27464
rect 7887 27424 7932 27452
rect 7926 27412 7932 27424
rect 7984 27412 7990 27464
rect 8018 27412 8024 27464
rect 8076 27452 8082 27464
rect 8956 27461 8984 27492
rect 11256 27492 15568 27520
rect 8159 27455 8217 27461
rect 8076 27424 8121 27452
rect 8076 27412 8082 27424
rect 8159 27421 8171 27455
rect 8205 27452 8217 27455
rect 8941 27455 8999 27461
rect 8205 27421 8239 27452
rect 8159 27415 8239 27421
rect 8941 27421 8953 27455
rect 8987 27452 8999 27455
rect 10502 27452 10508 27464
rect 8987 27424 10508 27452
rect 8987 27421 8999 27424
rect 8941 27415 8999 27421
rect 8211 27384 8239 27415
rect 10502 27412 10508 27424
rect 10560 27412 10566 27464
rect 10870 27452 10876 27464
rect 10831 27424 10876 27452
rect 10870 27412 10876 27424
rect 10928 27412 10934 27464
rect 11021 27455 11079 27461
rect 11021 27421 11033 27455
rect 11067 27452 11079 27455
rect 11256 27452 11284 27492
rect 15562 27480 15568 27492
rect 15620 27480 15626 27532
rect 16209 27523 16267 27529
rect 16209 27489 16221 27523
rect 16255 27520 16267 27523
rect 16574 27520 16580 27532
rect 16255 27492 16580 27520
rect 16255 27489 16267 27492
rect 16209 27483 16267 27489
rect 16574 27480 16580 27492
rect 16632 27480 16638 27532
rect 17770 27480 17776 27532
rect 17828 27520 17834 27532
rect 21468 27520 21496 27551
rect 25130 27548 25136 27600
rect 25188 27588 25194 27600
rect 25225 27591 25283 27597
rect 25225 27588 25237 27591
rect 25188 27560 25237 27588
rect 25188 27548 25194 27560
rect 25225 27557 25237 27560
rect 25271 27557 25283 27591
rect 25332 27588 25360 27628
rect 25976 27628 26280 27656
rect 25976 27588 26004 27628
rect 26142 27588 26148 27600
rect 25332 27560 26004 27588
rect 26103 27560 26148 27588
rect 25225 27551 25283 27557
rect 26142 27548 26148 27560
rect 26200 27548 26206 27600
rect 26252 27588 26280 27628
rect 27706 27588 27712 27600
rect 26252 27560 27712 27588
rect 27706 27548 27712 27560
rect 27764 27548 27770 27600
rect 30745 27591 30803 27597
rect 30745 27557 30757 27591
rect 30791 27588 30803 27591
rect 32490 27588 32496 27600
rect 30791 27560 32496 27588
rect 30791 27557 30803 27560
rect 30745 27551 30803 27557
rect 32490 27548 32496 27560
rect 32548 27548 32554 27600
rect 17828 27492 21496 27520
rect 17828 27480 17834 27492
rect 22094 27480 22100 27532
rect 22152 27520 22158 27532
rect 22281 27523 22339 27529
rect 22281 27520 22293 27523
rect 22152 27492 22293 27520
rect 22152 27480 22158 27492
rect 22281 27489 22293 27492
rect 22327 27489 22339 27523
rect 27801 27523 27859 27529
rect 27801 27520 27813 27523
rect 22281 27483 22339 27489
rect 24412 27492 27813 27520
rect 11067 27424 11284 27452
rect 11379 27455 11437 27461
rect 11067 27421 11079 27424
rect 11021 27415 11079 27421
rect 11379 27421 11391 27455
rect 11425 27452 11437 27455
rect 11882 27452 11888 27464
rect 11425 27424 11888 27452
rect 11425 27421 11437 27424
rect 11379 27415 11437 27421
rect 11882 27412 11888 27424
rect 11940 27412 11946 27464
rect 12713 27455 12771 27461
rect 12713 27421 12725 27455
rect 12759 27452 12771 27455
rect 12759 27424 12940 27452
rect 12759 27421 12771 27424
rect 12713 27415 12771 27421
rect 12912 27396 12940 27424
rect 12986 27412 12992 27464
rect 13044 27452 13050 27464
rect 13357 27455 13415 27461
rect 13357 27452 13369 27455
rect 13044 27424 13369 27452
rect 13044 27412 13050 27424
rect 13357 27421 13369 27424
rect 13403 27421 13415 27455
rect 13357 27415 13415 27421
rect 14093 27455 14151 27461
rect 14093 27421 14105 27455
rect 14139 27452 14151 27455
rect 14182 27452 14188 27464
rect 14139 27424 14188 27452
rect 14139 27421 14151 27424
rect 14093 27415 14151 27421
rect 14182 27412 14188 27424
rect 14240 27412 14246 27464
rect 14277 27455 14335 27461
rect 14277 27421 14289 27455
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27421 14427 27455
rect 14369 27415 14427 27421
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27452 14519 27455
rect 15194 27452 15200 27464
rect 14507 27424 15200 27452
rect 14507 27421 14519 27424
rect 14461 27415 14519 27421
rect 7208 27356 8239 27384
rect 8389 27387 8447 27393
rect 8389 27353 8401 27387
rect 8435 27384 8447 27387
rect 9186 27387 9244 27393
rect 9186 27384 9198 27387
rect 8435 27356 9198 27384
rect 8435 27353 8447 27356
rect 8389 27347 8447 27353
rect 9186 27353 9198 27356
rect 9232 27353 9244 27387
rect 11146 27384 11152 27396
rect 11107 27356 11152 27384
rect 9186 27347 9244 27353
rect 11146 27344 11152 27356
rect 11204 27344 11210 27396
rect 11241 27387 11299 27393
rect 11241 27353 11253 27387
rect 11287 27384 11299 27387
rect 11287 27356 11376 27384
rect 11287 27353 11299 27356
rect 11241 27347 11299 27353
rect 2314 27276 2320 27328
rect 2372 27276 2378 27328
rect 7374 27276 7380 27328
rect 7432 27316 7438 27328
rect 8018 27316 8024 27328
rect 7432 27288 8024 27316
rect 7432 27276 7438 27288
rect 8018 27276 8024 27288
rect 8076 27276 8082 27328
rect 8202 27276 8208 27328
rect 8260 27316 8266 27328
rect 11348 27316 11376 27356
rect 12894 27344 12900 27396
rect 12952 27384 12958 27396
rect 13173 27387 13231 27393
rect 13173 27384 13185 27387
rect 12952 27356 13185 27384
rect 12952 27344 12958 27356
rect 13173 27353 13185 27356
rect 13219 27353 13231 27387
rect 13173 27347 13231 27353
rect 13541 27387 13599 27393
rect 13541 27353 13553 27387
rect 13587 27384 13599 27387
rect 14292 27384 14320 27415
rect 13587 27356 14320 27384
rect 13587 27353 13599 27356
rect 13541 27347 13599 27353
rect 8260 27288 11376 27316
rect 8260 27276 8266 27288
rect 12066 27276 12072 27328
rect 12124 27316 12130 27328
rect 12529 27319 12587 27325
rect 12529 27316 12541 27319
rect 12124 27288 12541 27316
rect 12124 27276 12130 27288
rect 12529 27285 12541 27288
rect 12575 27285 12587 27319
rect 12529 27279 12587 27285
rect 14090 27276 14096 27328
rect 14148 27316 14154 27328
rect 14384 27316 14412 27415
rect 15194 27412 15200 27424
rect 15252 27412 15258 27464
rect 16298 27412 16304 27464
rect 16356 27452 16362 27464
rect 16485 27455 16543 27461
rect 16485 27452 16497 27455
rect 16356 27424 16497 27452
rect 16356 27412 16362 27424
rect 16485 27421 16497 27424
rect 16531 27421 16543 27455
rect 16485 27415 16543 27421
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 18233 27455 18291 27461
rect 18233 27452 18245 27455
rect 18012 27424 18245 27452
rect 18012 27412 18018 27424
rect 18233 27421 18245 27424
rect 18279 27421 18291 27455
rect 18506 27452 18512 27464
rect 18467 27424 18512 27452
rect 18233 27415 18291 27421
rect 18506 27412 18512 27424
rect 18564 27452 18570 27464
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 18564 27424 21281 27452
rect 18564 27412 18570 27424
rect 21269 27421 21281 27424
rect 21315 27421 21327 27455
rect 22002 27452 22008 27464
rect 21963 27424 22008 27452
rect 21269 27415 21327 27421
rect 16574 27344 16580 27396
rect 16632 27384 16638 27396
rect 17586 27384 17592 27396
rect 16632 27356 17592 27384
rect 16632 27344 16638 27356
rect 17586 27344 17592 27356
rect 17644 27384 17650 27396
rect 19245 27387 19303 27393
rect 19245 27384 19257 27387
rect 17644 27356 19257 27384
rect 17644 27344 17650 27356
rect 19245 27353 19257 27356
rect 19291 27353 19303 27387
rect 19426 27384 19432 27396
rect 19387 27356 19432 27384
rect 19245 27347 19303 27353
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 21284 27384 21312 27415
rect 22002 27412 22008 27424
rect 22060 27412 22066 27464
rect 24412 27384 24440 27492
rect 27801 27489 27813 27492
rect 27847 27520 27859 27523
rect 27982 27520 27988 27532
rect 27847 27492 27988 27520
rect 27847 27489 27859 27492
rect 27801 27483 27859 27489
rect 27982 27480 27988 27492
rect 28040 27480 28046 27532
rect 30558 27520 30564 27532
rect 30392 27492 30564 27520
rect 25590 27412 25596 27464
rect 25648 27452 25654 27464
rect 25961 27455 26019 27461
rect 25961 27452 25973 27455
rect 25648 27424 25973 27452
rect 25648 27412 25654 27424
rect 25961 27421 25973 27424
rect 26007 27421 26019 27455
rect 28074 27452 28080 27464
rect 28035 27424 28080 27452
rect 25961 27415 26019 27421
rect 28074 27412 28080 27424
rect 28132 27452 28138 27464
rect 30101 27455 30159 27461
rect 30101 27452 30113 27455
rect 28132 27424 30113 27452
rect 28132 27412 28138 27424
rect 30101 27421 30113 27424
rect 30147 27421 30159 27455
rect 30282 27452 30288 27464
rect 30243 27424 30288 27452
rect 30101 27415 30159 27421
rect 30282 27412 30288 27424
rect 30340 27412 30346 27464
rect 30392 27461 30420 27492
rect 30558 27480 30564 27492
rect 30616 27520 30622 27532
rect 30616 27492 30788 27520
rect 30616 27480 30622 27492
rect 30760 27464 30788 27492
rect 30377 27455 30435 27461
rect 30377 27421 30389 27455
rect 30423 27421 30435 27455
rect 30377 27415 30435 27421
rect 30469 27455 30527 27461
rect 30469 27421 30481 27455
rect 30515 27421 30527 27455
rect 30469 27415 30527 27421
rect 24578 27384 24584 27396
rect 21284 27356 24440 27384
rect 24539 27356 24584 27384
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 24765 27387 24823 27393
rect 24765 27353 24777 27387
rect 24811 27384 24823 27387
rect 24854 27384 24860 27396
rect 24811 27356 24860 27384
rect 24811 27353 24823 27356
rect 24765 27347 24823 27353
rect 24854 27344 24860 27356
rect 24912 27384 24918 27396
rect 25777 27387 25835 27393
rect 25777 27384 25789 27387
rect 24912 27356 25789 27384
rect 24912 27344 24918 27356
rect 25777 27353 25789 27356
rect 25823 27384 25835 27387
rect 26142 27384 26148 27396
rect 25823 27356 26148 27384
rect 25823 27353 25835 27356
rect 25777 27347 25835 27353
rect 26142 27344 26148 27356
rect 26200 27344 26206 27396
rect 26326 27344 26332 27396
rect 26384 27384 26390 27396
rect 29549 27387 29607 27393
rect 29549 27384 29561 27387
rect 26384 27356 29561 27384
rect 26384 27344 26390 27356
rect 29549 27353 29561 27356
rect 29595 27384 29607 27387
rect 30484 27384 30512 27415
rect 30742 27412 30748 27464
rect 30800 27412 30806 27464
rect 29595 27356 30512 27384
rect 29595 27353 29607 27356
rect 29549 27347 29607 27353
rect 14148 27288 14412 27316
rect 14148 27276 14154 27288
rect 18230 27276 18236 27328
rect 18288 27316 18294 27328
rect 19613 27319 19671 27325
rect 19613 27316 19625 27319
rect 18288 27288 19625 27316
rect 18288 27276 18294 27288
rect 19613 27285 19625 27288
rect 19659 27285 19671 27319
rect 19613 27279 19671 27285
rect 25222 27276 25228 27328
rect 25280 27316 25286 27328
rect 25682 27316 25688 27328
rect 25280 27288 25688 27316
rect 25280 27276 25286 27288
rect 25682 27276 25688 27288
rect 25740 27316 25746 27328
rect 26694 27316 26700 27328
rect 25740 27288 26700 27316
rect 25740 27276 25746 27288
rect 26694 27276 26700 27288
rect 26752 27276 26758 27328
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 6546 27112 6552 27124
rect 6507 27084 6552 27112
rect 6546 27072 6552 27084
rect 6604 27072 6610 27124
rect 10226 27072 10232 27124
rect 10284 27112 10290 27124
rect 10870 27112 10876 27124
rect 10284 27084 10732 27112
rect 10831 27084 10876 27112
rect 10284 27072 10290 27084
rect 2961 27047 3019 27053
rect 2961 27013 2973 27047
rect 3007 27044 3019 27047
rect 3666 27047 3724 27053
rect 3666 27044 3678 27047
rect 3007 27016 3678 27044
rect 3007 27013 3019 27016
rect 2961 27007 3019 27013
rect 3666 27013 3678 27016
rect 3712 27013 3724 27047
rect 3666 27007 3724 27013
rect 10134 27004 10140 27056
rect 10192 27044 10198 27056
rect 10505 27047 10563 27053
rect 10505 27044 10517 27047
rect 10192 27016 10517 27044
rect 10192 27004 10198 27016
rect 10505 27013 10517 27016
rect 10551 27013 10563 27047
rect 10704 27044 10732 27084
rect 10870 27072 10876 27084
rect 10928 27072 10934 27124
rect 16117 27115 16175 27121
rect 16117 27081 16129 27115
rect 16163 27112 16175 27115
rect 16574 27112 16580 27124
rect 16163 27084 16580 27112
rect 16163 27081 16175 27084
rect 16117 27075 16175 27081
rect 16574 27072 16580 27084
rect 16632 27072 16638 27124
rect 20438 27112 20444 27124
rect 20399 27084 20444 27112
rect 20438 27072 20444 27084
rect 20496 27112 20502 27124
rect 23109 27115 23167 27121
rect 23109 27112 23121 27115
rect 20496 27084 23121 27112
rect 20496 27072 20502 27084
rect 23109 27081 23121 27084
rect 23155 27112 23167 27115
rect 23566 27112 23572 27124
rect 23155 27084 23572 27112
rect 23155 27081 23167 27084
rect 23109 27075 23167 27081
rect 23566 27072 23572 27084
rect 23624 27112 23630 27124
rect 29178 27112 29184 27124
rect 23624 27084 29184 27112
rect 23624 27072 23630 27084
rect 29178 27072 29184 27084
rect 29236 27072 29242 27124
rect 29362 27112 29368 27124
rect 29323 27084 29368 27112
rect 29362 27072 29368 27084
rect 29420 27072 29426 27124
rect 30282 27072 30288 27124
rect 30340 27112 30346 27124
rect 30377 27115 30435 27121
rect 30377 27112 30389 27115
rect 30340 27084 30389 27112
rect 30340 27072 30346 27084
rect 30377 27081 30389 27084
rect 30423 27081 30435 27115
rect 30377 27075 30435 27081
rect 18138 27044 18144 27056
rect 10704 27016 12756 27044
rect 18099 27016 18144 27044
rect 10505 27007 10563 27013
rect 2314 26976 2320 26988
rect 2275 26948 2320 26976
rect 2314 26936 2320 26948
rect 2372 26936 2378 26988
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 2593 26979 2651 26985
rect 2593 26945 2605 26979
rect 2639 26945 2651 26979
rect 2593 26939 2651 26945
rect 2685 26979 2743 26985
rect 2685 26945 2697 26979
rect 2731 26976 2743 26979
rect 3418 26976 3424 26988
rect 2731 26948 3280 26976
rect 3379 26948 3424 26976
rect 2731 26945 2743 26948
rect 2685 26939 2743 26945
rect 2608 26908 2636 26939
rect 2866 26908 2872 26920
rect 2608 26880 2872 26908
rect 2866 26868 2872 26880
rect 2924 26868 2930 26920
rect 3252 26908 3280 26948
rect 3418 26936 3424 26948
rect 3476 26936 3482 26988
rect 6825 26979 6883 26985
rect 6825 26976 6837 26979
rect 3528 26948 6837 26976
rect 3528 26908 3556 26948
rect 6825 26945 6837 26948
rect 6871 26945 6883 26979
rect 6825 26939 6883 26945
rect 6917 26979 6975 26985
rect 6917 26945 6929 26979
rect 6963 26945 6975 26979
rect 6917 26939 6975 26945
rect 3252 26880 3556 26908
rect 6840 26840 6868 26939
rect 6932 26908 6960 26939
rect 7006 26936 7012 26988
rect 7064 26976 7070 26988
rect 7193 26979 7251 26985
rect 7064 26948 7109 26976
rect 7064 26936 7070 26948
rect 7193 26945 7205 26979
rect 7239 26976 7251 26979
rect 7282 26976 7288 26988
rect 7239 26948 7288 26976
rect 7239 26945 7251 26948
rect 7193 26939 7251 26945
rect 7282 26936 7288 26948
rect 7340 26976 7346 26988
rect 7653 26979 7711 26985
rect 7653 26976 7665 26979
rect 7340 26948 7665 26976
rect 7340 26936 7346 26948
rect 7653 26945 7665 26948
rect 7699 26945 7711 26979
rect 7653 26939 7711 26945
rect 9674 26936 9680 26988
rect 9732 26976 9738 26988
rect 10321 26979 10379 26985
rect 10321 26976 10333 26979
rect 9732 26948 10333 26976
rect 9732 26936 9738 26948
rect 10321 26945 10333 26948
rect 10367 26945 10379 26979
rect 10321 26939 10379 26945
rect 10597 26979 10655 26985
rect 10597 26945 10609 26979
rect 10643 26945 10655 26979
rect 10597 26939 10655 26945
rect 7374 26908 7380 26920
rect 6932 26880 7380 26908
rect 7374 26868 7380 26880
rect 7432 26868 7438 26920
rect 7466 26868 7472 26920
rect 7524 26908 7530 26920
rect 10612 26908 10640 26939
rect 10686 26936 10692 26988
rect 10744 26976 10750 26988
rect 12728 26985 12756 27016
rect 18138 27004 18144 27016
rect 18196 27004 18202 27056
rect 20990 27004 20996 27056
rect 21048 27044 21054 27056
rect 22005 27047 22063 27053
rect 22005 27044 22017 27047
rect 21048 27016 22017 27044
rect 21048 27004 21054 27016
rect 22005 27013 22017 27016
rect 22051 27013 22063 27047
rect 22005 27007 22063 27013
rect 23753 27047 23811 27053
rect 23753 27013 23765 27047
rect 23799 27044 23811 27047
rect 24394 27044 24400 27056
rect 23799 27016 24400 27044
rect 23799 27013 23811 27016
rect 23753 27007 23811 27013
rect 24394 27004 24400 27016
rect 24452 27004 24458 27056
rect 25130 27004 25136 27056
rect 25188 27044 25194 27056
rect 26326 27044 26332 27056
rect 25188 27016 26332 27044
rect 25188 27004 25194 27016
rect 12713 26979 12771 26985
rect 10744 26948 10789 26976
rect 10744 26936 10750 26948
rect 12713 26945 12725 26979
rect 12759 26976 12771 26979
rect 13998 26976 14004 26988
rect 12759 26948 14004 26976
rect 12759 26945 12771 26948
rect 12713 26939 12771 26945
rect 13998 26936 14004 26948
rect 14056 26936 14062 26988
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 14185 26979 14243 26985
rect 14185 26976 14197 26979
rect 14148 26948 14197 26976
rect 14148 26936 14154 26948
rect 14185 26945 14197 26948
rect 14231 26945 14243 26979
rect 15930 26976 15936 26988
rect 15891 26948 15936 26976
rect 14185 26939 14243 26945
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 20162 26936 20168 26988
rect 20220 26976 20226 26988
rect 20533 26979 20591 26985
rect 20533 26976 20545 26979
rect 20220 26948 20545 26976
rect 20220 26936 20226 26948
rect 20533 26945 20545 26948
rect 20579 26976 20591 26979
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 20579 26948 21097 26976
rect 20579 26945 20591 26948
rect 20533 26939 20591 26945
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 21174 26936 21180 26988
rect 21232 26976 21238 26988
rect 21818 26976 21824 26988
rect 21232 26948 21824 26976
rect 21232 26936 21238 26948
rect 21818 26936 21824 26948
rect 21876 26936 21882 26988
rect 23198 26936 23204 26988
rect 23256 26976 23262 26988
rect 23937 26979 23995 26985
rect 23937 26976 23949 26979
rect 23256 26948 23949 26976
rect 23256 26936 23262 26948
rect 23937 26945 23949 26948
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 7524 26880 10640 26908
rect 12069 26911 12127 26917
rect 7524 26868 7530 26880
rect 12069 26877 12081 26911
rect 12115 26908 12127 26911
rect 12529 26911 12587 26917
rect 12529 26908 12541 26911
rect 12115 26880 12541 26908
rect 12115 26877 12127 26880
rect 12069 26871 12127 26877
rect 12529 26877 12541 26880
rect 12575 26908 12587 26911
rect 13630 26908 13636 26920
rect 12575 26880 13636 26908
rect 12575 26877 12587 26880
rect 12529 26871 12587 26877
rect 13630 26868 13636 26880
rect 13688 26868 13694 26920
rect 13906 26908 13912 26920
rect 13867 26880 13912 26908
rect 13906 26868 13912 26880
rect 13964 26868 13970 26920
rect 16298 26868 16304 26920
rect 16356 26908 16362 26920
rect 16669 26911 16727 26917
rect 16669 26908 16681 26911
rect 16356 26880 16681 26908
rect 16356 26868 16362 26880
rect 16669 26877 16681 26880
rect 16715 26877 16727 26911
rect 16669 26871 16727 26877
rect 16945 26911 17003 26917
rect 16945 26877 16957 26911
rect 16991 26908 17003 26911
rect 17862 26908 17868 26920
rect 16991 26880 17868 26908
rect 16991 26877 17003 26880
rect 16945 26871 17003 26877
rect 17862 26868 17868 26880
rect 17920 26868 17926 26920
rect 23952 26908 23980 26939
rect 24026 26936 24032 26988
rect 24084 26976 24090 26988
rect 24949 26979 25007 26985
rect 24949 26976 24961 26979
rect 24084 26948 24961 26976
rect 24084 26936 24090 26948
rect 24949 26945 24961 26948
rect 24995 26945 25007 26979
rect 25222 26976 25228 26988
rect 25183 26948 25228 26976
rect 24949 26939 25007 26945
rect 25222 26936 25228 26948
rect 25280 26936 25286 26988
rect 25774 26936 25780 26988
rect 25832 26985 25838 26988
rect 26169 26985 26197 27016
rect 26326 27004 26332 27016
rect 26384 27004 26390 27056
rect 26421 27047 26479 27053
rect 26421 27013 26433 27047
rect 26467 27044 26479 27047
rect 26467 27016 27384 27044
rect 26467 27013 26479 27016
rect 26421 27007 26479 27013
rect 25832 26976 25841 26985
rect 25940 26979 25998 26985
rect 25832 26948 25877 26976
rect 25832 26939 25841 26948
rect 25940 26945 25952 26979
rect 25986 26976 25998 26979
rect 26053 26979 26111 26985
rect 25986 26945 26004 26976
rect 25940 26939 26004 26945
rect 26053 26945 26065 26979
rect 26099 26945 26111 26979
rect 26053 26939 26111 26945
rect 26165 26979 26223 26985
rect 26165 26945 26177 26979
rect 26211 26945 26223 26979
rect 27356 26976 27384 27016
rect 27614 27004 27620 27056
rect 27672 27044 27678 27056
rect 28166 27044 28172 27056
rect 27672 27016 28172 27044
rect 27672 27004 27678 27016
rect 28166 27004 28172 27016
rect 28224 27044 28230 27056
rect 28997 27047 29055 27053
rect 28224 27016 28580 27044
rect 28224 27004 28230 27016
rect 28552 26985 28580 27016
rect 28997 27013 29009 27047
rect 29043 27044 29055 27047
rect 29086 27044 29092 27056
rect 29043 27016 29092 27044
rect 29043 27013 29055 27016
rect 28997 27007 29055 27013
rect 29086 27004 29092 27016
rect 29144 27044 29150 27056
rect 30009 27047 30067 27053
rect 30009 27044 30021 27047
rect 29144 27016 30021 27044
rect 29144 27004 29150 27016
rect 30009 27013 30021 27016
rect 30055 27044 30067 27047
rect 30834 27044 30840 27056
rect 30055 27016 30840 27044
rect 30055 27013 30067 27016
rect 30009 27007 30067 27013
rect 30834 27004 30840 27016
rect 30892 27004 30898 27056
rect 32122 27044 32128 27056
rect 31726 27016 32128 27044
rect 28270 26979 28328 26985
rect 28270 26976 28282 26979
rect 27356 26948 28282 26976
rect 26165 26939 26223 26945
rect 28270 26945 28282 26948
rect 28316 26945 28328 26979
rect 28270 26939 28328 26945
rect 28537 26979 28595 26985
rect 28537 26945 28549 26979
rect 28583 26945 28595 26979
rect 28537 26939 28595 26945
rect 29181 26979 29239 26985
rect 29181 26945 29193 26979
rect 29227 26976 29239 26979
rect 29914 26976 29920 26988
rect 29227 26948 29920 26976
rect 29227 26945 29239 26948
rect 29181 26939 29239 26945
rect 25832 26936 25838 26939
rect 24854 26908 24860 26920
rect 23952 26880 24860 26908
rect 24854 26868 24860 26880
rect 24912 26868 24918 26920
rect 9122 26840 9128 26852
rect 6840 26812 9128 26840
rect 9122 26800 9128 26812
rect 9180 26800 9186 26852
rect 9490 26800 9496 26852
rect 9548 26840 9554 26852
rect 11882 26840 11888 26852
rect 9548 26812 11888 26840
rect 9548 26800 9554 26812
rect 11882 26800 11888 26812
rect 11940 26800 11946 26852
rect 25976 26840 26004 26939
rect 26068 26908 26096 26939
rect 29914 26936 29920 26948
rect 29972 26936 29978 26988
rect 30193 26979 30251 26985
rect 30193 26945 30205 26979
rect 30239 26976 30251 26979
rect 31726 26976 31754 27016
rect 32122 27004 32128 27016
rect 32180 27004 32186 27056
rect 30239 26948 31754 26976
rect 30239 26945 30251 26948
rect 30193 26939 30251 26945
rect 26326 26908 26332 26920
rect 26068 26880 26332 26908
rect 26326 26868 26332 26880
rect 26384 26868 26390 26920
rect 29638 26868 29644 26920
rect 29696 26908 29702 26920
rect 30208 26908 30236 26939
rect 29696 26880 30236 26908
rect 29696 26868 29702 26880
rect 26602 26840 26608 26852
rect 25976 26812 26608 26840
rect 26602 26800 26608 26812
rect 26660 26800 26666 26852
rect 3694 26732 3700 26784
rect 3752 26772 3758 26784
rect 4801 26775 4859 26781
rect 4801 26772 4813 26775
rect 3752 26744 4813 26772
rect 3752 26732 3758 26744
rect 4801 26741 4813 26744
rect 4847 26772 4859 26775
rect 10410 26772 10416 26784
rect 4847 26744 10416 26772
rect 4847 26741 4859 26744
rect 4801 26735 4859 26741
rect 10410 26732 10416 26744
rect 10468 26732 10474 26784
rect 12894 26772 12900 26784
rect 12855 26744 12900 26772
rect 12894 26732 12900 26744
rect 12952 26732 12958 26784
rect 14921 26775 14979 26781
rect 14921 26741 14933 26775
rect 14967 26772 14979 26775
rect 15194 26772 15200 26784
rect 14967 26744 15200 26772
rect 14967 26741 14979 26744
rect 14921 26735 14979 26741
rect 15194 26732 15200 26744
rect 15252 26772 15258 26784
rect 16022 26772 16028 26784
rect 15252 26744 16028 26772
rect 15252 26732 15258 26744
rect 16022 26732 16028 26744
rect 16080 26732 16086 26784
rect 18046 26732 18052 26784
rect 18104 26772 18110 26784
rect 19242 26772 19248 26784
rect 18104 26744 19248 26772
rect 18104 26732 18110 26744
rect 19242 26732 19248 26744
rect 19300 26772 19306 26784
rect 19429 26775 19487 26781
rect 19429 26772 19441 26775
rect 19300 26744 19441 26772
rect 19300 26732 19306 26744
rect 19429 26741 19441 26744
rect 19475 26741 19487 26775
rect 19429 26735 19487 26741
rect 22189 26775 22247 26781
rect 22189 26741 22201 26775
rect 22235 26772 22247 26775
rect 22646 26772 22652 26784
rect 22235 26744 22652 26772
rect 22235 26741 22247 26744
rect 22189 26735 22247 26741
rect 22646 26732 22652 26744
rect 22704 26732 22710 26784
rect 23382 26732 23388 26784
rect 23440 26772 23446 26784
rect 23569 26775 23627 26781
rect 23569 26772 23581 26775
rect 23440 26744 23581 26772
rect 23440 26732 23446 26744
rect 23569 26741 23581 26744
rect 23615 26741 23627 26775
rect 23569 26735 23627 26741
rect 26418 26732 26424 26784
rect 26476 26772 26482 26784
rect 27157 26775 27215 26781
rect 27157 26772 27169 26775
rect 26476 26744 27169 26772
rect 26476 26732 26482 26744
rect 27157 26741 27169 26744
rect 27203 26741 27215 26775
rect 27157 26735 27215 26741
rect 30929 26775 30987 26781
rect 30929 26741 30941 26775
rect 30975 26772 30987 26775
rect 31018 26772 31024 26784
rect 30975 26744 31024 26772
rect 30975 26741 30987 26744
rect 30929 26735 30987 26741
rect 31018 26732 31024 26744
rect 31076 26732 31082 26784
rect 67634 26772 67640 26784
rect 67595 26744 67640 26772
rect 67634 26732 67640 26744
rect 67692 26732 67698 26784
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 2498 26528 2504 26580
rect 2556 26568 2562 26580
rect 2593 26571 2651 26577
rect 2593 26568 2605 26571
rect 2556 26540 2605 26568
rect 2556 26528 2562 26540
rect 2593 26537 2605 26540
rect 2639 26537 2651 26571
rect 5166 26568 5172 26580
rect 5079 26540 5172 26568
rect 2593 26531 2651 26537
rect 5166 26528 5172 26540
rect 5224 26568 5230 26580
rect 7466 26568 7472 26580
rect 5224 26540 7472 26568
rect 5224 26528 5230 26540
rect 7466 26528 7472 26540
rect 7524 26528 7530 26580
rect 8202 26568 8208 26580
rect 8163 26540 8208 26568
rect 8202 26528 8208 26540
rect 8260 26528 8266 26580
rect 12158 26528 12164 26580
rect 12216 26568 12222 26580
rect 12802 26568 12808 26580
rect 12216 26540 12808 26568
rect 12216 26528 12222 26540
rect 12802 26528 12808 26540
rect 12860 26528 12866 26580
rect 14090 26528 14096 26580
rect 14148 26568 14154 26580
rect 14185 26571 14243 26577
rect 14185 26568 14197 26571
rect 14148 26540 14197 26568
rect 14148 26528 14154 26540
rect 14185 26537 14197 26540
rect 14231 26537 14243 26571
rect 25774 26568 25780 26580
rect 14185 26531 14243 26537
rect 23216 26540 25780 26568
rect 3694 26500 3700 26512
rect 2424 26472 3700 26500
rect 2424 26373 2452 26472
rect 3694 26460 3700 26472
rect 3752 26460 3758 26512
rect 10781 26503 10839 26509
rect 10781 26469 10793 26503
rect 10827 26500 10839 26503
rect 11882 26500 11888 26512
rect 10827 26472 11888 26500
rect 10827 26469 10839 26472
rect 10781 26463 10839 26469
rect 11882 26460 11888 26472
rect 11940 26460 11946 26512
rect 12618 26500 12624 26512
rect 12406 26472 12624 26500
rect 3418 26392 3424 26444
rect 3476 26432 3482 26444
rect 3786 26432 3792 26444
rect 3476 26404 3792 26432
rect 3476 26392 3482 26404
rect 3786 26392 3792 26404
rect 3844 26392 3850 26444
rect 12406 26432 12434 26472
rect 12618 26460 12624 26472
rect 12676 26460 12682 26512
rect 13078 26460 13084 26512
rect 13136 26500 13142 26512
rect 18506 26500 18512 26512
rect 13136 26472 16620 26500
rect 13136 26460 13142 26472
rect 10244 26404 12434 26432
rect 2409 26367 2467 26373
rect 2409 26333 2421 26367
rect 2455 26333 2467 26367
rect 3804 26364 3832 26392
rect 6822 26364 6828 26376
rect 3804 26336 6828 26364
rect 2409 26327 2467 26333
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 10244 26373 10272 26404
rect 10229 26367 10287 26373
rect 10229 26333 10241 26367
rect 10275 26333 10287 26367
rect 10505 26367 10563 26373
rect 10505 26364 10517 26367
rect 10229 26327 10287 26333
rect 10336 26336 10517 26364
rect 1762 26256 1768 26308
rect 1820 26296 1826 26308
rect 2225 26299 2283 26305
rect 2225 26296 2237 26299
rect 1820 26268 2237 26296
rect 1820 26256 1826 26268
rect 2225 26265 2237 26268
rect 2271 26265 2283 26299
rect 2225 26259 2283 26265
rect 3234 26256 3240 26308
rect 3292 26296 3298 26308
rect 4034 26299 4092 26305
rect 4034 26296 4046 26299
rect 3292 26268 4046 26296
rect 3292 26256 3298 26268
rect 4034 26265 4046 26268
rect 4080 26265 4092 26299
rect 4034 26259 4092 26265
rect 6914 26256 6920 26308
rect 6972 26296 6978 26308
rect 7070 26299 7128 26305
rect 7070 26296 7082 26299
rect 6972 26268 7082 26296
rect 6972 26256 6978 26268
rect 7070 26265 7082 26268
rect 7116 26265 7128 26299
rect 10336 26296 10364 26336
rect 10505 26333 10517 26336
rect 10551 26333 10563 26367
rect 10505 26327 10563 26333
rect 10594 26324 10600 26376
rect 10652 26364 10658 26376
rect 12345 26367 12403 26373
rect 10652 26336 10697 26364
rect 10652 26324 10658 26336
rect 12345 26333 12357 26367
rect 12391 26333 12403 26367
rect 12345 26327 12403 26333
rect 12437 26367 12495 26373
rect 12437 26333 12449 26367
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 7070 26259 7128 26265
rect 7208 26268 10364 26296
rect 5718 26188 5724 26240
rect 5776 26228 5782 26240
rect 7208 26228 7236 26268
rect 10410 26256 10416 26308
rect 10468 26296 10474 26308
rect 10468 26268 10513 26296
rect 10468 26256 10474 26268
rect 10686 26256 10692 26308
rect 10744 26296 10750 26308
rect 12069 26299 12127 26305
rect 12069 26296 12081 26299
rect 10744 26268 12081 26296
rect 10744 26256 10750 26268
rect 12069 26265 12081 26268
rect 12115 26265 12127 26299
rect 12069 26259 12127 26265
rect 5776 26200 7236 26228
rect 12360 26228 12388 26327
rect 12452 26296 12480 26327
rect 12526 26324 12532 26376
rect 12584 26364 12590 26376
rect 12713 26367 12771 26373
rect 12584 26336 12629 26364
rect 12584 26324 12590 26336
rect 12713 26333 12725 26367
rect 12759 26364 12771 26367
rect 12802 26364 12808 26376
rect 12759 26336 12808 26364
rect 12759 26333 12771 26336
rect 12713 26327 12771 26333
rect 12802 26324 12808 26336
rect 12860 26324 12866 26376
rect 12894 26324 12900 26376
rect 12952 26364 12958 26376
rect 13173 26367 13231 26373
rect 13173 26364 13185 26367
rect 12952 26336 13185 26364
rect 12952 26324 12958 26336
rect 13173 26333 13185 26336
rect 13219 26333 13231 26367
rect 13173 26327 13231 26333
rect 13998 26324 14004 26376
rect 14056 26364 14062 26376
rect 14093 26367 14151 26373
rect 14093 26364 14105 26367
rect 14056 26336 14105 26364
rect 14056 26324 14062 26336
rect 14093 26333 14105 26336
rect 14139 26333 14151 26367
rect 14093 26327 14151 26333
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 14737 26367 14795 26373
rect 14737 26333 14749 26367
rect 14783 26364 14795 26367
rect 14918 26364 14924 26376
rect 14783 26336 14924 26364
rect 14783 26333 14795 26336
rect 14737 26327 14795 26333
rect 13906 26296 13912 26308
rect 12452 26268 13912 26296
rect 13906 26256 13912 26268
rect 13964 26256 13970 26308
rect 14292 26296 14320 26327
rect 14918 26324 14924 26336
rect 14976 26324 14982 26376
rect 15010 26324 15016 26376
rect 15068 26364 15074 26376
rect 16025 26367 16083 26373
rect 16025 26364 16037 26367
rect 15068 26336 16037 26364
rect 15068 26324 15074 26336
rect 16025 26333 16037 26336
rect 16071 26333 16083 26367
rect 16025 26327 16083 26333
rect 16209 26367 16267 26373
rect 16209 26333 16221 26367
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 16224 26296 16252 26327
rect 16482 26296 16488 26308
rect 14292 26268 16488 26296
rect 16482 26256 16488 26268
rect 16540 26256 16546 26308
rect 16592 26296 16620 26472
rect 17788 26472 18512 26500
rect 17788 26432 17816 26472
rect 18506 26460 18512 26472
rect 18564 26500 18570 26512
rect 20990 26500 20996 26512
rect 18564 26472 20024 26500
rect 20951 26472 20996 26500
rect 18564 26460 18570 26472
rect 17512 26404 17816 26432
rect 16758 26324 16764 26376
rect 16816 26364 16822 26376
rect 17512 26373 17540 26404
rect 17862 26392 17868 26444
rect 17920 26432 17926 26444
rect 19996 26441 20024 26472
rect 20990 26460 20996 26472
rect 21048 26460 21054 26512
rect 19981 26435 20039 26441
rect 17920 26404 18368 26432
rect 17920 26392 17926 26404
rect 17313 26367 17371 26373
rect 17313 26364 17325 26367
rect 16816 26336 17325 26364
rect 16816 26324 16822 26336
rect 17313 26333 17325 26336
rect 17359 26333 17371 26367
rect 17313 26327 17371 26333
rect 17497 26367 17555 26373
rect 17497 26333 17509 26367
rect 17543 26333 17555 26367
rect 17497 26327 17555 26333
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 18012 26336 18061 26364
rect 18012 26324 18018 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 18230 26364 18236 26376
rect 18191 26336 18236 26364
rect 18049 26327 18107 26333
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 18340 26373 18368 26404
rect 19981 26401 19993 26435
rect 20027 26401 20039 26435
rect 19981 26395 20039 26401
rect 22373 26435 22431 26441
rect 22373 26401 22385 26435
rect 22419 26432 22431 26435
rect 22830 26432 22836 26444
rect 22419 26404 22836 26432
rect 22419 26401 22431 26404
rect 22373 26395 22431 26401
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 18325 26367 18383 26373
rect 18325 26333 18337 26367
rect 18371 26333 18383 26367
rect 18325 26327 18383 26333
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26364 18475 26367
rect 19702 26364 19708 26376
rect 18463 26336 19564 26364
rect 19663 26336 19708 26364
rect 18463 26333 18475 26336
rect 18417 26327 18475 26333
rect 16853 26299 16911 26305
rect 16853 26296 16865 26299
rect 16592 26268 16865 26296
rect 16853 26265 16865 26268
rect 16899 26296 16911 26299
rect 18432 26296 18460 26327
rect 16899 26268 18460 26296
rect 18693 26299 18751 26305
rect 16899 26265 16911 26268
rect 16853 26259 16911 26265
rect 18693 26265 18705 26299
rect 18739 26296 18751 26299
rect 19334 26296 19340 26308
rect 18739 26268 19340 26296
rect 18739 26265 18751 26268
rect 18693 26259 18751 26265
rect 19334 26256 19340 26268
rect 19392 26256 19398 26308
rect 19536 26296 19564 26336
rect 19702 26324 19708 26336
rect 19760 26324 19766 26376
rect 22738 26324 22744 26376
rect 22796 26364 22802 26376
rect 23216 26373 23244 26540
rect 25774 26528 25780 26540
rect 25832 26528 25838 26580
rect 26602 26568 26608 26580
rect 26563 26540 26608 26568
rect 26602 26528 26608 26540
rect 26660 26528 26666 26580
rect 27706 26568 27712 26580
rect 27667 26540 27712 26568
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 23382 26460 23388 26512
rect 23440 26460 23446 26512
rect 24394 26500 24400 26512
rect 24355 26472 24400 26500
rect 24394 26460 24400 26472
rect 24452 26460 24458 26512
rect 26694 26460 26700 26512
rect 26752 26500 26758 26512
rect 28445 26503 28503 26509
rect 28445 26500 28457 26503
rect 26752 26472 28457 26500
rect 26752 26460 26758 26472
rect 28445 26469 28457 26472
rect 28491 26500 28503 26503
rect 28491 26472 31754 26500
rect 28491 26469 28503 26472
rect 28445 26463 28503 26469
rect 23400 26432 23428 26460
rect 23750 26432 23756 26444
rect 23395 26404 23428 26432
rect 23479 26404 23756 26432
rect 23201 26367 23259 26373
rect 23395 26370 23423 26404
rect 23479 26373 23507 26404
rect 23750 26392 23756 26404
rect 23808 26392 23814 26444
rect 25774 26432 25780 26444
rect 25735 26404 25780 26432
rect 25774 26392 25780 26404
rect 25832 26392 25838 26444
rect 27706 26392 27712 26444
rect 27764 26432 27770 26444
rect 27764 26404 30236 26432
rect 27764 26392 27770 26404
rect 23201 26364 23213 26367
rect 22796 26336 23213 26364
rect 22796 26324 22802 26336
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 23364 26364 23423 26370
rect 23364 26330 23376 26364
rect 23410 26333 23423 26364
rect 23464 26367 23522 26373
rect 23464 26333 23476 26367
rect 23510 26333 23522 26367
rect 23410 26330 23422 26333
rect 23364 26324 23422 26330
rect 23464 26327 23522 26333
rect 23566 26324 23572 26376
rect 23624 26373 23630 26376
rect 23624 26367 23647 26373
rect 23635 26333 23647 26367
rect 23624 26327 23647 26333
rect 23624 26324 23630 26327
rect 26050 26324 26056 26376
rect 26108 26364 26114 26376
rect 30208 26373 30236 26404
rect 30742 26392 30748 26444
rect 30800 26432 30806 26444
rect 30800 26404 30972 26432
rect 30800 26392 30806 26404
rect 28997 26367 29055 26373
rect 28997 26364 29009 26367
rect 26108 26336 29009 26364
rect 26108 26324 26114 26336
rect 28997 26333 29009 26336
rect 29043 26364 29055 26367
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 29043 26336 29837 26364
rect 29043 26333 29055 26336
rect 28997 26327 29055 26333
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26333 29975 26367
rect 29917 26327 29975 26333
rect 30009 26367 30067 26373
rect 30009 26333 30021 26367
rect 30055 26333 30067 26367
rect 30009 26327 30067 26333
rect 30193 26367 30251 26373
rect 30193 26333 30205 26367
rect 30239 26333 30251 26367
rect 30650 26364 30656 26376
rect 30611 26336 30656 26364
rect 30193 26327 30251 26333
rect 19536 26268 22048 26296
rect 12434 26228 12440 26240
rect 12360 26200 12440 26228
rect 5776 26188 5782 26200
rect 12434 26188 12440 26200
rect 12492 26188 12498 26240
rect 12618 26188 12624 26240
rect 12676 26228 12682 26240
rect 13357 26231 13415 26237
rect 13357 26228 13369 26231
rect 12676 26200 13369 26228
rect 12676 26188 12682 26200
rect 13357 26197 13369 26200
rect 13403 26197 13415 26231
rect 13357 26191 13415 26197
rect 16209 26231 16267 26237
rect 16209 26197 16221 26231
rect 16255 26228 16267 26231
rect 16298 26228 16304 26240
rect 16255 26200 16304 26228
rect 16255 26197 16267 26200
rect 16209 26191 16267 26197
rect 16298 26188 16304 26200
rect 16356 26188 16362 26240
rect 18782 26188 18788 26240
rect 18840 26228 18846 26240
rect 19702 26228 19708 26240
rect 18840 26200 19708 26228
rect 18840 26188 18846 26200
rect 19702 26188 19708 26200
rect 19760 26188 19766 26240
rect 22020 26228 22048 26268
rect 22094 26256 22100 26308
rect 22152 26305 22158 26308
rect 22152 26296 22164 26305
rect 23845 26299 23903 26305
rect 22152 26268 22197 26296
rect 22152 26259 22164 26268
rect 23845 26265 23857 26299
rect 23891 26296 23903 26299
rect 25510 26299 25568 26305
rect 25510 26296 25522 26299
rect 23891 26268 25522 26296
rect 23891 26265 23903 26268
rect 23845 26259 23903 26265
rect 25510 26265 25522 26268
rect 25556 26265 25568 26299
rect 25510 26259 25568 26265
rect 22152 26256 22158 26259
rect 26142 26256 26148 26308
rect 26200 26296 26206 26308
rect 26237 26299 26295 26305
rect 26237 26296 26249 26299
rect 26200 26268 26249 26296
rect 26200 26256 26206 26268
rect 26237 26265 26249 26268
rect 26283 26265 26295 26299
rect 26418 26296 26424 26308
rect 26379 26268 26424 26296
rect 26237 26259 26295 26265
rect 26418 26256 26424 26268
rect 26476 26256 26482 26308
rect 27062 26296 27068 26308
rect 27023 26268 27068 26296
rect 27062 26256 27068 26268
rect 27120 26296 27126 26308
rect 28261 26299 28319 26305
rect 28261 26296 28273 26299
rect 27120 26268 28273 26296
rect 27120 26256 27126 26268
rect 28261 26265 28273 26268
rect 28307 26265 28319 26299
rect 28261 26259 28319 26265
rect 29730 26256 29736 26308
rect 29788 26296 29794 26308
rect 29932 26296 29960 26327
rect 29788 26268 29960 26296
rect 30024 26296 30052 26327
rect 30650 26324 30656 26336
rect 30708 26324 30714 26376
rect 30834 26364 30840 26376
rect 30795 26336 30840 26364
rect 30834 26324 30840 26336
rect 30892 26324 30898 26376
rect 30944 26373 30972 26404
rect 30929 26367 30987 26373
rect 30929 26333 30941 26367
rect 30975 26333 30987 26367
rect 30929 26327 30987 26333
rect 31018 26324 31024 26376
rect 31076 26364 31082 26376
rect 31726 26364 31754 26472
rect 33137 26435 33195 26441
rect 33137 26401 33149 26435
rect 33183 26432 33195 26435
rect 33502 26432 33508 26444
rect 33183 26404 33508 26432
rect 33183 26401 33195 26404
rect 33137 26395 33195 26401
rect 33502 26392 33508 26404
rect 33560 26392 33566 26444
rect 34054 26364 34060 26376
rect 31076 26336 31121 26364
rect 31726 26336 34060 26364
rect 31076 26324 31082 26336
rect 34054 26324 34060 26336
rect 34112 26324 34118 26376
rect 31202 26296 31208 26308
rect 30024 26268 31208 26296
rect 29788 26256 29794 26268
rect 31202 26256 31208 26268
rect 31260 26256 31266 26308
rect 31297 26299 31355 26305
rect 31297 26265 31309 26299
rect 31343 26296 31355 26299
rect 32870 26299 32928 26305
rect 32870 26296 32882 26299
rect 31343 26268 32882 26296
rect 31343 26265 31355 26268
rect 31297 26259 31355 26265
rect 32870 26265 32882 26268
rect 32916 26265 32928 26299
rect 32870 26259 32928 26265
rect 24762 26228 24768 26240
rect 22020 26200 24768 26228
rect 24762 26188 24768 26200
rect 24820 26188 24826 26240
rect 29546 26228 29552 26240
rect 29507 26200 29552 26228
rect 29546 26188 29552 26200
rect 29604 26188 29610 26240
rect 31757 26231 31815 26237
rect 31757 26197 31769 26231
rect 31803 26228 31815 26231
rect 31846 26228 31852 26240
rect 31803 26200 31852 26228
rect 31803 26197 31815 26200
rect 31757 26191 31815 26197
rect 31846 26188 31852 26200
rect 31904 26188 31910 26240
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 3234 26024 3240 26036
rect 3195 25996 3240 26024
rect 3234 25984 3240 25996
rect 3292 25984 3298 26036
rect 6822 25984 6828 26036
rect 6880 25984 6886 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 12897 26027 12955 26033
rect 12897 26024 12909 26027
rect 12492 25996 12909 26024
rect 12492 25984 12498 25996
rect 12897 25993 12909 25996
rect 12943 26024 12955 26027
rect 13078 26024 13084 26036
rect 12943 25996 13084 26024
rect 12943 25993 12955 25996
rect 12897 25987 12955 25993
rect 13078 25984 13084 25996
rect 13136 25984 13142 26036
rect 15930 25984 15936 26036
rect 15988 25984 15994 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 22189 26027 22247 26033
rect 22189 26024 22201 26027
rect 22152 25996 22201 26024
rect 22152 25984 22158 25996
rect 22189 25993 22201 25996
rect 22235 25993 22247 26027
rect 22189 25987 22247 25993
rect 25774 25984 25780 26036
rect 25832 26024 25838 26036
rect 25961 26027 26019 26033
rect 25961 26024 25973 26027
rect 25832 25996 25973 26024
rect 25832 25984 25838 25996
rect 25961 25993 25973 25996
rect 26007 26024 26019 26027
rect 27798 26024 27804 26036
rect 26007 25996 27804 26024
rect 26007 25993 26019 25996
rect 25961 25987 26019 25993
rect 27798 25984 27804 25996
rect 27856 25984 27862 26036
rect 30834 25984 30840 26036
rect 30892 26024 30898 26036
rect 31481 26027 31539 26033
rect 31481 26024 31493 26027
rect 30892 25996 31493 26024
rect 30892 25984 30898 25996
rect 31481 25993 31493 25996
rect 31527 25993 31539 26027
rect 31481 25987 31539 25993
rect 33502 25984 33508 26036
rect 33560 26024 33566 26036
rect 34422 26024 34428 26036
rect 33560 25996 34428 26024
rect 33560 25984 33566 25996
rect 34422 25984 34428 25996
rect 34480 26024 34486 26036
rect 34885 26027 34943 26033
rect 34885 26024 34897 26027
rect 34480 25996 34897 26024
rect 34480 25984 34486 25996
rect 34885 25993 34897 25996
rect 34931 25993 34943 26027
rect 34885 25987 34943 25993
rect 1762 25956 1768 25968
rect 1723 25928 1768 25956
rect 1762 25916 1768 25928
rect 1820 25916 1826 25968
rect 1949 25959 2007 25965
rect 1949 25925 1961 25959
rect 1995 25956 2007 25959
rect 5166 25956 5172 25968
rect 1995 25928 5172 25956
rect 1995 25925 2007 25928
rect 1949 25919 2007 25925
rect 5166 25916 5172 25928
rect 5224 25916 5230 25968
rect 6840 25956 6868 25984
rect 8472 25959 8530 25965
rect 6840 25928 8248 25956
rect 2314 25848 2320 25900
rect 2372 25888 2378 25900
rect 2593 25891 2651 25897
rect 2593 25888 2605 25891
rect 2372 25860 2605 25888
rect 2372 25848 2378 25860
rect 2593 25857 2605 25860
rect 2639 25857 2651 25891
rect 2593 25851 2651 25857
rect 2777 25891 2835 25897
rect 2777 25857 2789 25891
rect 2823 25857 2835 25891
rect 2777 25851 2835 25857
rect 2133 25823 2191 25829
rect 2133 25789 2145 25823
rect 2179 25820 2191 25823
rect 2792 25820 2820 25851
rect 2866 25848 2872 25900
rect 2924 25888 2930 25900
rect 3007 25891 3065 25897
rect 2924 25860 2969 25888
rect 2924 25848 2930 25860
rect 3007 25857 3019 25891
rect 3053 25888 3065 25891
rect 3789 25891 3847 25897
rect 3789 25888 3801 25891
rect 3053 25860 3801 25888
rect 3053 25857 3065 25860
rect 3007 25851 3065 25857
rect 3789 25857 3801 25860
rect 3835 25888 3847 25891
rect 5813 25891 5871 25897
rect 5813 25888 5825 25891
rect 3835 25860 5825 25888
rect 3835 25857 3847 25860
rect 3789 25851 3847 25857
rect 5813 25857 5825 25860
rect 5859 25888 5871 25891
rect 6638 25888 6644 25900
rect 5859 25860 6644 25888
rect 5859 25857 5871 25860
rect 5813 25851 5871 25857
rect 6638 25848 6644 25860
rect 6696 25848 6702 25900
rect 6733 25891 6791 25897
rect 6733 25857 6745 25891
rect 6779 25857 6791 25891
rect 6733 25851 6791 25857
rect 2179 25792 2820 25820
rect 6748 25820 6776 25851
rect 6822 25848 6828 25900
rect 6880 25888 6886 25900
rect 6880 25860 6925 25888
rect 6880 25848 6886 25860
rect 7006 25848 7012 25900
rect 7064 25888 7070 25900
rect 7742 25888 7748 25900
rect 7064 25860 7748 25888
rect 7064 25848 7070 25860
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 8220 25897 8248 25928
rect 8472 25925 8484 25959
rect 8518 25956 8530 25959
rect 10686 25956 10692 25968
rect 8518 25928 10692 25956
rect 8518 25925 8530 25928
rect 8472 25919 8530 25925
rect 10686 25916 10692 25928
rect 10744 25916 10750 25968
rect 11517 25959 11575 25965
rect 11517 25925 11529 25959
rect 11563 25956 11575 25959
rect 15197 25959 15255 25965
rect 11563 25928 12020 25956
rect 11563 25925 11575 25928
rect 11517 25919 11575 25925
rect 8205 25891 8263 25897
rect 8205 25857 8217 25891
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11992 25888 12020 25928
rect 15197 25925 15209 25959
rect 15243 25956 15255 25959
rect 15749 25959 15807 25965
rect 15749 25956 15761 25959
rect 15243 25928 15761 25956
rect 15243 25925 15255 25928
rect 15197 25919 15255 25925
rect 15749 25925 15761 25928
rect 15795 25956 15807 25959
rect 15948 25956 15976 25984
rect 15795 25928 15976 25956
rect 15795 25925 15807 25928
rect 15749 25919 15807 25925
rect 16022 25916 16028 25968
rect 16080 25956 16086 25968
rect 16850 25956 16856 25968
rect 16080 25928 16856 25956
rect 16080 25916 16086 25928
rect 16850 25916 16856 25928
rect 16908 25956 16914 25968
rect 28074 25956 28080 25968
rect 16908 25928 21312 25956
rect 16908 25916 16914 25928
rect 12618 25888 12624 25900
rect 11992 25860 12624 25888
rect 11701 25851 11759 25857
rect 7374 25820 7380 25832
rect 6748 25792 7380 25820
rect 2179 25789 2191 25792
rect 2133 25783 2191 25789
rect 7374 25780 7380 25792
rect 7432 25780 7438 25832
rect 9585 25755 9643 25761
rect 9585 25721 9597 25755
rect 9631 25752 9643 25755
rect 10226 25752 10232 25764
rect 9631 25724 10232 25752
rect 9631 25721 9643 25724
rect 9585 25715 9643 25721
rect 10226 25712 10232 25724
rect 10284 25752 10290 25764
rect 11716 25752 11744 25851
rect 12618 25848 12624 25860
rect 12676 25848 12682 25900
rect 13817 25891 13875 25897
rect 13817 25857 13829 25891
rect 13863 25888 13875 25891
rect 13998 25888 14004 25900
rect 13863 25860 14004 25888
rect 13863 25857 13875 25860
rect 13817 25851 13875 25857
rect 13998 25848 14004 25860
rect 14056 25848 14062 25900
rect 15010 25888 15016 25900
rect 14971 25860 15016 25888
rect 15010 25848 15016 25860
rect 15068 25848 15074 25900
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25857 15991 25891
rect 15933 25851 15991 25857
rect 11885 25823 11943 25829
rect 11885 25789 11897 25823
rect 11931 25820 11943 25823
rect 12526 25820 12532 25832
rect 11931 25792 12532 25820
rect 11931 25789 11943 25792
rect 11885 25783 11943 25789
rect 12526 25780 12532 25792
rect 12584 25780 12590 25832
rect 12986 25780 12992 25832
rect 13044 25820 13050 25832
rect 13541 25823 13599 25829
rect 13541 25820 13553 25823
rect 13044 25792 13553 25820
rect 13044 25780 13050 25792
rect 13541 25789 13553 25792
rect 13587 25789 13599 25823
rect 14826 25820 14832 25832
rect 14787 25792 14832 25820
rect 13541 25783 13599 25789
rect 14826 25780 14832 25792
rect 14884 25780 14890 25832
rect 10284 25724 11744 25752
rect 10284 25712 10290 25724
rect 13998 25712 14004 25764
rect 14056 25752 14062 25764
rect 15948 25752 15976 25851
rect 16666 25848 16672 25900
rect 16724 25888 16730 25900
rect 18334 25891 18392 25897
rect 18334 25888 18346 25891
rect 16724 25860 18346 25888
rect 16724 25848 16730 25860
rect 18334 25857 18346 25860
rect 18380 25857 18392 25891
rect 18334 25851 18392 25857
rect 19334 25848 19340 25900
rect 19392 25888 19398 25900
rect 21284 25897 21312 25928
rect 22848 25928 28080 25956
rect 19501 25891 19559 25897
rect 19501 25888 19513 25891
rect 19392 25860 19513 25888
rect 19392 25848 19398 25860
rect 19501 25857 19513 25860
rect 19547 25857 19559 25891
rect 19501 25851 19559 25857
rect 21269 25891 21327 25897
rect 21269 25857 21281 25891
rect 21315 25888 21327 25891
rect 22462 25888 22468 25900
rect 21315 25860 22468 25888
rect 21315 25857 21327 25860
rect 21269 25851 21327 25857
rect 22462 25848 22468 25860
rect 22520 25848 22526 25900
rect 22557 25891 22615 25897
rect 22557 25857 22569 25891
rect 22603 25857 22615 25891
rect 22557 25851 22615 25857
rect 18601 25823 18659 25829
rect 18601 25789 18613 25823
rect 18647 25820 18659 25823
rect 19242 25820 19248 25832
rect 18647 25792 19248 25820
rect 18647 25789 18659 25792
rect 18601 25783 18659 25789
rect 19242 25780 19248 25792
rect 19300 25780 19306 25832
rect 22002 25780 22008 25832
rect 22060 25820 22066 25832
rect 22572 25820 22600 25851
rect 22646 25848 22652 25900
rect 22704 25888 22710 25900
rect 22848 25897 22876 25928
rect 28074 25916 28080 25928
rect 28132 25916 28138 25968
rect 29546 25965 29552 25968
rect 29540 25956 29552 25965
rect 29507 25928 29552 25956
rect 29540 25919 29552 25928
rect 29546 25916 29552 25919
rect 29604 25916 29610 25968
rect 30668 25928 32536 25956
rect 30668 25900 30696 25928
rect 32508 25900 32536 25928
rect 22833 25891 22891 25897
rect 22704 25860 22749 25888
rect 22704 25848 22710 25860
rect 22833 25857 22845 25891
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23569 25891 23627 25897
rect 23569 25857 23581 25891
rect 23615 25888 23627 25891
rect 23750 25888 23756 25900
rect 23615 25860 23756 25888
rect 23615 25857 23627 25860
rect 23569 25851 23627 25857
rect 23750 25848 23756 25860
rect 23808 25848 23814 25900
rect 24673 25891 24731 25897
rect 24673 25857 24685 25891
rect 24719 25888 24731 25891
rect 26234 25888 26240 25900
rect 24719 25860 26240 25888
rect 24719 25857 24731 25860
rect 24673 25851 24731 25857
rect 26234 25848 26240 25860
rect 26292 25888 26298 25900
rect 27982 25888 27988 25900
rect 26292 25860 27108 25888
rect 27943 25860 27988 25888
rect 26292 25848 26298 25860
rect 23290 25820 23296 25832
rect 22060 25792 22600 25820
rect 23251 25792 23296 25820
rect 22060 25780 22066 25792
rect 23290 25780 23296 25792
rect 23348 25780 23354 25832
rect 17221 25755 17279 25761
rect 17221 25752 17233 25755
rect 14056 25724 17233 25752
rect 14056 25712 14062 25724
rect 17221 25721 17233 25724
rect 17267 25721 17279 25755
rect 17221 25715 17279 25721
rect 6365 25687 6423 25693
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 6914 25684 6920 25696
rect 6411 25656 6920 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 6914 25644 6920 25656
rect 6972 25644 6978 25696
rect 16117 25687 16175 25693
rect 16117 25653 16129 25687
rect 16163 25684 16175 25687
rect 16206 25684 16212 25696
rect 16163 25656 16212 25684
rect 16163 25653 16175 25656
rect 16117 25647 16175 25653
rect 16206 25644 16212 25656
rect 16264 25644 16270 25696
rect 16390 25644 16396 25696
rect 16448 25684 16454 25696
rect 19426 25684 19432 25696
rect 16448 25656 19432 25684
rect 16448 25644 16454 25656
rect 19426 25644 19432 25656
rect 19484 25684 19490 25696
rect 27080 25693 27108 25860
rect 27982 25848 27988 25860
rect 28040 25848 28046 25900
rect 28166 25848 28172 25900
rect 28224 25888 28230 25900
rect 29273 25891 29331 25897
rect 29273 25888 29285 25891
rect 28224 25860 29285 25888
rect 28224 25848 28230 25860
rect 29273 25857 29285 25860
rect 29319 25857 29331 25891
rect 30650 25888 30656 25900
rect 29273 25851 29331 25857
rect 29380 25860 30656 25888
rect 28261 25823 28319 25829
rect 28261 25789 28273 25823
rect 28307 25820 28319 25823
rect 29380 25820 29408 25860
rect 30650 25848 30656 25860
rect 30708 25848 30714 25900
rect 30926 25848 30932 25900
rect 30984 25888 30990 25900
rect 31113 25891 31171 25897
rect 31113 25888 31125 25891
rect 30984 25860 31125 25888
rect 30984 25848 30990 25860
rect 31113 25857 31125 25860
rect 31159 25857 31171 25891
rect 31113 25851 31171 25857
rect 31297 25891 31355 25897
rect 31297 25857 31309 25891
rect 31343 25888 31355 25891
rect 31846 25888 31852 25900
rect 31343 25860 31852 25888
rect 31343 25857 31355 25860
rect 31297 25851 31355 25857
rect 31846 25848 31852 25860
rect 31904 25848 31910 25900
rect 32490 25888 32496 25900
rect 32403 25860 32496 25888
rect 32490 25848 32496 25860
rect 32548 25848 32554 25900
rect 32674 25888 32680 25900
rect 32635 25860 32680 25888
rect 32674 25848 32680 25860
rect 32732 25848 32738 25900
rect 32769 25891 32827 25897
rect 32769 25857 32781 25891
rect 32815 25857 32827 25891
rect 32769 25851 32827 25857
rect 28307 25792 29408 25820
rect 32784 25820 32812 25851
rect 32858 25848 32864 25900
rect 32916 25888 32922 25900
rect 33597 25891 33655 25897
rect 32916 25860 32961 25888
rect 32916 25848 32922 25860
rect 33597 25857 33609 25891
rect 33643 25888 33655 25891
rect 34698 25888 34704 25900
rect 33643 25860 34704 25888
rect 33643 25857 33655 25860
rect 33597 25851 33655 25857
rect 32950 25820 32956 25832
rect 32784 25792 32956 25820
rect 28307 25789 28319 25792
rect 28261 25783 28319 25789
rect 32950 25780 32956 25792
rect 33008 25780 33014 25832
rect 33612 25752 33640 25851
rect 34698 25848 34704 25860
rect 34756 25848 34762 25900
rect 30208 25724 33640 25752
rect 20625 25687 20683 25693
rect 20625 25684 20637 25687
rect 19484 25656 20637 25684
rect 19484 25644 19490 25656
rect 20625 25653 20637 25656
rect 20671 25653 20683 25687
rect 20625 25647 20683 25653
rect 27065 25687 27123 25693
rect 27065 25653 27077 25687
rect 27111 25684 27123 25687
rect 30208 25684 30236 25724
rect 27111 25656 30236 25684
rect 30653 25687 30711 25693
rect 27111 25653 27123 25656
rect 27065 25647 27123 25653
rect 30653 25653 30665 25687
rect 30699 25684 30711 25687
rect 31570 25684 31576 25696
rect 30699 25656 31576 25684
rect 30699 25653 30711 25656
rect 30653 25647 30711 25653
rect 31570 25644 31576 25656
rect 31628 25644 31634 25696
rect 33134 25684 33140 25696
rect 33095 25656 33140 25684
rect 33134 25644 33140 25656
rect 33192 25644 33198 25696
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 5718 25480 5724 25492
rect 5679 25452 5724 25480
rect 5718 25440 5724 25452
rect 5776 25440 5782 25492
rect 6733 25483 6791 25489
rect 6733 25449 6745 25483
rect 6779 25480 6791 25483
rect 6822 25480 6828 25492
rect 6779 25452 6828 25480
rect 6779 25449 6791 25452
rect 6733 25443 6791 25449
rect 6822 25440 6828 25452
rect 6880 25440 6886 25492
rect 16666 25480 16672 25492
rect 16627 25452 16672 25480
rect 16666 25440 16672 25452
rect 16724 25440 16730 25492
rect 20625 25483 20683 25489
rect 20625 25480 20637 25483
rect 19168 25452 20637 25480
rect 12250 25372 12256 25424
rect 12308 25412 12314 25424
rect 18598 25412 18604 25424
rect 12308 25384 18604 25412
rect 12308 25372 12314 25384
rect 18598 25372 18604 25384
rect 18656 25372 18662 25424
rect 18693 25415 18751 25421
rect 18693 25381 18705 25415
rect 18739 25412 18751 25415
rect 18782 25412 18788 25424
rect 18739 25384 18788 25412
rect 18739 25381 18751 25384
rect 18693 25375 18751 25381
rect 18782 25372 18788 25384
rect 18840 25412 18846 25424
rect 19058 25412 19064 25424
rect 18840 25384 19064 25412
rect 18840 25372 18846 25384
rect 19058 25372 19064 25384
rect 19116 25372 19122 25424
rect 3786 25304 3792 25356
rect 3844 25344 3850 25356
rect 4341 25347 4399 25353
rect 4341 25344 4353 25347
rect 3844 25316 4353 25344
rect 3844 25304 3850 25316
rect 4341 25313 4353 25316
rect 4387 25313 4399 25347
rect 10502 25344 10508 25356
rect 10463 25316 10508 25344
rect 4341 25307 4399 25313
rect 10502 25304 10508 25316
rect 10560 25304 10566 25356
rect 11698 25304 11704 25356
rect 11756 25344 11762 25356
rect 19168 25344 19196 25452
rect 20625 25449 20637 25452
rect 20671 25449 20683 25483
rect 20625 25443 20683 25449
rect 21913 25483 21971 25489
rect 21913 25449 21925 25483
rect 21959 25480 21971 25483
rect 23198 25480 23204 25492
rect 21959 25452 23204 25480
rect 21959 25449 21971 25452
rect 21913 25443 21971 25449
rect 23198 25440 23204 25452
rect 23256 25440 23262 25492
rect 31202 25440 31208 25492
rect 31260 25480 31266 25492
rect 31297 25483 31355 25489
rect 31297 25480 31309 25483
rect 31260 25452 31309 25480
rect 31260 25440 31266 25452
rect 31297 25449 31309 25452
rect 31343 25449 31355 25483
rect 31297 25443 31355 25449
rect 32674 25440 32680 25492
rect 32732 25480 32738 25492
rect 32769 25483 32827 25489
rect 32769 25480 32781 25483
rect 32732 25452 32781 25480
rect 32732 25440 32738 25452
rect 32769 25449 32781 25452
rect 32815 25449 32827 25483
rect 32769 25443 32827 25449
rect 20898 25372 20904 25424
rect 20956 25412 20962 25424
rect 26234 25412 26240 25424
rect 20956 25384 26240 25412
rect 20956 25372 20962 25384
rect 26234 25372 26240 25384
rect 26292 25372 26298 25424
rect 26789 25415 26847 25421
rect 26789 25381 26801 25415
rect 26835 25381 26847 25415
rect 26789 25375 26847 25381
rect 23658 25344 23664 25356
rect 11756 25316 19196 25344
rect 22388 25316 23664 25344
rect 11756 25304 11762 25316
rect 2314 25236 2320 25288
rect 2372 25276 2378 25288
rect 2593 25279 2651 25285
rect 2593 25276 2605 25279
rect 2372 25248 2605 25276
rect 2372 25236 2378 25248
rect 2593 25245 2605 25248
rect 2639 25245 2651 25279
rect 2593 25239 2651 25245
rect 2777 25279 2835 25285
rect 2777 25245 2789 25279
rect 2823 25245 2835 25279
rect 2777 25239 2835 25245
rect 2792 25140 2820 25239
rect 2866 25236 2872 25288
rect 2924 25276 2930 25288
rect 3007 25279 3065 25285
rect 2924 25248 2969 25276
rect 2924 25236 2930 25248
rect 3007 25245 3019 25279
rect 3053 25276 3065 25279
rect 3881 25279 3939 25285
rect 3881 25276 3893 25279
rect 3053 25248 3893 25276
rect 3053 25245 3065 25248
rect 3007 25239 3065 25245
rect 3881 25245 3893 25248
rect 3927 25276 3939 25279
rect 5626 25276 5632 25288
rect 3927 25248 5632 25276
rect 3927 25245 3939 25248
rect 3881 25239 3939 25245
rect 5626 25236 5632 25248
rect 5684 25236 5690 25288
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 8202 25276 8208 25288
rect 6963 25248 8208 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 8202 25236 8208 25248
rect 8260 25236 8266 25288
rect 14277 25279 14335 25285
rect 14277 25245 14289 25279
rect 14323 25276 14335 25279
rect 14458 25276 14464 25288
rect 14323 25248 14464 25276
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 16025 25279 16083 25285
rect 16025 25245 16037 25279
rect 16071 25245 16083 25279
rect 16206 25276 16212 25288
rect 16167 25248 16212 25276
rect 16025 25239 16083 25245
rect 3237 25211 3295 25217
rect 3237 25177 3249 25211
rect 3283 25208 3295 25211
rect 4586 25211 4644 25217
rect 4586 25208 4598 25211
rect 3283 25180 4598 25208
rect 3283 25177 3295 25180
rect 3237 25171 3295 25177
rect 4586 25177 4598 25180
rect 4632 25177 4644 25211
rect 7098 25208 7104 25220
rect 7059 25180 7104 25208
rect 4586 25171 4644 25177
rect 7098 25168 7104 25180
rect 7156 25168 7162 25220
rect 10772 25211 10830 25217
rect 10772 25177 10784 25211
rect 10818 25208 10830 25211
rect 12342 25208 12348 25220
rect 10818 25180 12348 25208
rect 10818 25177 10830 25180
rect 10772 25171 10830 25177
rect 12342 25168 12348 25180
rect 12400 25168 12406 25220
rect 12618 25168 12624 25220
rect 12676 25208 12682 25220
rect 14093 25211 14151 25217
rect 14093 25208 14105 25211
rect 12676 25180 14105 25208
rect 12676 25168 12682 25180
rect 14093 25177 14105 25180
rect 14139 25177 14151 25211
rect 14826 25208 14832 25220
rect 14093 25171 14151 25177
rect 14200 25180 14832 25208
rect 2866 25140 2872 25152
rect 2792 25112 2872 25140
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 11885 25143 11943 25149
rect 11885 25109 11897 25143
rect 11931 25140 11943 25143
rect 12434 25140 12440 25152
rect 11931 25112 12440 25140
rect 11931 25109 11943 25112
rect 11885 25103 11943 25109
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 13446 25140 13452 25152
rect 13407 25112 13452 25140
rect 13446 25100 13452 25112
rect 13504 25100 13510 25152
rect 13814 25100 13820 25152
rect 13872 25140 13878 25152
rect 14200 25140 14228 25180
rect 14826 25168 14832 25180
rect 14884 25208 14890 25220
rect 14921 25211 14979 25217
rect 14921 25208 14933 25211
rect 14884 25180 14933 25208
rect 14884 25168 14890 25180
rect 14921 25177 14933 25180
rect 14967 25177 14979 25211
rect 16040 25208 16068 25239
rect 16206 25236 16212 25248
rect 16264 25236 16270 25288
rect 16298 25236 16304 25288
rect 16356 25276 16362 25288
rect 16439 25279 16497 25285
rect 16356 25248 16401 25276
rect 16356 25236 16362 25248
rect 16439 25245 16451 25279
rect 16485 25276 16497 25279
rect 16850 25276 16856 25288
rect 16485 25248 16856 25276
rect 16485 25245 16497 25248
rect 16439 25239 16497 25245
rect 16850 25236 16856 25248
rect 16908 25236 16914 25288
rect 17586 25276 17592 25288
rect 17547 25248 17592 25276
rect 17586 25236 17592 25248
rect 17644 25236 17650 25288
rect 17788 25285 17816 25316
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25245 17831 25279
rect 19242 25276 19248 25288
rect 19203 25248 19248 25276
rect 17773 25239 17831 25245
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25276 21787 25279
rect 21910 25276 21916 25288
rect 21775 25248 21916 25276
rect 21775 25245 21787 25248
rect 21729 25239 21787 25245
rect 21910 25236 21916 25248
rect 21968 25236 21974 25288
rect 22388 25285 22416 25316
rect 23658 25304 23664 25316
rect 23716 25304 23722 25356
rect 26050 25344 26056 25356
rect 23768 25316 26056 25344
rect 22373 25279 22431 25285
rect 22373 25245 22385 25279
rect 22419 25245 22431 25279
rect 22554 25276 22560 25288
rect 22515 25248 22560 25276
rect 22373 25239 22431 25245
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 22646 25236 22652 25288
rect 22704 25276 22710 25288
rect 22787 25279 22845 25285
rect 22704 25248 22749 25276
rect 22704 25236 22710 25248
rect 22787 25245 22799 25279
rect 22833 25276 22845 25279
rect 23768 25276 23796 25316
rect 26050 25304 26056 25316
rect 26108 25304 26114 25356
rect 22833 25248 23796 25276
rect 22833 25245 22845 25248
rect 22787 25239 22845 25245
rect 16758 25208 16764 25220
rect 16040 25180 16764 25208
rect 14921 25171 14979 25177
rect 16758 25168 16764 25180
rect 16816 25168 16822 25220
rect 19334 25168 19340 25220
rect 19392 25208 19398 25220
rect 19490 25211 19548 25217
rect 19490 25208 19502 25211
rect 19392 25180 19502 25208
rect 19392 25168 19398 25180
rect 19490 25177 19502 25180
rect 19536 25177 19548 25211
rect 19490 25171 19548 25177
rect 20530 25168 20536 25220
rect 20588 25208 20594 25220
rect 21269 25211 21327 25217
rect 21269 25208 21281 25211
rect 20588 25180 21281 25208
rect 20588 25168 20594 25180
rect 21269 25177 21281 25180
rect 21315 25208 21327 25211
rect 22802 25208 22830 25239
rect 25222 25236 25228 25288
rect 25280 25276 25286 25288
rect 25501 25279 25559 25285
rect 25501 25276 25513 25279
rect 25280 25248 25513 25276
rect 25280 25236 25286 25248
rect 25501 25245 25513 25248
rect 25547 25245 25559 25279
rect 25501 25239 25559 25245
rect 25682 25236 25688 25288
rect 25740 25276 25746 25288
rect 25777 25279 25835 25285
rect 25777 25276 25789 25279
rect 25740 25248 25789 25276
rect 25740 25236 25746 25248
rect 25777 25245 25789 25248
rect 25823 25245 25835 25279
rect 26804 25276 26832 25375
rect 28166 25344 28172 25356
rect 28127 25316 28172 25344
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 29825 25347 29883 25353
rect 29825 25313 29837 25347
rect 29871 25344 29883 25347
rect 30742 25344 30748 25356
rect 29871 25316 30748 25344
rect 29871 25313 29883 25316
rect 29825 25307 29883 25313
rect 30742 25304 30748 25316
rect 30800 25304 30806 25356
rect 34422 25304 34428 25356
rect 34480 25344 34486 25356
rect 35437 25347 35495 25353
rect 35437 25344 35449 25347
rect 34480 25316 35449 25344
rect 34480 25304 34486 25316
rect 35437 25313 35449 25316
rect 35483 25313 35495 25347
rect 35437 25307 35495 25313
rect 29546 25276 29552 25288
rect 25777 25239 25835 25245
rect 25864 25248 26832 25276
rect 29507 25248 29552 25276
rect 23474 25208 23480 25220
rect 21315 25180 22830 25208
rect 23435 25180 23480 25208
rect 21315 25177 21327 25180
rect 21269 25171 21327 25177
rect 23474 25168 23480 25180
rect 23532 25168 23538 25220
rect 23661 25211 23719 25217
rect 23661 25177 23673 25211
rect 23707 25208 23719 25211
rect 24026 25208 24032 25220
rect 23707 25180 24032 25208
rect 23707 25177 23719 25180
rect 23661 25171 23719 25177
rect 24026 25168 24032 25180
rect 24084 25208 24090 25220
rect 25864 25208 25892 25248
rect 29546 25236 29552 25248
rect 29604 25236 29610 25288
rect 31665 25279 31723 25285
rect 31665 25245 31677 25279
rect 31711 25276 31723 25279
rect 31711 25248 31800 25276
rect 31711 25245 31723 25248
rect 31665 25239 31723 25245
rect 31772 25220 31800 25248
rect 33134 25236 33140 25288
rect 33192 25276 33198 25288
rect 35693 25279 35751 25285
rect 35693 25276 35705 25279
rect 33192 25248 35705 25276
rect 33192 25236 33198 25248
rect 35693 25245 35705 25248
rect 35739 25245 35751 25279
rect 68094 25276 68100 25288
rect 68055 25248 68100 25276
rect 35693 25239 35751 25245
rect 68094 25236 68100 25248
rect 68152 25236 68158 25288
rect 24084 25180 25892 25208
rect 24084 25168 24090 25180
rect 26326 25168 26332 25220
rect 26384 25208 26390 25220
rect 27902 25211 27960 25217
rect 27902 25208 27914 25211
rect 26384 25180 27914 25208
rect 26384 25168 26390 25180
rect 27902 25177 27914 25180
rect 27948 25177 27960 25211
rect 27902 25171 27960 25177
rect 31481 25211 31539 25217
rect 31481 25177 31493 25211
rect 31527 25208 31539 25211
rect 31570 25208 31576 25220
rect 31527 25180 31576 25208
rect 31527 25177 31539 25180
rect 31481 25171 31539 25177
rect 31570 25168 31576 25180
rect 31628 25168 31634 25220
rect 31754 25168 31760 25220
rect 31812 25208 31818 25220
rect 32401 25211 32459 25217
rect 32401 25208 32413 25211
rect 31812 25180 32413 25208
rect 31812 25168 31818 25180
rect 32401 25177 32413 25180
rect 32447 25177 32459 25211
rect 32401 25171 32459 25177
rect 32585 25211 32643 25217
rect 32585 25177 32597 25211
rect 32631 25208 32643 25211
rect 32674 25208 32680 25220
rect 32631 25180 32680 25208
rect 32631 25177 32643 25180
rect 32585 25171 32643 25177
rect 32674 25168 32680 25180
rect 32732 25208 32738 25220
rect 32732 25180 36860 25208
rect 32732 25168 32738 25180
rect 13872 25112 14228 25140
rect 13872 25100 13878 25112
rect 14366 25100 14372 25152
rect 14424 25140 14430 25152
rect 14461 25143 14519 25149
rect 14461 25140 14473 25143
rect 14424 25112 14473 25140
rect 14424 25100 14430 25112
rect 14461 25109 14473 25112
rect 14507 25109 14519 25143
rect 14461 25103 14519 25109
rect 17957 25143 18015 25149
rect 17957 25109 17969 25143
rect 18003 25140 18015 25143
rect 18138 25140 18144 25152
rect 18003 25112 18144 25140
rect 18003 25109 18015 25112
rect 17957 25103 18015 25109
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 23017 25143 23075 25149
rect 23017 25109 23029 25143
rect 23063 25140 23075 25143
rect 23566 25140 23572 25152
rect 23063 25112 23572 25140
rect 23063 25109 23075 25112
rect 23017 25103 23075 25109
rect 23566 25100 23572 25112
rect 23624 25100 23630 25152
rect 23845 25143 23903 25149
rect 23845 25109 23857 25143
rect 23891 25140 23903 25143
rect 25498 25140 25504 25152
rect 23891 25112 25504 25140
rect 23891 25109 23903 25112
rect 23845 25103 23903 25109
rect 25498 25100 25504 25112
rect 25556 25100 25562 25152
rect 33505 25143 33563 25149
rect 33505 25109 33517 25143
rect 33551 25140 33563 25143
rect 34698 25140 34704 25152
rect 33551 25112 34704 25140
rect 33551 25109 33563 25112
rect 33505 25103 33563 25109
rect 34698 25100 34704 25112
rect 34756 25100 34762 25152
rect 36832 25149 36860 25180
rect 36817 25143 36875 25149
rect 36817 25109 36829 25143
rect 36863 25109 36875 25143
rect 36817 25103 36875 25109
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 2866 24936 2872 24948
rect 2827 24908 2872 24936
rect 2866 24896 2872 24908
rect 2924 24896 2930 24948
rect 11900 24908 13676 24936
rect 1762 24828 1768 24880
rect 1820 24868 1826 24880
rect 2501 24871 2559 24877
rect 2501 24868 2513 24871
rect 1820 24840 2513 24868
rect 1820 24828 1826 24840
rect 2501 24837 2513 24840
rect 2547 24837 2559 24871
rect 2501 24831 2559 24837
rect 2685 24803 2743 24809
rect 2685 24769 2697 24803
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 4157 24803 4215 24809
rect 4157 24769 4169 24803
rect 4203 24800 4215 24803
rect 4706 24800 4712 24812
rect 4203 24772 4712 24800
rect 4203 24769 4215 24772
rect 4157 24763 4215 24769
rect 2700 24732 2728 24763
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 5718 24732 5724 24744
rect 2700 24704 5724 24732
rect 5718 24692 5724 24704
rect 5776 24692 5782 24744
rect 6564 24732 6592 24763
rect 6730 24760 6736 24812
rect 6788 24800 6794 24812
rect 11900 24809 11928 24908
rect 13446 24828 13452 24880
rect 13504 24868 13510 24880
rect 13648 24868 13676 24908
rect 13906 24896 13912 24948
rect 13964 24896 13970 24948
rect 22189 24939 22247 24945
rect 22189 24905 22201 24939
rect 22235 24936 22247 24939
rect 22554 24936 22560 24948
rect 22235 24908 22560 24936
rect 22235 24905 22247 24908
rect 22189 24899 22247 24905
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 24762 24936 24768 24948
rect 24723 24908 24768 24936
rect 24762 24896 24768 24908
rect 24820 24936 24826 24948
rect 25130 24936 25136 24948
rect 24820 24908 25136 24936
rect 24820 24896 24826 24908
rect 25130 24896 25136 24908
rect 25188 24936 25194 24948
rect 25774 24936 25780 24948
rect 25188 24908 25780 24936
rect 25188 24896 25194 24908
rect 25774 24896 25780 24908
rect 25832 24936 25838 24948
rect 25832 24908 28994 24936
rect 25832 24896 25838 24908
rect 13924 24868 13952 24896
rect 13504 24840 13584 24868
rect 13504 24828 13510 24840
rect 8389 24803 8447 24809
rect 8389 24800 8401 24803
rect 6788 24772 8401 24800
rect 6788 24760 6794 24772
rect 8389 24769 8401 24772
rect 8435 24769 8447 24803
rect 8389 24763 8447 24769
rect 8656 24803 8714 24809
rect 8656 24769 8668 24803
rect 8702 24800 8714 24803
rect 11793 24803 11851 24809
rect 8702 24772 11560 24800
rect 8702 24769 8714 24772
rect 8656 24763 8714 24769
rect 7558 24732 7564 24744
rect 6564 24704 7564 24732
rect 7558 24692 7564 24704
rect 7616 24692 7622 24744
rect 7653 24735 7711 24741
rect 7653 24701 7665 24735
rect 7699 24701 7711 24735
rect 7653 24695 7711 24701
rect 4341 24667 4399 24673
rect 4341 24633 4353 24667
rect 4387 24664 4399 24667
rect 4798 24664 4804 24676
rect 4387 24636 4804 24664
rect 4387 24633 4399 24636
rect 4341 24627 4399 24633
rect 4798 24624 4804 24636
rect 4856 24664 4862 24676
rect 6365 24667 6423 24673
rect 4856 24636 5856 24664
rect 4856 24624 4862 24636
rect 4706 24556 4712 24608
rect 4764 24596 4770 24608
rect 4893 24599 4951 24605
rect 4893 24596 4905 24599
rect 4764 24568 4905 24596
rect 4764 24556 4770 24568
rect 4893 24565 4905 24568
rect 4939 24565 4951 24599
rect 5828 24596 5856 24636
rect 6365 24633 6377 24667
rect 6411 24664 6423 24667
rect 7098 24664 7104 24676
rect 6411 24636 7104 24664
rect 6411 24633 6423 24636
rect 6365 24627 6423 24633
rect 7098 24624 7104 24636
rect 7156 24624 7162 24676
rect 7374 24624 7380 24676
rect 7432 24664 7438 24676
rect 7668 24664 7696 24695
rect 7742 24692 7748 24744
rect 7800 24732 7806 24744
rect 11532 24741 11560 24772
rect 11793 24769 11805 24803
rect 11839 24769 11851 24803
rect 11793 24763 11851 24769
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24769 11943 24803
rect 11885 24763 11943 24769
rect 7929 24735 7987 24741
rect 7929 24732 7941 24735
rect 7800 24704 7941 24732
rect 7800 24692 7806 24704
rect 7929 24701 7941 24704
rect 7975 24701 7987 24735
rect 7929 24695 7987 24701
rect 11517 24735 11575 24741
rect 11517 24701 11529 24735
rect 11563 24701 11575 24735
rect 11517 24695 11575 24701
rect 7432 24636 7696 24664
rect 11808 24664 11836 24763
rect 11974 24760 11980 24812
rect 12032 24800 12038 24812
rect 12158 24800 12164 24812
rect 12032 24772 12077 24800
rect 12119 24772 12164 24800
rect 12032 24760 12038 24772
rect 12158 24760 12164 24772
rect 12216 24760 12222 24812
rect 13556 24809 13584 24840
rect 13648 24840 13952 24868
rect 13648 24809 13676 24840
rect 16942 24828 16948 24880
rect 17000 24868 17006 24880
rect 19245 24871 19303 24877
rect 19245 24868 19257 24871
rect 17000 24840 19257 24868
rect 17000 24828 17006 24840
rect 19245 24837 19257 24840
rect 19291 24837 19303 24871
rect 19245 24831 19303 24837
rect 25332 24840 25820 24868
rect 13541 24803 13599 24809
rect 13541 24769 13553 24803
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 13722 24760 13728 24812
rect 13780 24800 13786 24812
rect 13909 24803 13967 24809
rect 13780 24772 13825 24800
rect 13780 24760 13786 24772
rect 13909 24769 13921 24803
rect 13955 24769 13967 24803
rect 13909 24763 13967 24769
rect 12342 24692 12348 24744
rect 12400 24732 12406 24744
rect 13265 24735 13323 24741
rect 13265 24732 13277 24735
rect 12400 24704 13277 24732
rect 12400 24692 12406 24704
rect 13265 24701 13277 24704
rect 13311 24701 13323 24735
rect 13265 24695 13323 24701
rect 13354 24692 13360 24744
rect 13412 24732 13418 24744
rect 13924 24732 13952 24763
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 15850 24803 15908 24809
rect 15850 24800 15862 24803
rect 14884 24772 15862 24800
rect 14884 24760 14890 24772
rect 15850 24769 15862 24772
rect 15896 24769 15908 24803
rect 16850 24800 16856 24812
rect 16811 24772 16856 24800
rect 15850 24763 15908 24769
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17954 24800 17960 24812
rect 17915 24772 17960 24800
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 18138 24800 18144 24812
rect 18099 24772 18144 24800
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 18233 24803 18291 24809
rect 18233 24769 18245 24803
rect 18279 24769 18291 24803
rect 18233 24763 18291 24769
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24769 18383 24803
rect 19426 24800 19432 24812
rect 19387 24772 19432 24800
rect 18325 24763 18383 24769
rect 14182 24732 14188 24744
rect 13412 24704 14188 24732
rect 13412 24692 13418 24704
rect 14182 24692 14188 24704
rect 14240 24732 14246 24744
rect 14918 24732 14924 24744
rect 14240 24704 14924 24732
rect 14240 24692 14246 24704
rect 14918 24692 14924 24704
rect 14976 24692 14982 24744
rect 16114 24732 16120 24744
rect 16075 24704 16120 24732
rect 16114 24692 16120 24704
rect 16172 24692 16178 24744
rect 17494 24692 17500 24744
rect 17552 24732 17558 24744
rect 17862 24732 17868 24744
rect 17552 24704 17868 24732
rect 17552 24692 17558 24704
rect 17862 24692 17868 24704
rect 17920 24732 17926 24744
rect 18248 24732 18276 24763
rect 17920 24704 18276 24732
rect 17920 24692 17926 24704
rect 12713 24667 12771 24673
rect 12713 24664 12725 24667
rect 11808 24636 12725 24664
rect 7432 24624 7438 24636
rect 12713 24633 12725 24636
rect 12759 24664 12771 24667
rect 12759 24636 15240 24664
rect 12759 24633 12771 24636
rect 12713 24627 12771 24633
rect 6638 24596 6644 24608
rect 5828 24568 6644 24596
rect 4893 24559 4951 24565
rect 6638 24556 6644 24568
rect 6696 24556 6702 24608
rect 9582 24556 9588 24608
rect 9640 24596 9646 24608
rect 9769 24599 9827 24605
rect 9769 24596 9781 24599
rect 9640 24568 9781 24596
rect 9640 24556 9646 24568
rect 9769 24565 9781 24568
rect 9815 24565 9827 24599
rect 9769 24559 9827 24565
rect 14458 24556 14464 24608
rect 14516 24596 14522 24608
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14516 24568 14749 24596
rect 14516 24556 14522 24568
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 15212 24596 15240 24636
rect 18138 24624 18144 24676
rect 18196 24664 18202 24676
rect 18340 24664 18368 24763
rect 19426 24760 19432 24772
rect 19484 24760 19490 24812
rect 19978 24800 19984 24812
rect 19939 24772 19984 24800
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20165 24803 20223 24809
rect 20165 24769 20177 24803
rect 20211 24800 20223 24803
rect 20346 24800 20352 24812
rect 20211 24772 20352 24800
rect 20211 24769 20223 24772
rect 20165 24763 20223 24769
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 21082 24800 21088 24812
rect 21043 24772 21088 24800
rect 21082 24760 21088 24772
rect 21140 24760 21146 24812
rect 21821 24803 21879 24809
rect 21821 24769 21833 24803
rect 21867 24769 21879 24803
rect 22002 24800 22008 24812
rect 21963 24772 22008 24800
rect 21821 24763 21879 24769
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24732 18659 24735
rect 19334 24732 19340 24744
rect 18647 24704 19340 24732
rect 18647 24701 18659 24704
rect 18601 24695 18659 24701
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 21836 24732 21864 24763
rect 22002 24760 22008 24772
rect 22060 24760 22066 24812
rect 23474 24800 23480 24812
rect 22112 24772 23480 24800
rect 21836 24704 21956 24732
rect 19518 24664 19524 24676
rect 18196 24636 19524 24664
rect 18196 24624 18202 24636
rect 19518 24624 19524 24636
rect 19576 24664 19582 24676
rect 20898 24664 20904 24676
rect 19576 24636 20904 24664
rect 19576 24624 19582 24636
rect 20898 24624 20904 24636
rect 20956 24624 20962 24676
rect 21269 24667 21327 24673
rect 21269 24633 21281 24667
rect 21315 24664 21327 24667
rect 21928 24664 21956 24704
rect 22112 24664 22140 24772
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 23566 24760 23572 24812
rect 23624 24800 23630 24812
rect 23946 24803 24004 24809
rect 23946 24800 23958 24803
rect 23624 24772 23958 24800
rect 23624 24760 23630 24772
rect 23946 24769 23958 24772
rect 23992 24769 24004 24803
rect 24210 24800 24216 24812
rect 24171 24772 24216 24800
rect 23946 24763 24004 24769
rect 24210 24760 24216 24772
rect 24268 24760 24274 24812
rect 25222 24760 25228 24812
rect 25280 24800 25286 24812
rect 25332 24809 25360 24840
rect 25317 24803 25375 24809
rect 25317 24800 25329 24803
rect 25280 24772 25329 24800
rect 25280 24760 25286 24772
rect 25317 24769 25329 24772
rect 25363 24769 25375 24803
rect 25498 24800 25504 24812
rect 25459 24772 25504 24800
rect 25317 24763 25375 24769
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 25593 24803 25651 24809
rect 25593 24769 25605 24803
rect 25639 24769 25651 24803
rect 25593 24763 25651 24769
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25792 24800 25820 24840
rect 26234 24828 26240 24880
rect 26292 24868 26298 24880
rect 26292 24840 27384 24868
rect 26292 24828 26298 24840
rect 27356 24812 27384 24840
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 25792 24772 26985 24800
rect 25685 24763 25743 24769
rect 26973 24769 26985 24772
rect 27019 24769 27031 24803
rect 27154 24800 27160 24812
rect 27115 24772 27160 24800
rect 26973 24763 27031 24769
rect 21315 24636 22140 24664
rect 21315 24633 21327 24636
rect 21269 24627 21327 24633
rect 24210 24624 24216 24676
rect 24268 24664 24274 24676
rect 25498 24664 25504 24676
rect 24268 24636 25504 24664
rect 24268 24624 24274 24636
rect 25498 24624 25504 24636
rect 25556 24664 25562 24676
rect 25608 24664 25636 24763
rect 25700 24732 25728 24763
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 27249 24803 27307 24809
rect 27249 24769 27261 24803
rect 27295 24769 27307 24803
rect 27249 24763 27307 24769
rect 25774 24732 25780 24744
rect 25700 24704 25780 24732
rect 25774 24692 25780 24704
rect 25832 24692 25838 24744
rect 25961 24735 26019 24741
rect 25961 24701 25973 24735
rect 26007 24732 26019 24735
rect 26326 24732 26332 24744
rect 26007 24704 26332 24732
rect 26007 24701 26019 24704
rect 25961 24695 26019 24701
rect 26326 24692 26332 24704
rect 26384 24692 26390 24744
rect 27264 24664 27292 24763
rect 27338 24760 27344 24812
rect 27396 24800 27402 24812
rect 27396 24772 27489 24800
rect 27396 24760 27402 24772
rect 27706 24760 27712 24812
rect 27764 24800 27770 24812
rect 28077 24803 28135 24809
rect 28077 24800 28089 24803
rect 27764 24772 28089 24800
rect 27764 24760 27770 24772
rect 28077 24769 28089 24772
rect 28123 24800 28135 24803
rect 28350 24800 28356 24812
rect 28123 24772 28356 24800
rect 28123 24769 28135 24772
rect 28077 24763 28135 24769
rect 28350 24760 28356 24772
rect 28408 24760 28414 24812
rect 28966 24732 28994 24908
rect 30926 24896 30932 24948
rect 30984 24936 30990 24948
rect 31113 24939 31171 24945
rect 31113 24936 31125 24939
rect 30984 24908 31125 24936
rect 30984 24896 30990 24908
rect 31113 24905 31125 24908
rect 31159 24905 31171 24939
rect 32401 24939 32459 24945
rect 32401 24936 32413 24939
rect 31113 24899 31171 24905
rect 31726 24908 32413 24936
rect 30282 24800 30288 24812
rect 30243 24772 30288 24800
rect 30282 24760 30288 24772
rect 30340 24800 30346 24812
rect 30929 24803 30987 24809
rect 30929 24800 30941 24803
rect 30340 24772 30941 24800
rect 30340 24760 30346 24772
rect 30929 24769 30941 24772
rect 30975 24769 30987 24803
rect 30929 24763 30987 24769
rect 31726 24732 31754 24908
rect 32401 24905 32413 24908
rect 32447 24936 32459 24939
rect 32858 24936 32864 24948
rect 32447 24908 32864 24936
rect 32447 24905 32459 24908
rect 32401 24899 32459 24905
rect 32858 24896 32864 24908
rect 32916 24896 32922 24948
rect 32490 24760 32496 24812
rect 32548 24800 32554 24812
rect 33045 24803 33103 24809
rect 33045 24800 33057 24803
rect 32548 24772 33057 24800
rect 32548 24760 32554 24772
rect 33045 24769 33057 24772
rect 33091 24769 33103 24803
rect 33045 24763 33103 24769
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 33229 24803 33287 24809
rect 33229 24800 33241 24803
rect 33192 24772 33241 24800
rect 33192 24760 33198 24772
rect 33229 24769 33241 24772
rect 33275 24769 33287 24803
rect 33229 24763 33287 24769
rect 33321 24803 33379 24809
rect 33321 24769 33333 24803
rect 33367 24769 33379 24803
rect 33321 24763 33379 24769
rect 28966 24704 31754 24732
rect 32858 24692 32864 24744
rect 32916 24732 32922 24744
rect 33336 24732 33364 24763
rect 33410 24760 33416 24812
rect 33468 24800 33474 24812
rect 33468 24772 33513 24800
rect 33468 24760 33474 24772
rect 34422 24760 34428 24812
rect 34480 24800 34486 24812
rect 34701 24803 34759 24809
rect 34701 24800 34713 24803
rect 34480 24772 34713 24800
rect 34480 24760 34486 24772
rect 34701 24769 34713 24772
rect 34747 24769 34759 24803
rect 34957 24803 35015 24809
rect 34957 24800 34969 24803
rect 34701 24763 34759 24769
rect 34808 24772 34969 24800
rect 32916 24704 33364 24732
rect 33689 24735 33747 24741
rect 32916 24692 32922 24704
rect 33689 24701 33701 24735
rect 33735 24732 33747 24735
rect 34808 24732 34836 24772
rect 34957 24769 34969 24772
rect 35003 24769 35015 24803
rect 34957 24763 35015 24769
rect 33735 24704 34836 24732
rect 33735 24701 33747 24704
rect 33689 24695 33747 24701
rect 25556 24636 27292 24664
rect 30469 24667 30527 24673
rect 25556 24624 25562 24636
rect 30469 24633 30481 24667
rect 30515 24664 30527 24667
rect 31754 24664 31760 24676
rect 30515 24636 31760 24664
rect 30515 24633 30527 24636
rect 30469 24627 30527 24633
rect 31754 24624 31760 24636
rect 31812 24624 31818 24676
rect 18156 24596 18184 24624
rect 15212 24568 18184 24596
rect 14737 24559 14795 24565
rect 22002 24556 22008 24608
rect 22060 24596 22066 24608
rect 22833 24599 22891 24605
rect 22833 24596 22845 24599
rect 22060 24568 22845 24596
rect 22060 24556 22066 24568
rect 22833 24565 22845 24568
rect 22879 24565 22891 24599
rect 22833 24559 22891 24565
rect 27522 24556 27528 24608
rect 27580 24596 27586 24608
rect 27617 24599 27675 24605
rect 27617 24596 27629 24599
rect 27580 24568 27629 24596
rect 27580 24556 27586 24568
rect 27617 24565 27629 24568
rect 27663 24565 27675 24599
rect 27617 24559 27675 24565
rect 32950 24556 32956 24608
rect 33008 24596 33014 24608
rect 36081 24599 36139 24605
rect 36081 24596 36093 24599
rect 33008 24568 36093 24596
rect 33008 24556 33014 24568
rect 36081 24565 36093 24568
rect 36127 24565 36139 24599
rect 36081 24559 36139 24565
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 1762 24392 1768 24404
rect 1723 24364 1768 24392
rect 1762 24352 1768 24364
rect 1820 24352 1826 24404
rect 2958 24352 2964 24404
rect 3016 24401 3022 24404
rect 3016 24395 3065 24401
rect 3016 24361 3019 24395
rect 3053 24361 3065 24395
rect 3016 24355 3065 24361
rect 9401 24395 9459 24401
rect 9401 24361 9413 24395
rect 9447 24392 9459 24395
rect 11974 24392 11980 24404
rect 9447 24364 11980 24392
rect 9447 24361 9459 24364
rect 9401 24355 9459 24361
rect 3016 24352 3022 24355
rect 11974 24352 11980 24364
rect 12032 24352 12038 24404
rect 13173 24395 13231 24401
rect 13173 24361 13185 24395
rect 13219 24392 13231 24395
rect 13722 24392 13728 24404
rect 13219 24364 13728 24392
rect 13219 24361 13231 24364
rect 13173 24355 13231 24361
rect 13722 24352 13728 24364
rect 13780 24352 13786 24404
rect 14826 24392 14832 24404
rect 14787 24364 14832 24392
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 14918 24352 14924 24404
rect 14976 24392 14982 24404
rect 14976 24364 22094 24392
rect 14976 24352 14982 24364
rect 6638 24284 6644 24336
rect 6696 24324 6702 24336
rect 14550 24324 14556 24336
rect 6696 24296 14556 24324
rect 6696 24284 6702 24296
rect 14550 24284 14556 24296
rect 14608 24284 14614 24336
rect 16482 24284 16488 24336
rect 16540 24324 16546 24336
rect 22066 24324 22094 24364
rect 23290 24352 23296 24404
rect 23348 24392 23354 24404
rect 23385 24395 23443 24401
rect 23385 24392 23397 24395
rect 23348 24364 23397 24392
rect 23348 24352 23354 24364
rect 23385 24361 23397 24364
rect 23431 24361 23443 24395
rect 23385 24355 23443 24361
rect 25409 24395 25467 24401
rect 25409 24361 25421 24395
rect 25455 24392 25467 24395
rect 27154 24392 27160 24404
rect 25455 24364 27160 24392
rect 25455 24361 25467 24364
rect 25409 24355 25467 24361
rect 27154 24352 27160 24364
rect 27212 24352 27218 24404
rect 31757 24395 31815 24401
rect 31757 24392 31769 24395
rect 28552 24364 31769 24392
rect 22278 24324 22284 24336
rect 16540 24296 19840 24324
rect 22066 24296 22284 24324
rect 16540 24284 16546 24296
rect 5166 24216 5172 24268
rect 5224 24256 5230 24268
rect 5224 24228 10548 24256
rect 5224 24216 5230 24228
rect 1949 24191 2007 24197
rect 1949 24157 1961 24191
rect 1995 24157 2007 24191
rect 1949 24151 2007 24157
rect 3237 24191 3295 24197
rect 3237 24157 3249 24191
rect 3283 24157 3295 24191
rect 3237 24151 3295 24157
rect 1964 24120 1992 24151
rect 2498 24120 2504 24132
rect 1964 24092 2504 24120
rect 2498 24080 2504 24092
rect 2556 24080 2562 24132
rect 2866 24080 2872 24132
rect 2924 24120 2930 24132
rect 3252 24120 3280 24151
rect 3326 24148 3332 24200
rect 3384 24188 3390 24200
rect 3789 24191 3847 24197
rect 3789 24188 3801 24191
rect 3384 24160 3801 24188
rect 3384 24148 3390 24160
rect 3789 24157 3801 24160
rect 3835 24157 3847 24191
rect 3970 24188 3976 24200
rect 3931 24160 3976 24188
rect 3789 24151 3847 24157
rect 3970 24148 3976 24160
rect 4028 24148 4034 24200
rect 4065 24191 4123 24197
rect 4065 24157 4077 24191
rect 4111 24157 4123 24191
rect 4065 24151 4123 24157
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4893 24191 4951 24197
rect 4893 24188 4905 24191
rect 4203 24160 4905 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4893 24157 4905 24160
rect 4939 24188 4951 24191
rect 7834 24188 7840 24200
rect 4939 24160 7840 24188
rect 4939 24157 4951 24160
rect 4893 24151 4951 24157
rect 2924 24092 3280 24120
rect 2924 24080 2930 24092
rect 2682 24012 2688 24064
rect 2740 24052 2746 24064
rect 4080 24052 4108 24151
rect 7834 24148 7840 24160
rect 7892 24148 7898 24200
rect 9582 24188 9588 24200
rect 9543 24160 9588 24188
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 10226 24188 10232 24200
rect 10187 24160 10232 24188
rect 10226 24148 10232 24160
rect 10284 24148 10290 24200
rect 5537 24123 5595 24129
rect 5537 24089 5549 24123
rect 5583 24120 5595 24123
rect 6638 24120 6644 24132
rect 5583 24092 6644 24120
rect 5583 24089 5595 24092
rect 5537 24083 5595 24089
rect 6638 24080 6644 24092
rect 6696 24120 6702 24132
rect 7745 24123 7803 24129
rect 7745 24120 7757 24123
rect 6696 24092 7757 24120
rect 6696 24080 6702 24092
rect 7745 24089 7757 24092
rect 7791 24089 7803 24123
rect 7745 24083 7803 24089
rect 9769 24123 9827 24129
rect 9769 24089 9781 24123
rect 9815 24089 9827 24123
rect 9769 24083 9827 24089
rect 4430 24052 4436 24064
rect 2740 24024 4108 24052
rect 4391 24024 4436 24052
rect 2740 24012 2746 24024
rect 4430 24012 4436 24024
rect 4488 24012 4494 24064
rect 6730 24012 6736 24064
rect 6788 24052 6794 24064
rect 6825 24055 6883 24061
rect 6825 24052 6837 24055
rect 6788 24024 6837 24052
rect 6788 24012 6794 24024
rect 6825 24021 6837 24024
rect 6871 24021 6883 24055
rect 9784 24052 9812 24083
rect 10134 24080 10140 24132
rect 10192 24120 10198 24132
rect 10520 24129 10548 24228
rect 17494 24216 17500 24268
rect 17552 24256 17558 24268
rect 17552 24228 19564 24256
rect 17552 24216 17558 24228
rect 10594 24148 10600 24200
rect 10652 24188 10658 24200
rect 10652 24160 10697 24188
rect 10652 24148 10658 24160
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 12989 24191 13047 24197
rect 12989 24188 13001 24191
rect 12492 24160 13001 24188
rect 12492 24148 12498 24160
rect 12989 24157 13001 24160
rect 13035 24157 13047 24191
rect 12989 24151 13047 24157
rect 13354 24148 13360 24200
rect 13412 24188 13418 24200
rect 14173 24191 14231 24197
rect 14173 24188 14185 24191
rect 13412 24160 14185 24188
rect 13412 24148 13418 24160
rect 14173 24157 14185 24160
rect 14219 24157 14231 24191
rect 14366 24188 14372 24200
rect 14327 24160 14372 24188
rect 14173 24151 14231 24157
rect 14366 24148 14372 24160
rect 14424 24148 14430 24200
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24157 14611 24191
rect 14553 24151 14611 24157
rect 10413 24123 10471 24129
rect 10413 24120 10425 24123
rect 10192 24092 10425 24120
rect 10192 24080 10198 24092
rect 10413 24089 10425 24092
rect 10459 24089 10471 24123
rect 10413 24083 10471 24089
rect 10505 24123 10563 24129
rect 10505 24089 10517 24123
rect 10551 24089 10563 24123
rect 12618 24120 12624 24132
rect 10505 24083 10563 24089
rect 10704 24092 12624 24120
rect 10704 24052 10732 24092
rect 12618 24080 12624 24092
rect 12676 24120 12682 24132
rect 12805 24123 12863 24129
rect 12805 24120 12817 24123
rect 12676 24092 12817 24120
rect 12676 24080 12682 24092
rect 12805 24089 12817 24092
rect 12851 24120 12863 24123
rect 13170 24120 13176 24132
rect 12851 24092 13176 24120
rect 12851 24089 12863 24092
rect 12805 24083 12863 24089
rect 13170 24080 13176 24092
rect 13228 24080 13234 24132
rect 13906 24080 13912 24132
rect 13964 24120 13970 24132
rect 14476 24120 14504 24151
rect 13964 24092 14504 24120
rect 14568 24120 14596 24151
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 17129 24191 17187 24197
rect 17129 24188 17141 24191
rect 15252 24160 17141 24188
rect 15252 24148 15258 24160
rect 17129 24157 17141 24160
rect 17175 24157 17187 24191
rect 17129 24151 17187 24157
rect 17586 24148 17592 24200
rect 17644 24148 17650 24200
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 18012 24160 19257 24188
rect 18012 24148 18018 24160
rect 19245 24157 19257 24160
rect 19291 24157 19303 24191
rect 19426 24188 19432 24200
rect 19387 24160 19432 24188
rect 19245 24151 19303 24157
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 19536 24197 19564 24228
rect 19521 24191 19579 24197
rect 19521 24157 19533 24191
rect 19567 24157 19579 24191
rect 19521 24151 19579 24157
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 15289 24123 15347 24129
rect 15289 24120 15301 24123
rect 14568 24092 15301 24120
rect 13964 24080 13970 24092
rect 15289 24089 15301 24092
rect 15335 24120 15347 24123
rect 16850 24120 16856 24132
rect 15335 24092 16856 24120
rect 15335 24089 15347 24092
rect 15289 24083 15347 24089
rect 16850 24080 16856 24092
rect 16908 24080 16914 24132
rect 16945 24123 17003 24129
rect 16945 24089 16957 24123
rect 16991 24120 17003 24123
rect 17604 24120 17632 24148
rect 18230 24120 18236 24132
rect 16991 24092 18236 24120
rect 16991 24089 17003 24092
rect 16945 24083 17003 24089
rect 18230 24080 18236 24092
rect 18288 24080 18294 24132
rect 19150 24080 19156 24132
rect 19208 24120 19214 24132
rect 19628 24120 19656 24151
rect 19208 24092 19656 24120
rect 19812 24120 19840 24296
rect 22278 24284 22284 24296
rect 22336 24324 22342 24336
rect 23842 24324 23848 24336
rect 22336 24296 23848 24324
rect 22336 24284 22342 24296
rect 23842 24284 23848 24296
rect 23900 24284 23906 24336
rect 25682 24284 25688 24336
rect 25740 24324 25746 24336
rect 25869 24327 25927 24333
rect 25869 24324 25881 24327
rect 25740 24296 25881 24324
rect 25740 24284 25746 24296
rect 25869 24293 25881 24296
rect 25915 24293 25927 24327
rect 25869 24287 25927 24293
rect 21361 24259 21419 24265
rect 21361 24225 21373 24259
rect 21407 24256 21419 24259
rect 21818 24256 21824 24268
rect 21407 24228 21824 24256
rect 21407 24225 21419 24228
rect 21361 24219 21419 24225
rect 21818 24216 21824 24228
rect 21876 24256 21882 24268
rect 22833 24259 22891 24265
rect 22833 24256 22845 24259
rect 21876 24228 22845 24256
rect 21876 24216 21882 24228
rect 22833 24225 22845 24228
rect 22879 24225 22891 24259
rect 24210 24256 24216 24268
rect 22833 24219 22891 24225
rect 23124 24228 24216 24256
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 21269 24191 21327 24197
rect 21269 24188 21281 24191
rect 20956 24160 21281 24188
rect 20956 24148 20962 24160
rect 21269 24157 21281 24160
rect 21315 24157 21327 24191
rect 21269 24151 21327 24157
rect 21453 24191 21511 24197
rect 21453 24157 21465 24191
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24188 22615 24191
rect 22646 24188 22652 24200
rect 22603 24160 22652 24188
rect 22603 24157 22615 24160
rect 22557 24151 22615 24157
rect 21468 24120 21496 24151
rect 22646 24148 22652 24160
rect 22704 24188 22710 24200
rect 23124 24188 23152 24228
rect 24210 24216 24216 24228
rect 24268 24216 24274 24268
rect 27798 24256 27804 24268
rect 27759 24228 27804 24256
rect 27798 24216 27804 24228
rect 27856 24216 27862 24268
rect 22704 24160 23152 24188
rect 22704 24148 22710 24160
rect 23198 24148 23204 24200
rect 23256 24188 23262 24200
rect 23293 24191 23351 24197
rect 23293 24188 23305 24191
rect 23256 24160 23305 24188
rect 23256 24148 23262 24160
rect 23293 24157 23305 24160
rect 23339 24157 23351 24191
rect 23293 24151 23351 24157
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 23566 24188 23572 24200
rect 23523 24160 23572 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 24854 24148 24860 24200
rect 24912 24188 24918 24200
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 24912 24160 25053 24188
rect 24912 24148 24918 24160
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 27522 24148 27528 24200
rect 27580 24197 27586 24200
rect 27580 24188 27592 24197
rect 28350 24188 28356 24200
rect 27580 24160 27625 24188
rect 28311 24160 28356 24188
rect 27580 24151 27592 24160
rect 27580 24148 27586 24151
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 28552 24197 28580 24364
rect 31757 24361 31769 24364
rect 31803 24361 31815 24395
rect 33134 24392 33140 24404
rect 33095 24364 33140 24392
rect 31757 24355 31815 24361
rect 33134 24352 33140 24364
rect 33192 24352 33198 24404
rect 30558 24284 30564 24336
rect 30616 24324 30622 24336
rect 33410 24324 33416 24336
rect 30616 24296 33416 24324
rect 30616 24284 30622 24296
rect 33410 24284 33416 24296
rect 33468 24324 33474 24336
rect 33597 24327 33655 24333
rect 33597 24324 33609 24327
rect 33468 24296 33609 24324
rect 33468 24284 33474 24296
rect 33597 24293 33609 24296
rect 33643 24293 33655 24327
rect 33597 24287 33655 24293
rect 28902 24256 28908 24268
rect 28644 24228 28908 24256
rect 28644 24197 28672 24228
rect 28902 24216 28908 24228
rect 28960 24256 28966 24268
rect 29454 24256 29460 24268
rect 28960 24228 29460 24256
rect 28960 24216 28966 24228
rect 29454 24216 29460 24228
rect 29512 24216 29518 24268
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 28629 24191 28687 24197
rect 28629 24157 28641 24191
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 28721 24191 28779 24197
rect 28721 24157 28733 24191
rect 28767 24157 28779 24191
rect 28721 24151 28779 24157
rect 29549 24191 29607 24197
rect 29549 24157 29561 24191
rect 29595 24188 29607 24191
rect 31938 24188 31944 24200
rect 29595 24160 31944 24188
rect 29595 24157 29607 24160
rect 29549 24151 29607 24157
rect 23216 24120 23244 24148
rect 19812 24092 23244 24120
rect 19208 24080 19214 24092
rect 23750 24080 23756 24132
rect 23808 24120 23814 24132
rect 25225 24123 25283 24129
rect 23808 24092 24992 24120
rect 23808 24080 23814 24092
rect 9784 24024 10732 24052
rect 10781 24055 10839 24061
rect 6825 24015 6883 24021
rect 10781 24021 10793 24055
rect 10827 24052 10839 24055
rect 11146 24052 11152 24064
rect 10827 24024 11152 24052
rect 10827 24021 10839 24024
rect 10781 24015 10839 24021
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 11333 24055 11391 24061
rect 11333 24021 11345 24055
rect 11379 24052 11391 24055
rect 11514 24052 11520 24064
rect 11379 24024 11520 24052
rect 11379 24021 11391 24024
rect 11333 24015 11391 24021
rect 11514 24012 11520 24024
rect 11572 24012 11578 24064
rect 17313 24055 17371 24061
rect 17313 24021 17325 24055
rect 17359 24052 17371 24055
rect 17586 24052 17592 24064
rect 17359 24024 17592 24052
rect 17359 24021 17371 24024
rect 17313 24015 17371 24021
rect 17586 24012 17592 24024
rect 17644 24012 17650 24064
rect 18138 24052 18144 24064
rect 18099 24024 18144 24052
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 18693 24055 18751 24061
rect 18693 24021 18705 24055
rect 18739 24052 18751 24055
rect 19334 24052 19340 24064
rect 18739 24024 19340 24052
rect 18739 24021 18751 24024
rect 18693 24015 18751 24021
rect 19334 24012 19340 24024
rect 19392 24012 19398 24064
rect 19889 24055 19947 24061
rect 19889 24021 19901 24055
rect 19935 24052 19947 24055
rect 19978 24052 19984 24064
rect 19935 24024 19984 24052
rect 19935 24021 19947 24024
rect 19889 24015 19947 24021
rect 19978 24012 19984 24024
rect 20036 24012 20042 24064
rect 20346 24052 20352 24064
rect 20307 24024 20352 24052
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 24302 24012 24308 24064
rect 24360 24052 24366 24064
rect 24397 24055 24455 24061
rect 24397 24052 24409 24055
rect 24360 24024 24409 24052
rect 24360 24012 24366 24024
rect 24397 24021 24409 24024
rect 24443 24021 24455 24055
rect 24964 24052 24992 24092
rect 25225 24089 25237 24123
rect 25271 24120 25283 24123
rect 25271 24092 26464 24120
rect 25271 24089 25283 24092
rect 25225 24083 25283 24089
rect 25240 24052 25268 24083
rect 26436 24061 26464 24092
rect 28166 24080 28172 24132
rect 28224 24120 28230 24132
rect 28736 24120 28764 24151
rect 31938 24148 31944 24160
rect 31996 24188 32002 24200
rect 34422 24188 34428 24200
rect 31996 24160 34428 24188
rect 31996 24148 32002 24160
rect 34422 24148 34428 24160
rect 34480 24148 34486 24200
rect 68094 24188 68100 24200
rect 68055 24160 68100 24188
rect 68094 24148 68100 24160
rect 68152 24148 68158 24200
rect 28224 24092 28764 24120
rect 28997 24123 29055 24129
rect 28224 24080 28230 24092
rect 28997 24089 29009 24123
rect 29043 24120 29055 24123
rect 29794 24123 29852 24129
rect 29794 24120 29806 24123
rect 29043 24092 29806 24120
rect 29043 24089 29055 24092
rect 28997 24083 29055 24089
rect 29794 24089 29806 24092
rect 29840 24089 29852 24123
rect 29794 24083 29852 24089
rect 30282 24080 30288 24132
rect 30340 24120 30346 24132
rect 31389 24123 31447 24129
rect 31389 24120 31401 24123
rect 30340 24092 31401 24120
rect 30340 24080 30346 24092
rect 31389 24089 31401 24092
rect 31435 24089 31447 24123
rect 31389 24083 31447 24089
rect 31573 24123 31631 24129
rect 31573 24089 31585 24123
rect 31619 24089 31631 24123
rect 31573 24083 31631 24089
rect 24964 24024 25268 24052
rect 26421 24055 26479 24061
rect 24397 24015 24455 24021
rect 26421 24021 26433 24055
rect 26467 24021 26479 24055
rect 26421 24015 26479 24021
rect 27338 24012 27344 24064
rect 27396 24052 27402 24064
rect 30558 24052 30564 24064
rect 27396 24024 30564 24052
rect 27396 24012 27402 24024
rect 30558 24012 30564 24024
rect 30616 24012 30622 24064
rect 30929 24055 30987 24061
rect 30929 24021 30941 24055
rect 30975 24052 30987 24055
rect 31294 24052 31300 24064
rect 30975 24024 31300 24052
rect 30975 24021 30987 24024
rect 30929 24015 30987 24021
rect 31294 24012 31300 24024
rect 31352 24052 31358 24064
rect 31588 24052 31616 24083
rect 31662 24080 31668 24132
rect 31720 24120 31726 24132
rect 31720 24092 32720 24120
rect 31720 24080 31726 24092
rect 32214 24052 32220 24064
rect 31352 24024 31616 24052
rect 32175 24024 32220 24052
rect 31352 24012 31358 24024
rect 32214 24012 32220 24024
rect 32272 24012 32278 24064
rect 32692 24052 32720 24092
rect 32766 24080 32772 24132
rect 32824 24120 32830 24132
rect 32950 24120 32956 24132
rect 32824 24092 32869 24120
rect 32911 24092 32956 24120
rect 32824 24080 32830 24092
rect 32950 24080 32956 24092
rect 33008 24080 33014 24132
rect 36722 24052 36728 24064
rect 32692 24024 36728 24052
rect 36722 24012 36728 24024
rect 36780 24012 36786 24064
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 5626 23808 5632 23860
rect 5684 23848 5690 23860
rect 5721 23851 5779 23857
rect 5721 23848 5733 23851
rect 5684 23820 5733 23848
rect 5684 23808 5690 23820
rect 5721 23817 5733 23820
rect 5767 23817 5779 23851
rect 7098 23848 7104 23860
rect 5721 23811 5779 23817
rect 6564 23820 7104 23848
rect 4056 23783 4114 23789
rect 4056 23749 4068 23783
rect 4102 23780 4114 23783
rect 4430 23780 4436 23792
rect 4102 23752 4436 23780
rect 4102 23749 4114 23752
rect 4056 23743 4114 23749
rect 4430 23740 4436 23752
rect 4488 23740 4494 23792
rect 6564 23789 6592 23820
rect 7098 23808 7104 23820
rect 7156 23808 7162 23860
rect 8757 23851 8815 23857
rect 8757 23817 8769 23851
rect 8803 23848 8815 23851
rect 14642 23848 14648 23860
rect 8803 23820 11744 23848
rect 8803 23817 8815 23820
rect 8757 23811 8815 23817
rect 6549 23783 6607 23789
rect 6549 23749 6561 23783
rect 6595 23749 6607 23783
rect 6549 23743 6607 23749
rect 6733 23783 6791 23789
rect 6733 23749 6745 23783
rect 6779 23780 6791 23783
rect 8772 23780 8800 23811
rect 6779 23752 8800 23780
rect 6779 23749 6791 23752
rect 6733 23743 6791 23749
rect 2314 23712 2320 23724
rect 2275 23684 2320 23712
rect 2314 23672 2320 23684
rect 2372 23672 2378 23724
rect 3786 23712 3792 23724
rect 3747 23684 3792 23712
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 6822 23672 6828 23724
rect 6880 23712 6886 23724
rect 7377 23715 7435 23721
rect 7377 23712 7389 23715
rect 6880 23684 7389 23712
rect 6880 23672 6886 23684
rect 7377 23681 7389 23684
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 7466 23672 7472 23724
rect 7524 23712 7530 23724
rect 7633 23715 7691 23721
rect 7633 23712 7645 23715
rect 7524 23684 7645 23712
rect 7524 23672 7530 23684
rect 7633 23681 7645 23684
rect 7679 23681 7691 23715
rect 7633 23675 7691 23681
rect 9582 23672 9588 23724
rect 9640 23712 9646 23724
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 9640 23684 9965 23712
rect 9640 23672 9646 23684
rect 9953 23681 9965 23684
rect 9999 23681 10011 23715
rect 10134 23712 10140 23724
rect 10095 23684 10140 23712
rect 9953 23675 10011 23681
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23681 10287 23715
rect 10229 23675 10287 23681
rect 10321 23715 10379 23721
rect 10321 23681 10333 23715
rect 10367 23712 10379 23715
rect 10594 23712 10600 23724
rect 10367 23684 10600 23712
rect 10367 23681 10379 23684
rect 10321 23675 10379 23681
rect 2593 23647 2651 23653
rect 2593 23613 2605 23647
rect 2639 23644 2651 23647
rect 2639 23616 2774 23644
rect 2639 23613 2651 23616
rect 2593 23607 2651 23613
rect 2746 23508 2774 23616
rect 5166 23576 5172 23588
rect 5127 23548 5172 23576
rect 5166 23536 5172 23548
rect 5224 23536 5230 23588
rect 5626 23536 5632 23588
rect 5684 23576 5690 23588
rect 5684 23548 7052 23576
rect 5684 23536 5690 23548
rect 3142 23508 3148 23520
rect 2746 23480 3148 23508
rect 3142 23468 3148 23480
rect 3200 23468 3206 23520
rect 6914 23508 6920 23520
rect 6875 23480 6920 23508
rect 6914 23468 6920 23480
rect 6972 23468 6978 23520
rect 7024 23508 7052 23548
rect 10244 23508 10272 23675
rect 10594 23672 10600 23684
rect 10652 23672 10658 23724
rect 7024 23480 10272 23508
rect 10505 23511 10563 23517
rect 10505 23477 10517 23511
rect 10551 23508 10563 23511
rect 11606 23508 11612 23520
rect 10551 23480 11612 23508
rect 10551 23477 10563 23480
rect 10505 23471 10563 23477
rect 11606 23468 11612 23480
rect 11664 23468 11670 23520
rect 11716 23508 11744 23820
rect 12048 23820 14648 23848
rect 11882 23712 11888 23724
rect 11843 23684 11888 23712
rect 11882 23672 11888 23684
rect 11940 23672 11946 23724
rect 12048 23721 12076 23820
rect 14642 23808 14648 23820
rect 14700 23808 14706 23860
rect 14737 23851 14795 23857
rect 14737 23817 14749 23851
rect 14783 23848 14795 23851
rect 15194 23848 15200 23860
rect 14783 23820 15200 23848
rect 14783 23817 14795 23820
rect 14737 23811 14795 23817
rect 15194 23808 15200 23820
rect 15252 23808 15258 23860
rect 16022 23808 16028 23860
rect 16080 23848 16086 23860
rect 18601 23851 18659 23857
rect 16080 23820 18460 23848
rect 16080 23808 16086 23820
rect 13906 23780 13912 23792
rect 13648 23752 13912 23780
rect 12033 23715 12091 23721
rect 12033 23681 12045 23715
rect 12079 23681 12091 23715
rect 12033 23675 12091 23681
rect 12161 23715 12219 23721
rect 12161 23681 12173 23715
rect 12207 23681 12219 23715
rect 12161 23675 12219 23681
rect 12253 23715 12311 23721
rect 12253 23681 12265 23715
rect 12299 23681 12311 23715
rect 12253 23675 12311 23681
rect 12176 23588 12204 23675
rect 12158 23536 12164 23588
rect 12216 23536 12222 23588
rect 12268 23508 12296 23675
rect 12342 23672 12348 23724
rect 12400 23721 12406 23724
rect 12400 23712 12408 23721
rect 13354 23712 13360 23724
rect 12400 23684 12445 23712
rect 13315 23684 13360 23712
rect 12400 23675 12408 23684
rect 12400 23672 12406 23675
rect 13354 23672 13360 23684
rect 13412 23672 13418 23724
rect 13538 23712 13544 23724
rect 13499 23684 13544 23712
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 13648 23721 13676 23752
rect 13906 23740 13912 23752
rect 13964 23740 13970 23792
rect 18432 23789 18460 23820
rect 18601 23817 18613 23851
rect 18647 23848 18659 23851
rect 19426 23848 19432 23860
rect 18647 23820 19432 23848
rect 18647 23817 18659 23820
rect 18601 23811 18659 23817
rect 19426 23808 19432 23820
rect 19484 23808 19490 23860
rect 20717 23851 20775 23857
rect 20717 23848 20729 23851
rect 19536 23820 20729 23848
rect 15872 23783 15930 23789
rect 15872 23749 15884 23783
rect 15918 23780 15930 23783
rect 17129 23783 17187 23789
rect 17129 23780 17141 23783
rect 15918 23752 17141 23780
rect 15918 23749 15930 23752
rect 15872 23743 15930 23749
rect 17129 23749 17141 23752
rect 17175 23749 17187 23783
rect 18417 23783 18475 23789
rect 17129 23743 17187 23749
rect 17236 23752 17816 23780
rect 13633 23715 13691 23721
rect 13633 23681 13645 23715
rect 13679 23681 13691 23715
rect 13633 23675 13691 23681
rect 13725 23715 13783 23721
rect 13725 23681 13737 23715
rect 13771 23712 13783 23715
rect 15470 23712 15476 23724
rect 13771 23684 15476 23712
rect 13771 23681 13783 23684
rect 13725 23675 13783 23681
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 16758 23672 16764 23724
rect 16816 23712 16822 23724
rect 17236 23712 17264 23752
rect 17402 23712 17408 23724
rect 16816 23684 17264 23712
rect 17363 23684 17408 23712
rect 16816 23672 16822 23684
rect 17402 23672 17408 23684
rect 17460 23672 17466 23724
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23681 17555 23715
rect 17497 23675 17555 23681
rect 16114 23644 16120 23656
rect 16075 23616 16120 23644
rect 16114 23604 16120 23616
rect 16172 23604 16178 23656
rect 17512 23588 17540 23675
rect 17586 23672 17592 23724
rect 17644 23712 17650 23724
rect 17788 23721 17816 23752
rect 18417 23749 18429 23783
rect 18463 23780 18475 23783
rect 19536 23780 19564 23820
rect 20717 23817 20729 23820
rect 20763 23817 20775 23851
rect 22278 23848 22284 23860
rect 22239 23820 22284 23848
rect 20717 23811 20775 23817
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 23474 23848 23480 23860
rect 22940 23820 23480 23848
rect 18463 23752 19564 23780
rect 19604 23783 19662 23789
rect 18463 23749 18475 23752
rect 18417 23743 18475 23749
rect 19604 23749 19616 23783
rect 19650 23780 19662 23783
rect 19978 23780 19984 23792
rect 19650 23752 19984 23780
rect 19650 23749 19662 23752
rect 19604 23743 19662 23749
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 20346 23740 20352 23792
rect 20404 23780 20410 23792
rect 20990 23780 20996 23792
rect 20404 23752 20996 23780
rect 20404 23740 20410 23752
rect 20990 23740 20996 23752
rect 21048 23740 21054 23792
rect 22940 23789 22968 23820
rect 23474 23808 23480 23820
rect 23532 23848 23538 23860
rect 24854 23848 24860 23860
rect 23532 23820 24860 23848
rect 23532 23808 23538 23820
rect 24854 23808 24860 23820
rect 24912 23808 24918 23860
rect 28166 23848 28172 23860
rect 28127 23820 28172 23848
rect 28166 23808 28172 23820
rect 28224 23808 28230 23860
rect 31754 23848 31760 23860
rect 31220 23820 31760 23848
rect 22925 23783 22983 23789
rect 22925 23749 22937 23783
rect 22971 23749 22983 23783
rect 22925 23743 22983 23749
rect 23768 23752 24900 23780
rect 17773 23715 17831 23721
rect 17644 23684 17689 23712
rect 17644 23672 17650 23684
rect 17773 23681 17785 23715
rect 17819 23681 17831 23715
rect 18230 23712 18236 23724
rect 18191 23684 18236 23712
rect 17773 23675 17831 23681
rect 18230 23672 18236 23684
rect 18288 23672 18294 23724
rect 21174 23672 21180 23724
rect 21232 23712 21238 23724
rect 22373 23715 22431 23721
rect 22373 23712 22385 23715
rect 21232 23684 22385 23712
rect 21232 23672 21238 23684
rect 22373 23681 22385 23684
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 23109 23715 23167 23721
rect 23109 23681 23121 23715
rect 23155 23681 23167 23715
rect 23109 23675 23167 23681
rect 19242 23604 19248 23656
rect 19300 23644 19306 23656
rect 19337 23647 19395 23653
rect 19337 23644 19349 23647
rect 19300 23616 19349 23644
rect 19300 23604 19306 23616
rect 19337 23613 19349 23616
rect 19383 23613 19395 23647
rect 19337 23607 19395 23613
rect 14001 23579 14059 23585
rect 14001 23545 14013 23579
rect 14047 23576 14059 23579
rect 14047 23548 15240 23576
rect 14047 23545 14059 23548
rect 14001 23539 14059 23545
rect 15212 23520 15240 23548
rect 17494 23536 17500 23588
rect 17552 23536 17558 23588
rect 12526 23508 12532 23520
rect 11716 23480 12296 23508
rect 12487 23480 12532 23508
rect 12526 23468 12532 23480
rect 12584 23468 12590 23520
rect 15194 23468 15200 23520
rect 15252 23468 15258 23520
rect 16114 23468 16120 23520
rect 16172 23508 16178 23520
rect 19352 23508 19380 23607
rect 21726 23604 21732 23656
rect 21784 23644 21790 23656
rect 23124 23644 23152 23675
rect 23658 23672 23664 23724
rect 23716 23712 23722 23724
rect 23768 23721 23796 23752
rect 23753 23715 23811 23721
rect 23753 23712 23765 23715
rect 23716 23684 23765 23712
rect 23716 23672 23722 23684
rect 23753 23681 23765 23684
rect 23799 23681 23811 23715
rect 23753 23675 23811 23681
rect 23937 23715 23995 23721
rect 23937 23681 23949 23715
rect 23983 23681 23995 23715
rect 23937 23675 23995 23681
rect 24029 23715 24087 23721
rect 24029 23681 24041 23715
rect 24075 23681 24087 23715
rect 24029 23675 24087 23681
rect 24121 23715 24179 23721
rect 24121 23681 24133 23715
rect 24167 23712 24179 23715
rect 24302 23712 24308 23724
rect 24167 23684 24308 23712
rect 24167 23681 24179 23684
rect 24121 23675 24179 23681
rect 21784 23616 23152 23644
rect 23293 23647 23351 23653
rect 21784 23604 21790 23616
rect 23293 23613 23305 23647
rect 23339 23644 23351 23647
rect 23952 23644 23980 23675
rect 23339 23616 23980 23644
rect 24044 23644 24072 23675
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 24872 23712 24900 23752
rect 26970 23740 26976 23792
rect 27028 23780 27034 23792
rect 27798 23780 27804 23792
rect 27028 23752 27804 23780
rect 27028 23740 27034 23752
rect 27798 23740 27804 23752
rect 27856 23740 27862 23792
rect 31220 23789 31248 23820
rect 31754 23808 31760 23820
rect 31812 23848 31818 23860
rect 32490 23848 32496 23860
rect 31812 23820 32496 23848
rect 31812 23808 31818 23820
rect 32490 23808 32496 23820
rect 32548 23808 32554 23860
rect 33686 23848 33692 23860
rect 32600 23820 33692 23848
rect 31205 23783 31263 23789
rect 31205 23749 31217 23783
rect 31251 23749 31263 23783
rect 31205 23743 31263 23749
rect 25222 23712 25228 23724
rect 24872 23684 25228 23712
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 25497 23721 25503 23724
rect 25388 23715 25446 23721
rect 25388 23712 25400 23715
rect 25332 23684 25400 23712
rect 24210 23644 24216 23656
rect 24044 23616 24216 23644
rect 23339 23613 23351 23616
rect 23293 23607 23351 23613
rect 24210 23604 24216 23616
rect 24268 23604 24274 23656
rect 24320 23576 24348 23672
rect 25038 23604 25044 23656
rect 25096 23644 25102 23656
rect 25332 23644 25360 23684
rect 25388 23681 25400 23684
rect 25434 23681 25446 23715
rect 25388 23675 25446 23681
rect 25488 23715 25503 23721
rect 25488 23681 25500 23715
rect 25488 23675 25503 23681
rect 25497 23672 25503 23675
rect 25555 23672 25561 23724
rect 25613 23715 25671 23721
rect 25613 23681 25625 23715
rect 25659 23712 25671 23715
rect 29546 23712 29552 23724
rect 25659 23681 25682 23712
rect 29507 23684 29552 23712
rect 25613 23675 25682 23681
rect 25096 23616 25360 23644
rect 25654 23644 25682 23675
rect 29546 23672 29552 23684
rect 29604 23672 29610 23724
rect 29730 23672 29736 23724
rect 29788 23712 29794 23724
rect 29825 23715 29883 23721
rect 29825 23712 29837 23715
rect 29788 23684 29837 23712
rect 29788 23672 29794 23684
rect 29825 23681 29837 23684
rect 29871 23681 29883 23715
rect 29825 23675 29883 23681
rect 31389 23715 31447 23721
rect 31389 23681 31401 23715
rect 31435 23712 31447 23715
rect 31478 23712 31484 23724
rect 31435 23684 31484 23712
rect 31435 23681 31447 23684
rect 31389 23675 31447 23681
rect 25774 23644 25780 23656
rect 25654 23616 25780 23644
rect 25096 23604 25102 23616
rect 25774 23604 25780 23616
rect 25832 23644 25838 23656
rect 27154 23644 27160 23656
rect 25832 23616 27160 23644
rect 25832 23604 25838 23616
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 29840 23644 29868 23675
rect 31478 23672 31484 23684
rect 31536 23712 31542 23724
rect 31662 23712 31668 23724
rect 31536 23684 31668 23712
rect 31536 23672 31542 23684
rect 31662 23672 31668 23684
rect 31720 23672 31726 23724
rect 32398 23712 32404 23724
rect 32359 23684 32404 23712
rect 32398 23672 32404 23684
rect 32456 23672 32462 23724
rect 32600 23721 32628 23820
rect 33686 23808 33692 23820
rect 33744 23808 33750 23860
rect 33778 23808 33784 23860
rect 33836 23848 33842 23860
rect 36722 23848 36728 23860
rect 33836 23820 35020 23848
rect 36683 23820 36728 23848
rect 33836 23808 33842 23820
rect 32858 23780 32864 23792
rect 32692 23752 32864 23780
rect 32692 23721 32720 23752
rect 32858 23740 32864 23752
rect 32916 23740 32922 23792
rect 33045 23783 33103 23789
rect 33045 23749 33057 23783
rect 33091 23749 33103 23783
rect 33045 23743 33103 23749
rect 32585 23715 32643 23721
rect 32585 23681 32597 23715
rect 32631 23681 32643 23715
rect 32585 23675 32643 23681
rect 32677 23715 32735 23721
rect 32677 23681 32689 23715
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 32769 23715 32827 23721
rect 32769 23681 32781 23715
rect 32815 23681 32827 23715
rect 33060 23712 33088 23743
rect 34422 23740 34428 23792
rect 34480 23780 34486 23792
rect 34992 23780 35020 23820
rect 36722 23808 36728 23820
rect 36780 23808 36786 23860
rect 35590 23783 35648 23789
rect 35590 23780 35602 23783
rect 34480 23752 34928 23780
rect 34992 23752 35602 23780
rect 34480 23740 34486 23752
rect 34900 23721 34928 23752
rect 35590 23749 35602 23752
rect 35636 23749 35648 23783
rect 35590 23743 35648 23749
rect 34618 23715 34676 23721
rect 34618 23712 34630 23715
rect 33060 23684 34630 23712
rect 32769 23675 32827 23681
rect 34618 23681 34630 23684
rect 34664 23681 34676 23715
rect 34618 23675 34676 23681
rect 34885 23715 34943 23721
rect 34885 23681 34897 23715
rect 34931 23712 34943 23715
rect 35345 23715 35403 23721
rect 35345 23712 35357 23715
rect 34931 23684 35357 23712
rect 34931 23681 34943 23684
rect 34885 23675 34943 23681
rect 35345 23681 35357 23684
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 32122 23644 32128 23656
rect 29840 23616 32128 23644
rect 32122 23604 32128 23616
rect 32180 23644 32186 23656
rect 32692 23644 32720 23675
rect 32180 23616 32720 23644
rect 32180 23604 32186 23616
rect 30466 23576 30472 23588
rect 24320 23548 30472 23576
rect 30466 23536 30472 23548
rect 30524 23536 30530 23588
rect 32214 23576 32220 23588
rect 30576 23548 32220 23576
rect 21174 23508 21180 23520
rect 16172 23480 19380 23508
rect 21135 23480 21180 23508
rect 16172 23468 16178 23480
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 24397 23511 24455 23517
rect 24397 23477 24409 23511
rect 24443 23508 24455 23511
rect 25682 23508 25688 23520
rect 24443 23480 25688 23508
rect 24443 23477 24455 23480
rect 24397 23471 24455 23477
rect 25682 23468 25688 23480
rect 25740 23468 25746 23520
rect 25869 23511 25927 23517
rect 25869 23477 25881 23511
rect 25915 23508 25927 23511
rect 27062 23508 27068 23520
rect 25915 23480 27068 23508
rect 25915 23477 25927 23480
rect 25869 23471 25927 23477
rect 27062 23468 27068 23480
rect 27120 23468 27126 23520
rect 27154 23468 27160 23520
rect 27212 23508 27218 23520
rect 27798 23508 27804 23520
rect 27212 23480 27804 23508
rect 27212 23468 27218 23480
rect 27798 23468 27804 23480
rect 27856 23508 27862 23520
rect 30576 23508 30604 23548
rect 32214 23536 32220 23548
rect 32272 23576 32278 23588
rect 32784 23576 32812 23675
rect 32272 23548 32812 23576
rect 32272 23536 32278 23548
rect 27856 23480 30604 23508
rect 31573 23511 31631 23517
rect 27856 23468 27862 23480
rect 31573 23477 31585 23511
rect 31619 23508 31631 23511
rect 32398 23508 32404 23520
rect 31619 23480 32404 23508
rect 31619 23477 31631 23480
rect 31573 23471 31631 23477
rect 32398 23468 32404 23480
rect 32456 23468 32462 23520
rect 32582 23468 32588 23520
rect 32640 23508 32646 23520
rect 32766 23508 32772 23520
rect 32640 23480 32772 23508
rect 32640 23468 32646 23480
rect 32766 23468 32772 23480
rect 32824 23468 32830 23520
rect 33410 23468 33416 23520
rect 33468 23508 33474 23520
rect 33505 23511 33563 23517
rect 33505 23508 33517 23511
rect 33468 23480 33517 23508
rect 33468 23468 33474 23480
rect 33505 23477 33517 23480
rect 33551 23477 33563 23511
rect 33505 23471 33563 23477
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 5626 23304 5632 23316
rect 5587 23276 5632 23304
rect 5626 23264 5632 23276
rect 5684 23264 5690 23316
rect 6365 23307 6423 23313
rect 6365 23273 6377 23307
rect 6411 23304 6423 23307
rect 7466 23304 7472 23316
rect 6411 23276 7472 23304
rect 6411 23273 6423 23276
rect 6365 23267 6423 23273
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 11517 23307 11575 23313
rect 11517 23273 11529 23307
rect 11563 23304 11575 23307
rect 12066 23304 12072 23316
rect 11563 23276 12072 23304
rect 11563 23273 11575 23276
rect 11517 23267 11575 23273
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 16666 23304 16672 23316
rect 14608 23276 16672 23304
rect 14608 23264 14614 23276
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 16850 23264 16856 23316
rect 16908 23304 16914 23316
rect 17770 23304 17776 23316
rect 16908 23276 17776 23304
rect 16908 23264 16914 23276
rect 17770 23264 17776 23276
rect 17828 23304 17834 23316
rect 19150 23304 19156 23316
rect 17828 23276 19156 23304
rect 17828 23264 17834 23276
rect 19150 23264 19156 23276
rect 19208 23304 19214 23316
rect 19334 23304 19340 23316
rect 19208 23276 19340 23304
rect 19208 23264 19214 23276
rect 19334 23264 19340 23276
rect 19392 23304 19398 23316
rect 21082 23304 21088 23316
rect 19392 23276 19485 23304
rect 21043 23276 21088 23304
rect 19392 23264 19398 23276
rect 21082 23264 21088 23276
rect 21140 23264 21146 23316
rect 21910 23304 21916 23316
rect 21871 23276 21916 23304
rect 21910 23264 21916 23276
rect 21968 23304 21974 23316
rect 22922 23304 22928 23316
rect 21968 23276 22928 23304
rect 21968 23264 21974 23276
rect 22922 23264 22928 23276
rect 22980 23264 22986 23316
rect 25038 23264 25044 23316
rect 25096 23304 25102 23316
rect 25225 23307 25283 23313
rect 25225 23304 25237 23307
rect 25096 23276 25237 23304
rect 25096 23264 25102 23276
rect 25225 23273 25237 23276
rect 25271 23273 25283 23307
rect 28902 23304 28908 23316
rect 25225 23267 25283 23273
rect 25516 23276 27936 23304
rect 28863 23276 28908 23304
rect 6822 23196 6828 23248
rect 6880 23236 6886 23248
rect 6880 23208 7696 23236
rect 6880 23196 6886 23208
rect 3326 23168 3332 23180
rect 2148 23140 3332 23168
rect 1578 23060 1584 23112
rect 1636 23100 1642 23112
rect 2148 23109 2176 23140
rect 3326 23128 3332 23140
rect 3384 23128 3390 23180
rect 3786 23128 3792 23180
rect 3844 23168 3850 23180
rect 4249 23171 4307 23177
rect 4249 23168 4261 23171
rect 3844 23140 4261 23168
rect 3844 23128 3850 23140
rect 4249 23137 4261 23140
rect 4295 23137 4307 23171
rect 7374 23168 7380 23180
rect 4249 23131 4307 23137
rect 6748 23140 7380 23168
rect 2133 23103 2191 23109
rect 2133 23100 2145 23103
rect 1636 23072 2145 23100
rect 1636 23060 1642 23072
rect 2133 23069 2145 23072
rect 2179 23069 2191 23103
rect 2314 23100 2320 23112
rect 2275 23072 2320 23100
rect 2133 23063 2191 23069
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23069 2467 23103
rect 2409 23063 2467 23069
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23100 2559 23103
rect 2958 23100 2964 23112
rect 2547 23072 2964 23100
rect 2547 23069 2559 23072
rect 2501 23063 2559 23069
rect 2424 23032 2452 23063
rect 2958 23060 2964 23072
rect 3016 23060 3022 23112
rect 5534 23060 5540 23112
rect 5592 23100 5598 23112
rect 5718 23100 5724 23112
rect 5592 23072 5724 23100
rect 5592 23060 5598 23072
rect 5718 23060 5724 23072
rect 5776 23100 5782 23112
rect 6748 23109 6776 23140
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 6641 23103 6699 23109
rect 6641 23100 6653 23103
rect 5776 23072 6653 23100
rect 5776 23060 5782 23072
rect 6641 23069 6653 23072
rect 6687 23069 6699 23103
rect 6641 23063 6699 23069
rect 6733 23103 6791 23109
rect 6733 23069 6745 23103
rect 6779 23069 6791 23103
rect 6733 23063 6791 23069
rect 6825 23103 6883 23109
rect 6825 23069 6837 23103
rect 6871 23100 6883 23103
rect 6914 23100 6920 23112
rect 6871 23072 6920 23100
rect 6871 23069 6883 23072
rect 6825 23063 6883 23069
rect 6914 23060 6920 23072
rect 6972 23060 6978 23112
rect 7006 23060 7012 23112
rect 7064 23100 7070 23112
rect 7466 23100 7472 23112
rect 7064 23072 7472 23100
rect 7064 23060 7070 23072
rect 7466 23060 7472 23072
rect 7524 23060 7530 23112
rect 7668 23109 7696 23208
rect 7742 23196 7748 23248
rect 7800 23236 7806 23248
rect 9033 23239 9091 23245
rect 9033 23236 9045 23239
rect 7800 23208 9045 23236
rect 7800 23196 7806 23208
rect 9033 23205 9045 23208
rect 9079 23205 9091 23239
rect 14458 23236 14464 23248
rect 9033 23199 9091 23205
rect 10980 23208 14464 23236
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 8036 23140 9689 23168
rect 8036 23112 8064 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 10134 23128 10140 23180
rect 10192 23168 10198 23180
rect 10192 23140 10824 23168
rect 10192 23128 10198 23140
rect 7653 23103 7711 23109
rect 7653 23069 7665 23103
rect 7699 23069 7711 23103
rect 7653 23063 7711 23069
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23069 7803 23103
rect 7745 23063 7803 23069
rect 2682 23032 2688 23044
rect 2424 23004 2688 23032
rect 2682 22992 2688 23004
rect 2740 22992 2746 23044
rect 2777 23035 2835 23041
rect 2777 23001 2789 23035
rect 2823 23032 2835 23035
rect 4494 23035 4552 23041
rect 4494 23032 4506 23035
rect 2823 23004 4506 23032
rect 2823 23001 2835 23004
rect 2777 22995 2835 23001
rect 4494 23001 4506 23004
rect 4540 23001 4552 23035
rect 4494 22995 4552 23001
rect 4614 22992 4620 23044
rect 4672 23032 4678 23044
rect 4672 23004 5764 23032
rect 4672 22992 4678 23004
rect 2498 22924 2504 22976
rect 2556 22964 2562 22976
rect 5442 22964 5448 22976
rect 2556 22936 5448 22964
rect 2556 22924 2562 22936
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 5736 22964 5764 23004
rect 7098 22992 7104 23044
rect 7156 23032 7162 23044
rect 7760 23032 7788 23063
rect 7834 23060 7840 23112
rect 7892 23100 7898 23112
rect 8018 23100 8024 23112
rect 7892 23072 8024 23100
rect 7892 23060 7898 23072
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8904 23072 8953 23100
rect 8904 23060 8910 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9490 23100 9496 23112
rect 9171 23072 9496 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9490 23060 9496 23072
rect 9548 23060 9554 23112
rect 10594 23100 10600 23112
rect 10555 23072 10600 23100
rect 10594 23060 10600 23072
rect 10652 23060 10658 23112
rect 10796 23041 10824 23140
rect 10980 23109 11008 23208
rect 14458 23196 14464 23208
rect 14516 23196 14522 23248
rect 21174 23236 21180 23248
rect 17144 23208 21180 23236
rect 12986 23168 12992 23180
rect 12947 23140 12992 23168
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23168 15531 23171
rect 16114 23168 16120 23180
rect 15519 23140 16120 23168
rect 15519 23137 15531 23140
rect 15473 23131 15531 23137
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 10965 23103 11023 23109
rect 10965 23069 10977 23103
rect 11011 23069 11023 23103
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 10965 23063 11023 23069
rect 11072 23072 12725 23100
rect 10689 23035 10747 23041
rect 10689 23032 10701 23035
rect 7156 23004 7788 23032
rect 7852 23004 10701 23032
rect 7156 22992 7162 23004
rect 7852 22964 7880 23004
rect 10689 23001 10701 23004
rect 10735 23001 10747 23035
rect 10689 22995 10747 23001
rect 10781 23035 10839 23041
rect 10781 23001 10793 23035
rect 10827 23032 10839 23035
rect 11072 23032 11100 23072
rect 12713 23069 12725 23072
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 15194 23060 15200 23112
rect 15252 23109 15258 23112
rect 15252 23100 15264 23109
rect 15252 23072 15297 23100
rect 15252 23063 15264 23072
rect 15252 23060 15258 23063
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17037 23103 17095 23109
rect 17037 23100 17049 23103
rect 16816 23072 17049 23100
rect 16816 23060 16822 23072
rect 17037 23069 17049 23072
rect 17083 23069 17095 23103
rect 17037 23063 17095 23069
rect 10827 23004 11100 23032
rect 10827 23001 10839 23004
rect 10781 22995 10839 23001
rect 11514 22992 11520 23044
rect 11572 23032 11578 23044
rect 11609 23035 11667 23041
rect 11609 23032 11621 23035
rect 11572 23004 11621 23032
rect 11572 22992 11578 23004
rect 11609 23001 11621 23004
rect 11655 23032 11667 23035
rect 11655 23004 14964 23032
rect 11655 23001 11667 23004
rect 11609 22995 11667 23001
rect 5736 22936 7880 22964
rect 8113 22967 8171 22973
rect 8113 22933 8125 22967
rect 8159 22964 8171 22967
rect 8202 22964 8208 22976
rect 8159 22936 8208 22964
rect 8159 22933 8171 22936
rect 8113 22927 8171 22933
rect 8202 22924 8208 22936
rect 8260 22924 8266 22976
rect 10413 22967 10471 22973
rect 10413 22933 10425 22967
rect 10459 22964 10471 22967
rect 13262 22964 13268 22976
rect 10459 22936 13268 22964
rect 10459 22933 10471 22936
rect 10413 22927 10471 22933
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 13354 22924 13360 22976
rect 13412 22964 13418 22976
rect 14093 22967 14151 22973
rect 14093 22964 14105 22967
rect 13412 22936 14105 22964
rect 13412 22924 13418 22936
rect 14093 22933 14105 22936
rect 14139 22933 14151 22967
rect 14936 22964 14964 23004
rect 17144 22964 17172 23208
rect 21174 23196 21180 23208
rect 21232 23196 21238 23248
rect 23198 23196 23204 23248
rect 23256 23236 23262 23248
rect 23293 23239 23351 23245
rect 23293 23236 23305 23239
rect 23256 23208 23305 23236
rect 23256 23196 23262 23208
rect 23293 23205 23305 23208
rect 23339 23236 23351 23239
rect 25516 23236 25544 23276
rect 23339 23208 25544 23236
rect 27908 23236 27936 23276
rect 28902 23264 28908 23276
rect 28960 23264 28966 23316
rect 29917 23307 29975 23313
rect 29917 23273 29929 23307
rect 29963 23304 29975 23307
rect 30282 23304 30288 23316
rect 29963 23276 30288 23304
rect 29963 23273 29975 23276
rect 29917 23267 29975 23273
rect 30282 23264 30288 23276
rect 30340 23264 30346 23316
rect 33686 23304 33692 23316
rect 33647 23276 33692 23304
rect 33686 23264 33692 23276
rect 33744 23264 33750 23316
rect 32861 23239 32919 23245
rect 27908 23208 28856 23236
rect 23339 23205 23351 23208
rect 23293 23199 23351 23205
rect 17494 23168 17500 23180
rect 17328 23140 17500 23168
rect 17328 23109 17356 23140
rect 17494 23128 17500 23140
rect 17552 23128 17558 23180
rect 20257 23171 20315 23177
rect 20257 23137 20269 23171
rect 20303 23168 20315 23171
rect 20303 23140 21772 23168
rect 20303 23137 20315 23140
rect 20257 23131 20315 23137
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 17313 23103 17371 23109
rect 17313 23069 17325 23103
rect 17359 23069 17371 23103
rect 17313 23063 17371 23069
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23100 17463 23103
rect 17586 23100 17592 23112
rect 17451 23072 17592 23100
rect 17451 23069 17463 23072
rect 17405 23063 17463 23069
rect 17236 23032 17264 23063
rect 17586 23060 17592 23072
rect 17644 23060 17650 23112
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 18288 23072 18521 23100
rect 18288 23060 18294 23072
rect 18509 23069 18521 23072
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 20622 23060 20628 23112
rect 20680 23100 20686 23112
rect 20717 23103 20775 23109
rect 20717 23100 20729 23103
rect 20680 23072 20729 23100
rect 20680 23060 20686 23072
rect 20717 23069 20729 23072
rect 20763 23069 20775 23103
rect 20898 23100 20904 23112
rect 20859 23072 20904 23100
rect 20717 23063 20775 23069
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 21266 23060 21272 23112
rect 21324 23100 21330 23112
rect 21744 23109 21772 23140
rect 25498 23128 25504 23180
rect 25556 23168 25562 23180
rect 25685 23171 25743 23177
rect 25685 23168 25697 23171
rect 25556 23140 25697 23168
rect 25556 23128 25562 23140
rect 25685 23137 25697 23140
rect 25731 23168 25743 23171
rect 25774 23168 25780 23180
rect 25731 23140 25780 23168
rect 25731 23137 25743 23140
rect 25685 23131 25743 23137
rect 25774 23128 25780 23140
rect 25832 23128 25838 23180
rect 26970 23168 26976 23180
rect 26931 23140 26976 23168
rect 26970 23128 26976 23140
rect 27028 23128 27034 23180
rect 21545 23103 21603 23109
rect 21545 23100 21557 23103
rect 21324 23072 21557 23100
rect 21324 23060 21330 23072
rect 21545 23069 21557 23072
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22094 23100 22100 23112
rect 21775 23072 22100 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 22094 23060 22100 23072
rect 22152 23060 22158 23112
rect 23014 23060 23020 23112
rect 23072 23100 23078 23112
rect 23290 23100 23296 23112
rect 23072 23072 23296 23100
rect 23072 23060 23078 23072
rect 23290 23060 23296 23072
rect 23348 23060 23354 23112
rect 24854 23100 24860 23112
rect 24815 23072 24860 23100
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 27062 23060 27068 23112
rect 27120 23100 27126 23112
rect 28828 23109 28856 23208
rect 32861 23205 32873 23239
rect 32907 23236 32919 23239
rect 33778 23236 33784 23248
rect 32907 23208 33784 23236
rect 32907 23205 32919 23208
rect 32861 23199 32919 23205
rect 33778 23196 33784 23208
rect 33836 23196 33842 23248
rect 31757 23171 31815 23177
rect 29012 23140 29776 23168
rect 29012 23109 29040 23140
rect 27229 23103 27287 23109
rect 27229 23100 27241 23103
rect 27120 23072 27241 23100
rect 27120 23060 27126 23072
rect 27229 23069 27241 23072
rect 27275 23069 27287 23103
rect 27229 23063 27287 23069
rect 28813 23103 28871 23109
rect 28813 23069 28825 23103
rect 28859 23069 28871 23103
rect 28813 23063 28871 23069
rect 28997 23103 29055 23109
rect 28997 23069 29009 23103
rect 29043 23069 29055 23103
rect 29546 23100 29552 23112
rect 29507 23072 29552 23100
rect 28997 23063 29055 23069
rect 29546 23060 29552 23072
rect 29604 23060 29610 23112
rect 29748 23109 29776 23140
rect 31757 23137 31769 23171
rect 31803 23168 31815 23171
rect 31938 23168 31944 23180
rect 31803 23140 31944 23168
rect 31803 23137 31815 23140
rect 31757 23131 31815 23137
rect 31938 23128 31944 23140
rect 31996 23128 32002 23180
rect 29733 23103 29791 23109
rect 29733 23069 29745 23103
rect 29779 23100 29791 23103
rect 29914 23100 29920 23112
rect 29779 23072 29920 23100
rect 29779 23069 29791 23072
rect 29733 23063 29791 23069
rect 29914 23060 29920 23072
rect 29972 23060 29978 23112
rect 32214 23100 32220 23112
rect 32175 23072 32220 23100
rect 32214 23060 32220 23072
rect 32272 23060 32278 23112
rect 32398 23109 32404 23112
rect 32396 23100 32404 23109
rect 32359 23072 32404 23100
rect 32396 23063 32404 23072
rect 32398 23060 32404 23063
rect 32456 23060 32462 23112
rect 32496 23100 32554 23106
rect 32496 23066 32508 23100
rect 32542 23066 32554 23100
rect 32496 23060 32554 23066
rect 32582 23060 32588 23112
rect 32640 23100 32646 23112
rect 32640 23072 32685 23100
rect 32640 23060 32646 23072
rect 32766 23060 32772 23112
rect 32824 23100 32830 23112
rect 33321 23103 33379 23109
rect 33321 23100 33333 23103
rect 32824 23072 33333 23100
rect 32824 23060 32830 23072
rect 33321 23069 33333 23072
rect 33367 23069 33379 23103
rect 33321 23063 33379 23069
rect 18141 23035 18199 23041
rect 18141 23032 18153 23035
rect 17236 23004 18153 23032
rect 18141 23001 18153 23004
rect 18187 23001 18199 23035
rect 18322 23032 18328 23044
rect 18283 23004 18328 23032
rect 18141 22995 18199 23001
rect 18322 22992 18328 23004
rect 18380 22992 18386 23044
rect 21174 22992 21180 23044
rect 21232 23032 21238 23044
rect 21358 23032 21364 23044
rect 21232 23004 21364 23032
rect 21232 22992 21238 23004
rect 21358 22992 21364 23004
rect 21416 23032 21422 23044
rect 22002 23032 22008 23044
rect 21416 23004 22008 23032
rect 21416 22992 21422 23004
rect 22002 22992 22008 23004
rect 22060 23032 22066 23044
rect 22649 23035 22707 23041
rect 22649 23032 22661 23035
rect 22060 23004 22661 23032
rect 22060 22992 22066 23004
rect 22649 23001 22661 23004
rect 22695 23001 22707 23035
rect 23474 23032 23480 23044
rect 23435 23004 23480 23032
rect 22649 22995 22707 23001
rect 23474 22992 23480 23004
rect 23532 22992 23538 23044
rect 25041 23035 25099 23041
rect 25041 23001 25053 23035
rect 25087 23032 25099 23035
rect 25087 23004 28396 23032
rect 25087 23001 25099 23004
rect 25041 22995 25099 23001
rect 17678 22964 17684 22976
rect 14936 22936 17172 22964
rect 17639 22936 17684 22964
rect 14093 22927 14151 22933
rect 17678 22924 17684 22936
rect 17736 22924 17742 22976
rect 22738 22964 22744 22976
rect 22651 22936 22744 22964
rect 22738 22924 22744 22936
rect 22796 22964 22802 22976
rect 23658 22964 23664 22976
rect 22796 22936 23664 22964
rect 22796 22924 22802 22936
rect 23658 22924 23664 22936
rect 23716 22924 23722 22976
rect 24762 22924 24768 22976
rect 24820 22964 24826 22976
rect 25056 22964 25084 22995
rect 28368 22973 28396 23004
rect 30650 22992 30656 23044
rect 30708 23032 30714 23044
rect 31490 23035 31548 23041
rect 31490 23032 31502 23035
rect 30708 23004 31502 23032
rect 30708 22992 30714 23004
rect 31490 23001 31502 23004
rect 31536 23001 31548 23035
rect 31490 22995 31548 23001
rect 32122 22992 32128 23044
rect 32180 23032 32186 23044
rect 32508 23032 32536 23060
rect 32180 23004 32536 23032
rect 32180 22992 32186 23004
rect 33410 22992 33416 23044
rect 33468 23032 33474 23044
rect 33505 23035 33563 23041
rect 33505 23032 33517 23035
rect 33468 23004 33517 23032
rect 33468 22992 33474 23004
rect 33505 23001 33517 23004
rect 33551 23001 33563 23035
rect 33505 22995 33563 23001
rect 24820 22936 25084 22964
rect 28353 22967 28411 22973
rect 24820 22924 24826 22936
rect 28353 22933 28365 22967
rect 28399 22933 28411 22967
rect 28353 22927 28411 22933
rect 30098 22924 30104 22976
rect 30156 22964 30162 22976
rect 30377 22967 30435 22973
rect 30377 22964 30389 22967
rect 30156 22936 30389 22964
rect 30156 22924 30162 22936
rect 30377 22933 30389 22936
rect 30423 22933 30435 22967
rect 30377 22927 30435 22933
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 2501 22763 2559 22769
rect 2501 22729 2513 22763
rect 2547 22760 2559 22763
rect 3970 22760 3976 22772
rect 2547 22732 3976 22760
rect 2547 22729 2559 22732
rect 2501 22723 2559 22729
rect 3970 22720 3976 22732
rect 4028 22720 4034 22772
rect 4525 22763 4583 22769
rect 4525 22729 4537 22763
rect 4571 22760 4583 22763
rect 4614 22760 4620 22772
rect 4571 22732 4620 22760
rect 4571 22729 4583 22732
rect 4525 22723 4583 22729
rect 4614 22720 4620 22732
rect 4672 22720 4678 22772
rect 5442 22760 5448 22772
rect 5403 22732 5448 22760
rect 5442 22720 5448 22732
rect 5500 22720 5506 22772
rect 13538 22760 13544 22772
rect 11992 22732 12434 22760
rect 13499 22732 13544 22760
rect 3786 22692 3792 22704
rect 3160 22664 3792 22692
rect 2130 22624 2136 22636
rect 2091 22596 2136 22624
rect 2130 22584 2136 22596
rect 2188 22584 2194 22636
rect 3160 22633 3188 22664
rect 3786 22652 3792 22664
rect 3844 22652 3850 22704
rect 2317 22627 2375 22633
rect 2317 22593 2329 22627
rect 2363 22593 2375 22627
rect 2317 22587 2375 22593
rect 3145 22627 3203 22633
rect 3145 22593 3157 22627
rect 3191 22593 3203 22627
rect 3145 22587 3203 22593
rect 2332 22420 2360 22587
rect 3234 22584 3240 22636
rect 3292 22624 3298 22636
rect 3401 22627 3459 22633
rect 3401 22624 3413 22627
rect 3292 22596 3413 22624
rect 3292 22584 3298 22596
rect 3401 22593 3413 22596
rect 3447 22593 3459 22627
rect 3401 22587 3459 22593
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22593 5687 22627
rect 5629 22587 5687 22593
rect 5644 22488 5672 22587
rect 6730 22584 6736 22636
rect 6788 22624 6794 22636
rect 8202 22633 8208 22636
rect 7929 22627 7987 22633
rect 7929 22624 7941 22627
rect 6788 22596 7941 22624
rect 6788 22584 6794 22596
rect 7929 22593 7941 22596
rect 7975 22593 7987 22627
rect 8196 22624 8208 22633
rect 8163 22596 8208 22624
rect 7929 22587 7987 22593
rect 8196 22587 8208 22596
rect 8202 22584 8208 22587
rect 8260 22584 8266 22636
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 10652 22596 10701 22624
rect 10652 22584 10658 22596
rect 10689 22593 10701 22596
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 11146 22584 11152 22636
rect 11204 22624 11210 22636
rect 11992 22633 12020 22732
rect 12158 22692 12164 22704
rect 12119 22664 12164 22692
rect 12158 22652 12164 22664
rect 12216 22652 12222 22704
rect 12406 22692 12434 22732
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 17586 22720 17592 22772
rect 17644 22720 17650 22772
rect 18138 22760 18144 22772
rect 18051 22732 18144 22760
rect 18138 22720 18144 22732
rect 18196 22760 18202 22772
rect 18322 22760 18328 22772
rect 18196 22732 18328 22760
rect 18196 22720 18202 22732
rect 18322 22720 18328 22732
rect 18380 22720 18386 22772
rect 21266 22720 21272 22772
rect 21324 22760 21330 22772
rect 29365 22763 29423 22769
rect 29365 22760 29377 22763
rect 21324 22732 29377 22760
rect 21324 22720 21330 22732
rect 29365 22729 29377 22732
rect 29411 22760 29423 22763
rect 29546 22760 29552 22772
rect 29411 22732 29552 22760
rect 29411 22729 29423 22732
rect 29365 22723 29423 22729
rect 29546 22720 29552 22732
rect 29604 22720 29610 22772
rect 30466 22720 30472 22772
rect 30524 22760 30530 22772
rect 31481 22763 31539 22769
rect 31481 22760 31493 22763
rect 30524 22732 31493 22760
rect 30524 22720 30530 22732
rect 31481 22729 31493 22732
rect 31527 22760 31539 22763
rect 32582 22760 32588 22772
rect 31527 22732 32588 22760
rect 31527 22729 31539 22732
rect 31481 22723 31539 22729
rect 32582 22720 32588 22732
rect 32640 22720 32646 22772
rect 13170 22692 13176 22704
rect 12406 22664 13032 22692
rect 13131 22664 13176 22692
rect 11885 22627 11943 22633
rect 11885 22624 11897 22627
rect 11204 22596 11897 22624
rect 11204 22584 11210 22596
rect 11885 22593 11897 22596
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 11978 22627 12036 22633
rect 11978 22593 11990 22627
rect 12024 22593 12036 22627
rect 11978 22587 12036 22593
rect 12253 22627 12311 22633
rect 12253 22593 12265 22627
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 5813 22559 5871 22565
rect 5813 22525 5825 22559
rect 5859 22556 5871 22559
rect 5902 22556 5908 22568
rect 5859 22528 5908 22556
rect 5859 22525 5871 22528
rect 5813 22519 5871 22525
rect 5902 22516 5908 22528
rect 5960 22516 5966 22568
rect 7098 22516 7104 22568
rect 7156 22556 7162 22568
rect 7193 22559 7251 22565
rect 7193 22556 7205 22559
rect 7156 22528 7205 22556
rect 7156 22516 7162 22528
rect 7193 22525 7205 22528
rect 7239 22525 7251 22559
rect 7193 22519 7251 22525
rect 7469 22559 7527 22565
rect 7469 22525 7481 22559
rect 7515 22556 7527 22559
rect 7558 22556 7564 22568
rect 7515 22528 7564 22556
rect 7515 22525 7527 22528
rect 7469 22519 7527 22525
rect 7558 22516 7564 22528
rect 7616 22556 7622 22568
rect 7742 22556 7748 22568
rect 7616 22528 7748 22556
rect 7616 22516 7622 22528
rect 7742 22516 7748 22528
rect 7800 22516 7806 22568
rect 10962 22556 10968 22568
rect 10923 22528 10968 22556
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 7926 22488 7932 22500
rect 5644 22460 7932 22488
rect 7926 22448 7932 22460
rect 7984 22448 7990 22500
rect 9306 22488 9312 22500
rect 9219 22460 9312 22488
rect 9306 22448 9312 22460
rect 9364 22488 9370 22500
rect 12268 22488 12296 22587
rect 12342 22584 12348 22636
rect 12400 22633 12406 22636
rect 12400 22624 12408 22633
rect 12400 22596 12445 22624
rect 12400 22587 12408 22596
rect 12400 22584 12406 22587
rect 13004 22556 13032 22664
rect 13170 22652 13176 22664
rect 13228 22652 13234 22704
rect 13354 22692 13360 22704
rect 13315 22664 13360 22692
rect 13354 22652 13360 22664
rect 13412 22652 13418 22704
rect 13446 22652 13452 22704
rect 13504 22692 13510 22704
rect 17604 22692 17632 22720
rect 13504 22664 17632 22692
rect 13504 22652 13510 22664
rect 17678 22652 17684 22704
rect 17736 22692 17742 22704
rect 19254 22695 19312 22701
rect 19254 22692 19266 22695
rect 17736 22664 19266 22692
rect 17736 22652 17742 22664
rect 19254 22661 19266 22664
rect 19300 22661 19312 22695
rect 22002 22692 22008 22704
rect 21963 22664 22008 22692
rect 19254 22655 19312 22661
rect 22002 22652 22008 22664
rect 22060 22652 22066 22704
rect 30098 22652 30104 22704
rect 30156 22692 30162 22704
rect 30745 22695 30803 22701
rect 30745 22692 30757 22695
rect 30156 22664 30757 22692
rect 30156 22652 30162 22664
rect 30745 22661 30757 22664
rect 30791 22661 30803 22695
rect 32493 22695 32551 22701
rect 32493 22692 32505 22695
rect 30745 22655 30803 22661
rect 31726 22664 32505 22692
rect 31726 22636 31754 22664
rect 32493 22661 32505 22664
rect 32539 22661 32551 22695
rect 32493 22655 32551 22661
rect 14185 22627 14243 22633
rect 14185 22593 14197 22627
rect 14231 22624 14243 22627
rect 15470 22624 15476 22636
rect 14231 22596 15476 22624
rect 14231 22593 14243 22596
rect 14185 22587 14243 22593
rect 15470 22584 15476 22596
rect 15528 22624 15534 22636
rect 17402 22624 17408 22636
rect 15528 22596 17408 22624
rect 15528 22584 15534 22596
rect 17402 22584 17408 22596
rect 17460 22624 17466 22636
rect 17589 22627 17647 22633
rect 17589 22624 17601 22627
rect 17460 22596 17601 22624
rect 17460 22584 17466 22596
rect 17589 22593 17601 22596
rect 17635 22624 17647 22627
rect 20438 22624 20444 22636
rect 17635 22596 20444 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 20438 22584 20444 22596
rect 20496 22584 20502 22636
rect 20806 22584 20812 22636
rect 20864 22624 20870 22636
rect 24305 22627 24363 22633
rect 24305 22624 24317 22627
rect 20864 22596 24317 22624
rect 20864 22584 20870 22596
rect 24305 22593 24317 22596
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 24394 22584 24400 22636
rect 24452 22624 24458 22636
rect 24581 22627 24639 22633
rect 24452 22596 24497 22624
rect 24452 22584 24458 22596
rect 24581 22593 24593 22627
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 24673 22627 24731 22633
rect 24673 22593 24685 22627
rect 24719 22593 24731 22627
rect 24673 22587 24731 22593
rect 24811 22627 24869 22633
rect 24811 22593 24823 22627
rect 24857 22624 24869 22627
rect 24946 22624 24952 22636
rect 24857 22596 24952 22624
rect 24857 22593 24869 22596
rect 24811 22587 24869 22593
rect 16298 22556 16304 22568
rect 13004 22528 16304 22556
rect 16298 22516 16304 22528
rect 16356 22516 16362 22568
rect 19521 22559 19579 22565
rect 19521 22525 19533 22559
rect 19567 22556 19579 22559
rect 22002 22556 22008 22568
rect 19567 22528 22008 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 22002 22516 22008 22528
rect 22060 22516 22066 22568
rect 23198 22516 23204 22568
rect 23256 22556 23262 22568
rect 23293 22559 23351 22565
rect 23293 22556 23305 22559
rect 23256 22528 23305 22556
rect 23256 22516 23262 22528
rect 23293 22525 23305 22528
rect 23339 22525 23351 22559
rect 23293 22519 23351 22525
rect 9364 22460 12296 22488
rect 12529 22491 12587 22497
rect 9364 22448 9370 22460
rect 12529 22457 12541 22491
rect 12575 22488 12587 22491
rect 16390 22488 16396 22500
rect 12575 22460 16396 22488
rect 12575 22457 12587 22460
rect 12529 22451 12587 22457
rect 16390 22448 16396 22460
rect 16448 22448 16454 22500
rect 21269 22491 21327 22497
rect 21269 22457 21281 22491
rect 21315 22488 21327 22491
rect 22094 22488 22100 22500
rect 21315 22460 22100 22488
rect 21315 22457 21327 22460
rect 21269 22451 21327 22457
rect 22094 22448 22100 22460
rect 22152 22488 22158 22500
rect 23216 22488 23244 22516
rect 23566 22488 23572 22500
rect 22152 22460 23244 22488
rect 23400 22460 23572 22488
rect 22152 22448 22158 22460
rect 5166 22420 5172 22432
rect 2332 22392 5172 22420
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 7944 22420 7972 22448
rect 8110 22420 8116 22432
rect 7944 22392 8116 22420
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 13262 22380 13268 22432
rect 13320 22420 13326 22432
rect 15930 22420 15936 22432
rect 13320 22392 15936 22420
rect 13320 22380 13326 22392
rect 15930 22380 15936 22392
rect 15988 22380 15994 22432
rect 20622 22420 20628 22432
rect 20583 22392 20628 22420
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 23063 22423 23121 22429
rect 23063 22389 23075 22423
rect 23109 22420 23121 22423
rect 23400 22420 23428 22460
rect 23566 22448 23572 22460
rect 23624 22488 23630 22500
rect 24596 22488 24624 22587
rect 24688 22556 24716 22587
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 30561 22627 30619 22633
rect 30561 22593 30573 22627
rect 30607 22624 30619 22627
rect 31662 22624 31668 22636
rect 30607 22596 31668 22624
rect 30607 22593 30619 22596
rect 30561 22587 30619 22593
rect 31662 22584 31668 22596
rect 31720 22596 31754 22636
rect 32309 22627 32367 22633
rect 31720 22584 31726 22596
rect 32309 22593 32321 22627
rect 32355 22624 32367 22627
rect 33502 22624 33508 22636
rect 32355 22596 33508 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 32324 22556 32352 22587
rect 33502 22584 33508 22596
rect 33560 22584 33566 22636
rect 37277 22627 37335 22633
rect 37277 22593 37289 22627
rect 37323 22624 37335 22627
rect 37366 22624 37372 22636
rect 37323 22596 37372 22624
rect 37323 22593 37335 22596
rect 37277 22587 37335 22593
rect 37366 22584 37372 22596
rect 37424 22584 37430 22636
rect 37550 22633 37556 22636
rect 37544 22587 37556 22633
rect 37608 22624 37614 22636
rect 37608 22596 37644 22624
rect 37550 22584 37556 22587
rect 37608 22584 37614 22596
rect 24688 22528 32352 22556
rect 24670 22488 24676 22500
rect 23624 22460 24676 22488
rect 23624 22448 23630 22460
rect 24670 22448 24676 22460
rect 24728 22448 24734 22500
rect 67634 22488 67640 22500
rect 67595 22460 67640 22488
rect 67634 22448 67640 22460
rect 67692 22448 67698 22500
rect 23109 22392 23428 22420
rect 23109 22389 23121 22392
rect 23063 22383 23121 22389
rect 23474 22380 23480 22432
rect 23532 22420 23538 22432
rect 23753 22423 23811 22429
rect 23753 22420 23765 22423
rect 23532 22392 23765 22420
rect 23532 22380 23538 22392
rect 23753 22389 23765 22392
rect 23799 22389 23811 22423
rect 23753 22383 23811 22389
rect 24854 22380 24860 22432
rect 24912 22420 24918 22432
rect 24949 22423 25007 22429
rect 24949 22420 24961 22423
rect 24912 22392 24961 22420
rect 24912 22380 24918 22392
rect 24949 22389 24961 22392
rect 24995 22389 25007 22423
rect 24949 22383 25007 22389
rect 30929 22423 30987 22429
rect 30929 22389 30941 22423
rect 30975 22420 30987 22423
rect 31110 22420 31116 22432
rect 30975 22392 31116 22420
rect 30975 22389 30987 22392
rect 30929 22383 30987 22389
rect 31110 22380 31116 22392
rect 31168 22380 31174 22432
rect 32030 22380 32036 22432
rect 32088 22420 32094 22432
rect 32125 22423 32183 22429
rect 32125 22420 32137 22423
rect 32088 22392 32137 22420
rect 32088 22380 32094 22392
rect 32125 22389 32137 22392
rect 32171 22389 32183 22423
rect 32950 22420 32956 22432
rect 32911 22392 32956 22420
rect 32125 22383 32183 22389
rect 32950 22380 32956 22392
rect 33008 22380 33014 22432
rect 38654 22420 38660 22432
rect 38615 22392 38660 22420
rect 38654 22380 38660 22392
rect 38712 22380 38718 22432
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 2225 22219 2283 22225
rect 2225 22185 2237 22219
rect 2271 22216 2283 22219
rect 2314 22216 2320 22228
rect 2271 22188 2320 22216
rect 2271 22185 2283 22188
rect 2225 22179 2283 22185
rect 2314 22176 2320 22188
rect 2372 22176 2378 22228
rect 6730 22216 6736 22228
rect 5000 22188 6736 22216
rect 3786 22108 3792 22160
rect 3844 22148 3850 22160
rect 5000 22148 5028 22188
rect 6730 22176 6736 22188
rect 6788 22176 6794 22228
rect 11164 22188 12434 22216
rect 9490 22148 9496 22160
rect 3844 22120 5028 22148
rect 9451 22120 9496 22148
rect 3844 22108 3850 22120
rect 4614 22080 4620 22092
rect 1596 22052 4620 22080
rect 1596 22021 1624 22052
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 5000 22089 5028 22120
rect 9490 22108 9496 22120
rect 9548 22108 9554 22160
rect 10962 22108 10968 22160
rect 11020 22148 11026 22160
rect 11164 22148 11192 22188
rect 11020 22120 11192 22148
rect 11020 22108 11026 22120
rect 4985 22083 5043 22089
rect 4985 22049 4997 22083
rect 5031 22080 5043 22083
rect 6822 22080 6828 22092
rect 5031 22052 5065 22080
rect 6783 22052 6828 22080
rect 5031 22049 5043 22052
rect 4985 22043 5043 22049
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 9306 22080 9312 22092
rect 7024 22052 9312 22080
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 21981 1639 22015
rect 2130 22012 2136 22024
rect 1581 21975 1639 21981
rect 1780 21984 2136 22012
rect 1780 21956 1808 21984
rect 2130 21972 2136 21984
rect 2188 22012 2194 22024
rect 2593 22015 2651 22021
rect 2593 22012 2605 22015
rect 2188 21984 2605 22012
rect 2188 21972 2194 21984
rect 2593 21981 2605 21984
rect 2639 21981 2651 22015
rect 5626 22012 5632 22024
rect 2593 21975 2651 21981
rect 2746 21984 5632 22012
rect 1762 21944 1768 21956
rect 1723 21916 1768 21944
rect 1762 21904 1768 21916
rect 1820 21904 1826 21956
rect 2409 21947 2467 21953
rect 2409 21913 2421 21947
rect 2455 21944 2467 21947
rect 2746 21944 2774 21984
rect 5626 21972 5632 21984
rect 5684 21972 5690 22024
rect 7024 22021 7052 22052
rect 9306 22040 9312 22052
rect 9364 22040 9370 22092
rect 11164 22089 11192 22120
rect 12066 22108 12072 22160
rect 12124 22108 12130 22160
rect 12250 22148 12256 22160
rect 12211 22120 12256 22148
rect 12250 22108 12256 22120
rect 12308 22108 12314 22160
rect 12406 22148 12434 22188
rect 17586 22176 17592 22228
rect 17644 22216 17650 22228
rect 17773 22219 17831 22225
rect 17773 22216 17785 22219
rect 17644 22188 17785 22216
rect 17644 22176 17650 22188
rect 17773 22185 17785 22188
rect 17819 22185 17831 22219
rect 17773 22179 17831 22185
rect 12526 22148 12532 22160
rect 12406 22120 12532 22148
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 14182 22108 14188 22160
rect 14240 22148 14246 22160
rect 17788 22148 17816 22179
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 19705 22219 19763 22225
rect 19705 22216 19717 22219
rect 19484 22188 19717 22216
rect 19484 22176 19490 22188
rect 19705 22185 19717 22188
rect 19751 22185 19763 22219
rect 19705 22179 19763 22185
rect 20622 22176 20628 22228
rect 20680 22216 20686 22228
rect 23566 22216 23572 22228
rect 20680 22188 23572 22216
rect 20680 22176 20686 22188
rect 23566 22176 23572 22188
rect 23624 22176 23630 22228
rect 27338 22176 27344 22228
rect 27396 22216 27402 22228
rect 27614 22216 27620 22228
rect 27396 22188 27620 22216
rect 27396 22176 27402 22188
rect 27614 22176 27620 22188
rect 27672 22176 27678 22228
rect 20530 22148 20536 22160
rect 14240 22120 16344 22148
rect 17788 22120 20536 22148
rect 14240 22108 14246 22120
rect 11149 22083 11207 22089
rect 11149 22049 11161 22083
rect 11195 22049 11207 22083
rect 12084 22080 12112 22108
rect 14921 22083 14979 22089
rect 14921 22080 14933 22083
rect 11149 22043 11207 22049
rect 11900 22052 14933 22080
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 21981 7067 22015
rect 7009 21975 7067 21981
rect 7653 22015 7711 22021
rect 7653 21981 7665 22015
rect 7699 21981 7711 22015
rect 7653 21975 7711 21981
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 7926 22012 7932 22024
rect 7883 21984 7932 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 2455 21916 2774 21944
rect 2884 21916 3188 21944
rect 2455 21913 2467 21916
rect 2409 21907 2467 21913
rect 1397 21879 1455 21885
rect 1397 21845 1409 21879
rect 1443 21876 1455 21879
rect 1670 21876 1676 21888
rect 1443 21848 1676 21876
rect 1443 21845 1455 21848
rect 1397 21839 1455 21845
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 2774 21836 2780 21888
rect 2832 21876 2838 21888
rect 2884 21876 2912 21916
rect 3050 21876 3056 21888
rect 2832 21848 2912 21876
rect 3011 21848 3056 21876
rect 2832 21836 2838 21848
rect 3050 21836 3056 21848
rect 3108 21836 3114 21888
rect 3160 21876 3188 21916
rect 4614 21904 4620 21956
rect 4672 21944 4678 21956
rect 5230 21947 5288 21953
rect 5230 21944 5242 21947
rect 4672 21916 5242 21944
rect 4672 21904 4678 21916
rect 5230 21913 5242 21916
rect 5276 21913 5288 21947
rect 7190 21944 7196 21956
rect 5230 21907 5288 21913
rect 5368 21916 6684 21944
rect 7151 21916 7196 21944
rect 3326 21876 3332 21888
rect 3160 21848 3332 21876
rect 3326 21836 3332 21848
rect 3384 21876 3390 21888
rect 5368 21876 5396 21916
rect 3384 21848 5396 21876
rect 6365 21879 6423 21885
rect 3384 21836 3390 21848
rect 6365 21845 6377 21879
rect 6411 21876 6423 21879
rect 6546 21876 6552 21888
rect 6411 21848 6552 21876
rect 6411 21845 6423 21848
rect 6365 21839 6423 21845
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 6656 21876 6684 21916
rect 7190 21904 7196 21916
rect 7248 21904 7254 21956
rect 7668 21944 7696 21975
rect 7926 21972 7932 21984
rect 7984 22012 7990 22024
rect 10873 22015 10931 22021
rect 10873 22012 10885 22015
rect 7984 21984 10885 22012
rect 7984 21972 7990 21984
rect 10873 21981 10885 21984
rect 10919 21981 10931 22015
rect 11606 22012 11612 22024
rect 11567 21984 11612 22012
rect 10873 21975 10931 21981
rect 11606 21972 11612 21984
rect 11664 21972 11670 22024
rect 11698 21972 11704 22024
rect 11756 22012 11762 22024
rect 11900 22021 11928 22052
rect 14921 22049 14933 22052
rect 14967 22080 14979 22083
rect 15470 22080 15476 22092
rect 14967 22052 15476 22080
rect 14967 22049 14979 22052
rect 14921 22043 14979 22049
rect 15470 22040 15476 22052
rect 15528 22040 15534 22092
rect 11885 22015 11943 22021
rect 11756 21984 11801 22012
rect 11756 21972 11762 21984
rect 11885 21981 11897 22015
rect 11931 21981 11943 22015
rect 11885 21975 11943 21981
rect 12115 22015 12173 22021
rect 12115 21981 12127 22015
rect 12161 22012 12173 22015
rect 12342 22012 12348 22024
rect 12161 21984 12348 22012
rect 12161 21981 12173 21984
rect 12115 21975 12173 21981
rect 12342 21972 12348 21984
rect 12400 22012 12406 22024
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 12400 21984 13277 22012
rect 12400 21972 12406 21984
rect 13265 21981 13277 21984
rect 13311 22012 13323 22015
rect 13446 22012 13452 22024
rect 13311 21984 13452 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13446 21972 13452 21984
rect 13504 21972 13510 22024
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 21981 13599 22015
rect 14642 22012 14648 22024
rect 14603 21984 14648 22012
rect 13541 21975 13599 21981
rect 8846 21944 8852 21956
rect 7668 21916 8852 21944
rect 8846 21904 8852 21916
rect 8904 21904 8910 21956
rect 9677 21947 9735 21953
rect 9677 21913 9689 21947
rect 9723 21913 9735 21947
rect 9677 21907 9735 21913
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 6656 21848 7665 21876
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 9692 21876 9720 21907
rect 11974 21904 11980 21956
rect 12032 21944 12038 21956
rect 13556 21944 13584 21975
rect 14642 21972 14648 21984
rect 14700 21972 14706 22024
rect 15930 22012 15936 22024
rect 15891 21984 15936 22012
rect 15930 21972 15936 21984
rect 15988 21972 15994 22024
rect 16022 21972 16028 22024
rect 16080 22012 16086 22024
rect 16316 22021 16344 22120
rect 20530 22108 20536 22120
rect 20588 22148 20594 22160
rect 20990 22148 20996 22160
rect 20588 22120 20996 22148
rect 20588 22108 20594 22120
rect 20990 22108 20996 22120
rect 21048 22108 21054 22160
rect 23382 22148 23388 22160
rect 22388 22120 23388 22148
rect 20714 22080 20720 22092
rect 20272 22052 20720 22080
rect 20272 22021 20300 22052
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 22002 22080 22008 22092
rect 21836 22052 22008 22080
rect 21836 22024 21864 22052
rect 22002 22040 22008 22052
rect 22060 22080 22066 22092
rect 22186 22080 22192 22092
rect 22060 22052 22192 22080
rect 22060 22040 22066 22052
rect 22186 22040 22192 22052
rect 22244 22040 22250 22092
rect 16298 22015 16356 22021
rect 16080 21984 16125 22012
rect 16080 21972 16086 21984
rect 16298 21981 16310 22015
rect 16344 21981 16356 22015
rect 16298 21975 16356 21981
rect 16417 22015 16475 22021
rect 16417 21981 16429 22015
rect 16463 22012 16475 22015
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 16463 21981 16482 22012
rect 16417 21975 16482 21981
rect 14366 21944 14372 21956
rect 12032 21916 12077 21944
rect 13372 21916 14372 21944
rect 12032 21904 12038 21916
rect 13372 21876 13400 21916
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 14660 21944 14688 21972
rect 15010 21944 15016 21956
rect 14660 21916 15016 21944
rect 15010 21904 15016 21916
rect 15068 21904 15074 21956
rect 15470 21904 15476 21956
rect 15528 21944 15534 21956
rect 16209 21947 16267 21953
rect 16209 21944 16221 21947
rect 15528 21916 16221 21944
rect 15528 21904 15534 21916
rect 16209 21913 16221 21916
rect 16255 21913 16267 21947
rect 16209 21907 16267 21913
rect 9692 21848 13400 21876
rect 7653 21839 7711 21845
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 15746 21876 15752 21888
rect 13504 21848 15752 21876
rect 13504 21836 13510 21848
rect 15746 21836 15752 21848
rect 15804 21876 15810 21888
rect 16454 21876 16482 21975
rect 19306 21984 19625 22012
rect 18782 21944 18788 21956
rect 16592 21916 18788 21944
rect 16592 21885 16620 21916
rect 18782 21904 18788 21916
rect 18840 21904 18846 21956
rect 15804 21848 16482 21876
rect 16577 21879 16635 21885
rect 15804 21836 15810 21848
rect 16577 21845 16589 21879
rect 16623 21845 16635 21879
rect 16577 21839 16635 21845
rect 18506 21836 18512 21888
rect 18564 21876 18570 21888
rect 18601 21879 18659 21885
rect 18601 21876 18613 21879
rect 18564 21848 18613 21876
rect 18564 21836 18570 21848
rect 18601 21845 18613 21848
rect 18647 21876 18659 21879
rect 19306 21876 19334 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 20257 22015 20315 22021
rect 20257 21981 20269 22015
rect 20303 21981 20315 22015
rect 20625 22015 20683 22021
rect 20625 22012 20637 22015
rect 20257 21975 20315 21981
rect 20364 21984 20637 22012
rect 19426 21904 19432 21956
rect 19484 21944 19490 21956
rect 20364 21944 20392 21984
rect 20625 21981 20637 21984
rect 20671 21981 20683 22015
rect 20898 22012 20904 22024
rect 20625 21975 20683 21981
rect 20732 21984 20904 22012
rect 19484 21916 20392 21944
rect 20441 21947 20499 21953
rect 19484 21904 19490 21916
rect 20441 21913 20453 21947
rect 20487 21913 20499 21947
rect 20441 21907 20499 21913
rect 18647 21848 19334 21876
rect 20456 21876 20484 21907
rect 20530 21904 20536 21956
rect 20588 21944 20594 21956
rect 20588 21916 20633 21944
rect 20588 21904 20594 21916
rect 20732 21888 20760 21984
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 21818 21972 21824 22024
rect 21876 21972 21882 22024
rect 22094 22012 22100 22024
rect 22055 21984 22100 22012
rect 22094 21972 22100 21984
rect 22152 21972 22158 22024
rect 22278 22012 22284 22024
rect 22239 21984 22284 22012
rect 22278 21972 22284 21984
rect 22336 21972 22342 22024
rect 22388 22021 22416 22120
rect 23382 22108 23388 22120
rect 23440 22108 23446 22160
rect 22741 22083 22799 22089
rect 22741 22049 22753 22083
rect 22787 22049 22799 22083
rect 22741 22043 22799 22049
rect 22373 22015 22431 22021
rect 22373 21981 22385 22015
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 22520 21984 22565 22012
rect 22520 21972 22526 21984
rect 22646 21972 22652 22024
rect 22704 22012 22710 22024
rect 22756 22012 22784 22043
rect 22830 22040 22836 22092
rect 22888 22080 22894 22092
rect 25593 22083 25651 22089
rect 25593 22080 25605 22083
rect 22888 22052 25605 22080
rect 22888 22040 22894 22052
rect 25593 22049 25605 22052
rect 25639 22049 25651 22083
rect 25593 22043 25651 22049
rect 27448 22052 29960 22080
rect 23382 22012 23388 22024
rect 22704 21984 22784 22012
rect 23343 21984 23388 22012
rect 22704 21972 22710 21984
rect 23382 21972 23388 21984
rect 23440 21972 23446 22024
rect 24578 22021 24584 22024
rect 24397 22015 24455 22021
rect 24397 21981 24409 22015
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24545 22015 24584 22021
rect 24545 21981 24557 22015
rect 24545 21975 24584 21981
rect 20824 21916 22094 21944
rect 20714 21876 20720 21888
rect 20456 21848 20720 21876
rect 18647 21845 18659 21848
rect 18601 21839 18659 21845
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 20824 21885 20852 21916
rect 20809 21879 20867 21885
rect 20809 21845 20821 21879
rect 20855 21845 20867 21879
rect 20809 21839 20867 21845
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 21361 21879 21419 21885
rect 21361 21876 21373 21879
rect 21324 21848 21373 21876
rect 21324 21836 21330 21848
rect 21361 21845 21373 21848
rect 21407 21845 21419 21879
rect 22066 21876 22094 21916
rect 22186 21904 22192 21956
rect 22244 21944 22250 21956
rect 22554 21944 22560 21956
rect 22244 21916 22560 21944
rect 22244 21904 22250 21916
rect 22554 21904 22560 21916
rect 22612 21904 22618 21956
rect 24412 21944 24440 21975
rect 24578 21972 24584 21975
rect 24636 21972 24642 22024
rect 24946 22021 24952 22024
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 24903 22015 24952 22021
rect 24903 21981 24915 22015
rect 24949 21981 24952 22015
rect 24903 21975 24952 21981
rect 24670 21944 24676 21956
rect 22664 21916 24440 21944
rect 24631 21916 24676 21944
rect 22664 21876 22692 21916
rect 24670 21904 24676 21916
rect 24728 21904 24734 21956
rect 24780 21944 24808 21975
rect 24946 21972 24952 21975
rect 25004 21972 25010 22024
rect 25682 21972 25688 22024
rect 25740 22012 25746 22024
rect 25849 22015 25907 22021
rect 25849 22012 25861 22015
rect 25740 21984 25861 22012
rect 25740 21972 25746 21984
rect 25849 21981 25861 21984
rect 25895 21981 25907 22015
rect 25849 21975 25907 21981
rect 27448 21944 27476 22052
rect 28166 22012 28172 22024
rect 28127 21984 28172 22012
rect 28166 21972 28172 21984
rect 28224 21972 28230 22024
rect 28258 21972 28264 22024
rect 28316 22012 28322 22024
rect 28353 22015 28411 22021
rect 28353 22012 28365 22015
rect 28316 21984 28365 22012
rect 28316 21972 28322 21984
rect 28353 21981 28365 21984
rect 28399 21981 28411 22015
rect 28353 21975 28411 21981
rect 28442 21972 28448 22024
rect 28500 22012 28506 22024
rect 28583 22015 28641 22021
rect 28500 21984 28545 22012
rect 28500 21972 28506 21984
rect 28583 21981 28595 22015
rect 28629 21981 28641 22015
rect 29932 22012 29960 22052
rect 31386 22040 31392 22092
rect 31444 22080 31450 22092
rect 31444 22052 31892 22080
rect 31444 22040 31450 22052
rect 30098 22012 30104 22024
rect 29932 21984 30104 22012
rect 28583 21975 28641 21981
rect 24780 21916 27476 21944
rect 27614 21904 27620 21956
rect 27672 21944 27678 21956
rect 28598 21944 28626 21975
rect 30098 21972 30104 21984
rect 30156 21972 30162 22024
rect 30929 22015 30987 22021
rect 30929 21981 30941 22015
rect 30975 22012 30987 22015
rect 31754 22012 31760 22024
rect 30975 21984 31760 22012
rect 30975 21981 30987 21984
rect 30929 21975 30987 21981
rect 31754 21972 31760 21984
rect 31812 21972 31818 22024
rect 31864 22021 31892 22052
rect 32398 22040 32404 22092
rect 32456 22080 32462 22092
rect 33060 22080 33364 22094
rect 34057 22083 34115 22089
rect 34057 22080 34069 22083
rect 32456 22066 34069 22080
rect 32456 22052 33088 22066
rect 33336 22052 34069 22066
rect 32456 22040 32462 22052
rect 31849 22015 31907 22021
rect 31849 21981 31861 22015
rect 31895 21981 31907 22015
rect 32030 22012 32036 22024
rect 31991 21984 32036 22012
rect 31849 21975 31907 21981
rect 32030 21972 32036 21984
rect 32088 21972 32094 22024
rect 32125 22015 32183 22021
rect 32125 21981 32137 22015
rect 32171 21981 32183 22015
rect 32125 21975 32183 21981
rect 27672 21916 28626 21944
rect 28813 21947 28871 21953
rect 27672 21904 27678 21916
rect 28813 21913 28825 21947
rect 28859 21944 28871 21947
rect 30662 21947 30720 21953
rect 30662 21944 30674 21947
rect 28859 21916 30674 21944
rect 28859 21913 28871 21916
rect 28813 21907 28871 21913
rect 30662 21913 30674 21916
rect 30708 21913 30720 21947
rect 30662 21907 30720 21913
rect 31202 21904 31208 21956
rect 31260 21944 31266 21956
rect 32140 21944 32168 21975
rect 32214 21972 32220 22024
rect 32272 22012 32278 22024
rect 32968 22021 32996 22052
rect 34057 22049 34069 22052
rect 34103 22049 34115 22083
rect 34057 22043 34115 22049
rect 32953 22015 33011 22021
rect 32272 21984 32317 22012
rect 32272 21972 32278 21984
rect 32953 21981 32965 22015
rect 32999 22012 33011 22015
rect 33134 22012 33140 22024
rect 32999 21984 33033 22012
rect 33095 21984 33140 22012
rect 32999 21981 33011 21984
rect 32953 21975 33011 21981
rect 33134 21972 33140 21984
rect 33192 21972 33198 22024
rect 33229 22015 33287 22021
rect 33229 21981 33241 22015
rect 33275 21981 33287 22015
rect 33229 21975 33287 21981
rect 33244 21944 33272 21975
rect 33318 21972 33324 22024
rect 33376 22012 33382 22024
rect 34330 22012 34336 22024
rect 33376 21984 34336 22012
rect 33376 21972 33382 21984
rect 34330 21972 34336 21984
rect 34388 21972 34394 22024
rect 34514 21972 34520 22024
rect 34572 22012 34578 22024
rect 36265 22015 36323 22021
rect 36265 22012 36277 22015
rect 34572 21984 36277 22012
rect 34572 21972 34578 21984
rect 36265 21981 36277 21984
rect 36311 22012 36323 22015
rect 37458 22012 37464 22024
rect 36311 21984 37464 22012
rect 36311 21981 36323 21984
rect 36265 21975 36323 21981
rect 37458 21972 37464 21984
rect 37516 21972 37522 22024
rect 31260 21916 33272 21944
rect 33597 21947 33655 21953
rect 31260 21904 31266 21916
rect 33597 21913 33609 21947
rect 33643 21944 33655 21947
rect 35998 21947 36056 21953
rect 35998 21944 36010 21947
rect 33643 21916 36010 21944
rect 33643 21913 33655 21916
rect 33597 21907 33655 21913
rect 35998 21913 36010 21916
rect 36044 21913 36056 21947
rect 35998 21907 36056 21913
rect 22066 21848 22692 21876
rect 23293 21879 23351 21885
rect 21361 21839 21419 21845
rect 23293 21845 23305 21879
rect 23339 21876 23351 21879
rect 23382 21876 23388 21888
rect 23339 21848 23388 21876
rect 23339 21845 23351 21848
rect 23293 21839 23351 21845
rect 23382 21836 23388 21848
rect 23440 21836 23446 21888
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 25222 21876 25228 21888
rect 25087 21848 25228 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 25222 21836 25228 21848
rect 25280 21836 25286 21888
rect 26970 21876 26976 21888
rect 26931 21848 26976 21876
rect 26970 21836 26976 21848
rect 27028 21836 27034 21888
rect 27430 21836 27436 21888
rect 27488 21876 27494 21888
rect 29549 21879 29607 21885
rect 29549 21876 29561 21879
rect 27488 21848 29561 21876
rect 27488 21836 27494 21848
rect 29549 21845 29561 21848
rect 29595 21845 29607 21879
rect 29549 21839 29607 21845
rect 31386 21836 31392 21888
rect 31444 21876 31450 21888
rect 32398 21876 32404 21888
rect 31444 21848 32404 21876
rect 31444 21836 31450 21848
rect 32398 21836 32404 21848
rect 32456 21836 32462 21888
rect 32493 21879 32551 21885
rect 32493 21845 32505 21879
rect 32539 21876 32551 21879
rect 33962 21876 33968 21888
rect 32539 21848 33968 21876
rect 32539 21845 32551 21848
rect 32493 21839 32551 21845
rect 33962 21836 33968 21848
rect 34020 21836 34026 21888
rect 34882 21876 34888 21888
rect 34843 21848 34888 21876
rect 34882 21836 34888 21848
rect 34940 21836 34946 21888
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 3234 21672 3240 21684
rect 2271 21644 3240 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 4065 21675 4123 21681
rect 4065 21641 4077 21675
rect 4111 21672 4123 21675
rect 4111 21644 6500 21672
rect 4111 21641 4123 21644
rect 4065 21635 4123 21641
rect 1578 21536 1584 21548
rect 1539 21508 1584 21536
rect 1578 21496 1584 21508
rect 1636 21496 1642 21548
rect 1670 21496 1676 21548
rect 1728 21536 1734 21548
rect 1765 21539 1823 21545
rect 1765 21536 1777 21539
rect 1728 21508 1777 21536
rect 1728 21496 1734 21508
rect 1765 21505 1777 21508
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21505 1915 21539
rect 1857 21499 1915 21505
rect 1949 21539 2007 21545
rect 1949 21505 1961 21539
rect 1995 21536 2007 21539
rect 4080 21536 4108 21635
rect 5442 21564 5448 21616
rect 5500 21604 5506 21616
rect 6365 21607 6423 21613
rect 6365 21604 6377 21607
rect 5500 21576 6377 21604
rect 5500 21564 5506 21576
rect 6365 21573 6377 21576
rect 6411 21573 6423 21607
rect 6472 21604 6500 21644
rect 9398 21632 9404 21684
rect 9456 21672 9462 21684
rect 10226 21672 10232 21684
rect 9456 21644 10232 21672
rect 9456 21632 9462 21644
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 10594 21672 10600 21684
rect 10555 21644 10600 21672
rect 10594 21632 10600 21644
rect 10652 21632 10658 21684
rect 13725 21675 13783 21681
rect 13725 21641 13737 21675
rect 13771 21672 13783 21675
rect 15194 21672 15200 21684
rect 13771 21644 15200 21672
rect 13771 21641 13783 21644
rect 13725 21635 13783 21641
rect 15194 21632 15200 21644
rect 15252 21632 15258 21684
rect 16669 21675 16727 21681
rect 16669 21672 16681 21675
rect 15360 21644 16681 21672
rect 9490 21613 9496 21616
rect 9484 21604 9496 21613
rect 6472 21576 9240 21604
rect 9451 21576 9496 21604
rect 6365 21567 6423 21573
rect 6546 21536 6552 21548
rect 1995 21508 4108 21536
rect 6459 21508 6552 21536
rect 1995 21505 2007 21508
rect 1949 21499 2007 21505
rect 1872 21400 1900 21499
rect 6546 21496 6552 21508
rect 6604 21536 6610 21548
rect 7834 21536 7840 21548
rect 6604 21508 7840 21536
rect 6604 21496 6610 21508
rect 7834 21496 7840 21508
rect 7892 21496 7898 21548
rect 9212 21542 9240 21576
rect 9484 21567 9496 21576
rect 9490 21564 9496 21567
rect 9548 21564 9554 21616
rect 9582 21564 9588 21616
rect 9640 21604 9646 21616
rect 9640 21576 12434 21604
rect 9640 21564 9646 21576
rect 9212 21536 9444 21542
rect 11514 21536 11520 21548
rect 9212 21514 11520 21536
rect 9416 21508 11520 21514
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21468 2743 21471
rect 2774 21468 2780 21480
rect 2731 21440 2780 21468
rect 2731 21437 2743 21440
rect 2685 21431 2743 21437
rect 2774 21428 2780 21440
rect 2832 21428 2838 21480
rect 2961 21471 3019 21477
rect 2961 21437 2973 21471
rect 3007 21437 3019 21471
rect 2961 21431 3019 21437
rect 2314 21400 2320 21412
rect 1872 21372 2320 21400
rect 2314 21360 2320 21372
rect 2372 21400 2378 21412
rect 2976 21400 3004 21431
rect 9214 21428 9220 21480
rect 9272 21468 9278 21480
rect 9272 21440 9317 21468
rect 9272 21428 9278 21440
rect 2372 21372 3004 21400
rect 2372 21360 2378 21372
rect 2700 21344 2728 21372
rect 4798 21360 4804 21412
rect 4856 21400 4862 21412
rect 6733 21403 6791 21409
rect 6733 21400 6745 21403
rect 4856 21372 6745 21400
rect 4856 21360 4862 21372
rect 6733 21369 6745 21372
rect 6779 21369 6791 21403
rect 12406 21400 12434 21576
rect 13078 21564 13084 21616
rect 13136 21604 13142 21616
rect 13357 21607 13415 21613
rect 13357 21604 13369 21607
rect 13136 21576 13369 21604
rect 13136 21564 13142 21576
rect 13357 21573 13369 21576
rect 13403 21573 13415 21607
rect 13357 21567 13415 21573
rect 14553 21607 14611 21613
rect 14553 21573 14565 21607
rect 14599 21604 14611 21607
rect 15360 21604 15388 21644
rect 16669 21641 16681 21644
rect 16715 21672 16727 21675
rect 20901 21675 20959 21681
rect 16715 21644 20668 21672
rect 16715 21641 16727 21644
rect 16669 21635 16727 21641
rect 15470 21604 15476 21616
rect 14599 21576 15388 21604
rect 15431 21576 15476 21604
rect 14599 21573 14611 21576
rect 14553 21567 14611 21573
rect 15470 21564 15476 21576
rect 15528 21564 15534 21616
rect 16574 21564 16580 21616
rect 16632 21604 16638 21616
rect 20640 21613 20668 21644
rect 20901 21641 20913 21675
rect 20947 21672 20959 21675
rect 28258 21672 28264 21684
rect 20947 21644 25728 21672
rect 28219 21644 28264 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 19613 21607 19671 21613
rect 19613 21604 19625 21607
rect 16632 21576 19625 21604
rect 16632 21564 16638 21576
rect 19613 21573 19625 21576
rect 19659 21573 19671 21607
rect 19613 21567 19671 21573
rect 19705 21607 19763 21613
rect 19705 21573 19717 21607
rect 19751 21604 19763 21607
rect 20625 21607 20683 21613
rect 19751 21576 20576 21604
rect 19751 21573 19763 21576
rect 19705 21567 19763 21573
rect 20548 21548 20576 21576
rect 20625 21573 20637 21607
rect 20671 21573 20683 21607
rect 20625 21567 20683 21573
rect 22278 21564 22284 21616
rect 22336 21604 22342 21616
rect 23753 21607 23811 21613
rect 23753 21604 23765 21607
rect 22336 21576 23765 21604
rect 22336 21564 22342 21576
rect 23753 21573 23765 21576
rect 23799 21573 23811 21607
rect 23753 21567 23811 21573
rect 24670 21564 24676 21616
rect 24728 21604 24734 21616
rect 24728 21576 25452 21604
rect 24728 21564 24734 21576
rect 25424 21548 25452 21576
rect 13173 21539 13231 21545
rect 13173 21505 13185 21539
rect 13219 21536 13231 21539
rect 13262 21536 13268 21548
rect 13219 21508 13268 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 13464 21412 13492 21499
rect 13538 21496 13544 21548
rect 13596 21536 13602 21548
rect 14369 21539 14427 21545
rect 13596 21508 13641 21536
rect 13596 21496 13602 21508
rect 14369 21505 14381 21539
rect 14415 21505 14427 21539
rect 15194 21536 15200 21548
rect 15155 21508 15200 21536
rect 14369 21499 14427 21505
rect 14384 21468 14412 21499
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 15378 21545 15384 21548
rect 15345 21539 15384 21545
rect 15345 21505 15357 21539
rect 15345 21499 15384 21505
rect 15378 21496 15384 21499
rect 15436 21496 15442 21548
rect 15746 21545 15752 21548
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21505 15623 21539
rect 15565 21499 15623 21505
rect 15703 21539 15752 21545
rect 15703 21505 15715 21539
rect 15749 21505 15752 21539
rect 15703 21499 15752 21505
rect 14458 21468 14464 21480
rect 13648 21440 14464 21468
rect 12406 21372 13400 21400
rect 6733 21363 6791 21369
rect 2682 21292 2688 21344
rect 2740 21292 2746 21344
rect 5813 21335 5871 21341
rect 5813 21301 5825 21335
rect 5859 21332 5871 21335
rect 5902 21332 5908 21344
rect 5859 21304 5908 21332
rect 5859 21301 5871 21304
rect 5813 21295 5871 21301
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 9214 21292 9220 21344
rect 9272 21332 9278 21344
rect 9582 21332 9588 21344
rect 9272 21304 9588 21332
rect 9272 21292 9278 21304
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 12526 21292 12532 21344
rect 12584 21332 12590 21344
rect 13262 21332 13268 21344
rect 12584 21304 13268 21332
rect 12584 21292 12590 21304
rect 13262 21292 13268 21304
rect 13320 21292 13326 21344
rect 13372 21332 13400 21372
rect 13446 21360 13452 21412
rect 13504 21360 13510 21412
rect 13648 21332 13676 21440
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 15580 21468 15608 21499
rect 15746 21496 15752 21499
rect 15804 21496 15810 21548
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 17782 21539 17840 21545
rect 17782 21536 17794 21539
rect 15896 21508 17794 21536
rect 15896 21496 15902 21508
rect 17782 21505 17794 21508
rect 17828 21505 17840 21539
rect 17782 21499 17840 21505
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21536 18843 21539
rect 18874 21536 18880 21548
rect 18831 21508 18880 21536
rect 18831 21505 18843 21508
rect 18785 21499 18843 21505
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19484 21508 19533 21536
rect 19484 21496 19490 21508
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 20070 21536 20076 21548
rect 19935 21508 20076 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 20349 21539 20407 21545
rect 20349 21505 20361 21539
rect 20395 21505 20407 21539
rect 20530 21536 20536 21548
rect 20491 21508 20536 21536
rect 20349 21499 20407 21505
rect 18046 21468 18052 21480
rect 14568 21440 15608 21468
rect 18007 21440 18052 21468
rect 13372 21304 13676 21332
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 14568 21332 14596 21440
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 20364 21468 20392 21499
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 20717 21539 20775 21545
rect 20717 21505 20729 21539
rect 20763 21536 20775 21539
rect 20898 21536 20904 21548
rect 20763 21508 20904 21536
rect 20763 21505 20775 21508
rect 20717 21499 20775 21505
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 22922 21536 22928 21548
rect 22883 21508 22928 21536
rect 22922 21496 22928 21508
rect 22980 21536 22986 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 22980 21508 23397 21536
rect 22980 21496 22986 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21536 23627 21539
rect 23842 21536 23848 21548
rect 23615 21508 23848 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 24946 21496 24952 21548
rect 25004 21536 25010 21548
rect 25179 21539 25237 21545
rect 25179 21536 25191 21539
rect 25004 21508 25191 21536
rect 25004 21496 25010 21508
rect 25179 21505 25191 21508
rect 25225 21505 25237 21539
rect 25179 21499 25237 21505
rect 25317 21539 25375 21545
rect 25317 21505 25329 21539
rect 25363 21505 25375 21539
rect 25317 21499 25375 21505
rect 20364 21440 22600 21468
rect 18601 21403 18659 21409
rect 18601 21369 18613 21403
rect 18647 21400 18659 21403
rect 22462 21400 22468 21412
rect 18647 21372 22468 21400
rect 18647 21369 18659 21372
rect 18601 21363 18659 21369
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 22572 21400 22600 21440
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 25332 21468 25360 21499
rect 25406 21496 25412 21548
rect 25464 21536 25470 21548
rect 25590 21536 25596 21548
rect 25464 21508 25509 21536
rect 25551 21508 25596 21536
rect 25464 21496 25470 21508
rect 25590 21496 25596 21508
rect 25648 21496 25654 21548
rect 25700 21545 25728 21644
rect 28258 21632 28264 21644
rect 28316 21632 28322 21684
rect 30650 21672 30656 21684
rect 30611 21644 30656 21672
rect 30650 21632 30656 21644
rect 30708 21632 30714 21684
rect 32582 21672 32588 21684
rect 30944 21644 32588 21672
rect 27430 21564 27436 21616
rect 27488 21604 27494 21616
rect 28077 21607 28135 21613
rect 28077 21604 28089 21607
rect 27488 21576 28089 21604
rect 27488 21564 27494 21576
rect 28077 21573 28089 21576
rect 28123 21573 28135 21607
rect 28077 21567 28135 21573
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 27893 21539 27951 21545
rect 27893 21505 27905 21539
rect 27939 21536 27951 21539
rect 27982 21536 27988 21548
rect 27939 21508 27988 21536
rect 27939 21505 27951 21508
rect 27893 21499 27951 21505
rect 27982 21496 27988 21508
rect 28040 21496 28046 21548
rect 29270 21496 29276 21548
rect 29328 21536 29334 21548
rect 30944 21545 30972 21644
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 32677 21675 32735 21681
rect 32677 21641 32689 21675
rect 32723 21672 32735 21675
rect 33134 21672 33140 21684
rect 32723 21644 33140 21672
rect 32723 21641 32735 21644
rect 32677 21635 32735 21641
rect 33134 21632 33140 21644
rect 33192 21632 33198 21684
rect 33502 21672 33508 21684
rect 33463 21644 33508 21672
rect 33502 21632 33508 21644
rect 33560 21632 33566 21684
rect 34882 21672 34888 21684
rect 33612 21644 34888 21672
rect 31202 21604 31208 21616
rect 31036 21576 31208 21604
rect 31036 21545 31064 21576
rect 31202 21564 31208 21576
rect 31260 21564 31266 21616
rect 31662 21564 31668 21616
rect 31720 21604 31726 21616
rect 32309 21607 32367 21613
rect 32309 21604 32321 21607
rect 31720 21576 32321 21604
rect 31720 21564 31726 21576
rect 32309 21573 32321 21576
rect 32355 21573 32367 21607
rect 32309 21567 32367 21573
rect 32493 21607 32551 21613
rect 32493 21573 32505 21607
rect 32539 21604 32551 21607
rect 33612 21604 33640 21644
rect 34882 21632 34888 21644
rect 34940 21632 34946 21684
rect 36633 21675 36691 21681
rect 36633 21641 36645 21675
rect 36679 21672 36691 21675
rect 37550 21672 37556 21684
rect 36679 21644 37556 21672
rect 36679 21641 36691 21644
rect 36633 21635 36691 21641
rect 37550 21632 37556 21644
rect 37608 21632 37614 21684
rect 32539 21576 33640 21604
rect 32539 21573 32551 21576
rect 32493 21567 32551 21573
rect 29549 21539 29607 21545
rect 29549 21536 29561 21539
rect 29328 21508 29561 21536
rect 29328 21496 29334 21508
rect 29549 21505 29561 21508
rect 29595 21505 29607 21539
rect 29549 21499 29607 21505
rect 30193 21539 30251 21545
rect 30193 21505 30205 21539
rect 30239 21536 30251 21539
rect 30929 21539 30987 21545
rect 30929 21536 30941 21539
rect 30239 21508 30941 21536
rect 30239 21505 30251 21508
rect 30193 21499 30251 21505
rect 30929 21505 30941 21508
rect 30975 21505 30987 21539
rect 30929 21499 30987 21505
rect 31021 21539 31079 21545
rect 31021 21505 31033 21539
rect 31067 21505 31079 21539
rect 31021 21499 31079 21505
rect 31110 21496 31116 21548
rect 31168 21536 31174 21548
rect 31297 21539 31355 21545
rect 31168 21508 31213 21536
rect 31168 21496 31174 21508
rect 31297 21505 31309 21539
rect 31343 21536 31355 21539
rect 31386 21536 31392 21548
rect 31343 21508 31392 21536
rect 31343 21505 31355 21508
rect 31297 21499 31355 21505
rect 31386 21496 31392 21508
rect 31444 21496 31450 21548
rect 32508 21468 32536 21567
rect 33962 21564 33968 21616
rect 34020 21604 34026 21616
rect 34618 21607 34676 21613
rect 34618 21604 34630 21607
rect 34020 21576 34630 21604
rect 34020 21564 34026 21576
rect 34618 21573 34630 21576
rect 34664 21573 34676 21607
rect 34618 21567 34676 21573
rect 35529 21607 35587 21613
rect 35529 21573 35541 21607
rect 35575 21604 35587 21607
rect 39298 21604 39304 21616
rect 35575 21576 39304 21604
rect 35575 21573 35587 21576
rect 35529 21567 35587 21573
rect 34330 21496 34336 21548
rect 34388 21536 34394 21548
rect 35544 21536 35572 21567
rect 35986 21536 35992 21548
rect 34388 21508 35572 21536
rect 35947 21508 35992 21536
rect 34388 21496 34394 21508
rect 35986 21496 35992 21508
rect 36044 21496 36050 21548
rect 36170 21536 36176 21548
rect 36131 21508 36176 21536
rect 36170 21496 36176 21508
rect 36228 21496 36234 21548
rect 36262 21496 36268 21548
rect 36320 21536 36326 21548
rect 36403 21539 36461 21545
rect 36320 21508 36365 21536
rect 36320 21496 36326 21508
rect 36403 21505 36415 21539
rect 36449 21536 36461 21539
rect 36556 21536 36584 21576
rect 39298 21564 39304 21576
rect 39356 21564 39362 21616
rect 37458 21536 37464 21548
rect 36449 21508 36584 21536
rect 37419 21508 37464 21536
rect 36449 21505 36461 21508
rect 36403 21499 36461 21505
rect 37458 21496 37464 21508
rect 37516 21496 37522 21548
rect 37734 21545 37740 21548
rect 37728 21499 37740 21545
rect 37792 21536 37798 21548
rect 37792 21508 37828 21536
rect 37734 21496 37740 21499
rect 37792 21496 37798 21508
rect 22704 21440 22749 21468
rect 25332 21440 32536 21468
rect 34885 21471 34943 21477
rect 22704 21428 22710 21440
rect 34885 21437 34897 21471
rect 34931 21437 34943 21471
rect 34885 21431 34943 21437
rect 23106 21400 23112 21412
rect 22572 21372 23112 21400
rect 23106 21360 23112 21372
rect 23164 21360 23170 21412
rect 25498 21360 25504 21412
rect 25556 21400 25562 21412
rect 32950 21400 32956 21412
rect 25556 21372 29684 21400
rect 25556 21360 25562 21372
rect 13780 21304 14596 21332
rect 14737 21335 14795 21341
rect 13780 21292 13786 21304
rect 14737 21301 14749 21335
rect 14783 21332 14795 21335
rect 15378 21332 15384 21344
rect 14783 21304 15384 21332
rect 14783 21301 14795 21304
rect 14737 21295 14795 21301
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 15841 21335 15899 21341
rect 15841 21301 15853 21335
rect 15887 21332 15899 21335
rect 16574 21332 16580 21344
rect 15887 21304 16580 21332
rect 15887 21301 15899 21304
rect 15841 21295 15899 21301
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 19337 21335 19395 21341
rect 19337 21301 19349 21335
rect 19383 21332 19395 21335
rect 20806 21332 20812 21344
rect 19383 21304 20812 21332
rect 19383 21301 19395 21304
rect 19337 21295 19395 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 25038 21332 25044 21344
rect 24999 21304 25044 21332
rect 25038 21292 25044 21304
rect 25096 21292 25102 21344
rect 29656 21332 29684 21372
rect 31726 21372 32956 21400
rect 31726 21332 31754 21372
rect 32950 21360 32956 21372
rect 33008 21360 33014 21412
rect 29656 21304 31754 21332
rect 34514 21292 34520 21344
rect 34572 21332 34578 21344
rect 34900 21332 34928 21431
rect 38838 21332 38844 21344
rect 34572 21304 34928 21332
rect 38799 21304 38844 21332
rect 34572 21292 34578 21304
rect 38838 21292 38844 21304
rect 38896 21292 38902 21344
rect 67634 21332 67640 21344
rect 67595 21304 67640 21332
rect 67634 21292 67640 21304
rect 67692 21292 67698 21344
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 5169 21131 5227 21137
rect 5169 21128 5181 21131
rect 2056 21100 5181 21128
rect 2056 20933 2084 21100
rect 5169 21097 5181 21100
rect 5215 21128 5227 21131
rect 13446 21128 13452 21140
rect 5215 21100 13452 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 14458 21088 14464 21140
rect 14516 21128 14522 21140
rect 15562 21128 15568 21140
rect 14516 21100 15568 21128
rect 14516 21088 14522 21100
rect 15562 21088 15568 21100
rect 15620 21088 15626 21140
rect 15838 21128 15844 21140
rect 15799 21100 15844 21128
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 16206 21088 16212 21140
rect 16264 21128 16270 21140
rect 18506 21128 18512 21140
rect 16264 21100 18512 21128
rect 16264 21088 16270 21100
rect 18506 21088 18512 21100
rect 18564 21088 18570 21140
rect 19426 21088 19432 21140
rect 19484 21128 19490 21140
rect 20898 21128 20904 21140
rect 19484 21100 20904 21128
rect 19484 21088 19490 21100
rect 20898 21088 20904 21100
rect 20956 21088 20962 21140
rect 22462 21088 22468 21140
rect 22520 21128 22526 21140
rect 22741 21131 22799 21137
rect 22741 21128 22753 21131
rect 22520 21100 22753 21128
rect 22520 21088 22526 21100
rect 22741 21097 22753 21100
rect 22787 21097 22799 21131
rect 34054 21128 34060 21140
rect 34015 21100 34060 21128
rect 22741 21091 22799 21097
rect 34054 21088 34060 21100
rect 34112 21088 34118 21140
rect 35437 21131 35495 21137
rect 35437 21097 35449 21131
rect 35483 21128 35495 21131
rect 36170 21128 36176 21140
rect 35483 21100 36176 21128
rect 35483 21097 35495 21100
rect 35437 21091 35495 21097
rect 36170 21088 36176 21100
rect 36228 21088 36234 21140
rect 37734 21088 37740 21140
rect 37792 21128 37798 21140
rect 37829 21131 37887 21137
rect 37829 21128 37841 21131
rect 37792 21100 37841 21128
rect 37792 21088 37798 21100
rect 37829 21097 37841 21100
rect 37875 21097 37887 21131
rect 37829 21091 37887 21097
rect 8113 21063 8171 21069
rect 8113 21029 8125 21063
rect 8159 21029 8171 21063
rect 14182 21060 14188 21072
rect 8113 21023 8171 21029
rect 10428 21032 14188 21060
rect 6730 20992 6736 21004
rect 6691 20964 6736 20992
rect 6730 20952 6736 20964
rect 6788 20952 6794 21004
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20893 2099 20927
rect 2041 20887 2099 20893
rect 2498 20884 2504 20936
rect 2556 20924 2562 20936
rect 2869 20927 2927 20933
rect 2869 20924 2881 20927
rect 2556 20896 2881 20924
rect 2556 20884 2562 20896
rect 2869 20893 2881 20896
rect 2915 20893 2927 20927
rect 2869 20887 2927 20893
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20924 3847 20927
rect 3878 20924 3884 20936
rect 3835 20896 3884 20924
rect 3835 20893 3847 20896
rect 3789 20887 3847 20893
rect 3878 20884 3884 20896
rect 3936 20884 3942 20936
rect 8128 20924 8156 21023
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 8128 20896 9137 20924
rect 9125 20893 9137 20896
rect 9171 20893 9183 20927
rect 9306 20924 9312 20936
rect 9267 20896 9312 20924
rect 9125 20887 9183 20893
rect 1762 20816 1768 20868
rect 1820 20856 1826 20868
rect 1857 20859 1915 20865
rect 1857 20856 1869 20859
rect 1820 20828 1869 20856
rect 1820 20816 1826 20828
rect 1857 20825 1869 20828
rect 1903 20856 1915 20859
rect 1903 20828 2728 20856
rect 1903 20825 1915 20828
rect 1857 20819 1915 20825
rect 2222 20788 2228 20800
rect 2183 20760 2228 20788
rect 2222 20748 2228 20760
rect 2280 20748 2286 20800
rect 2700 20797 2728 20828
rect 3418 20816 3424 20868
rect 3476 20856 3482 20868
rect 4034 20859 4092 20865
rect 4034 20856 4046 20859
rect 3476 20828 4046 20856
rect 3476 20816 3482 20828
rect 4034 20825 4046 20828
rect 4080 20825 4092 20859
rect 4034 20819 4092 20825
rect 7000 20859 7058 20865
rect 7000 20825 7012 20859
rect 7046 20856 7058 20859
rect 7742 20856 7748 20868
rect 7046 20828 7748 20856
rect 7046 20825 7058 20828
rect 7000 20819 7058 20825
rect 7742 20816 7748 20828
rect 7800 20816 7806 20868
rect 7834 20816 7840 20868
rect 7892 20856 7898 20868
rect 9140 20856 9168 20887
rect 9306 20884 9312 20896
rect 9364 20884 9370 20936
rect 10226 20924 10232 20936
rect 10187 20896 10232 20924
rect 10226 20884 10232 20896
rect 10284 20884 10290 20936
rect 9674 20856 9680 20868
rect 7892 20828 9076 20856
rect 9140 20828 9680 20856
rect 7892 20816 7898 20828
rect 2685 20791 2743 20797
rect 2685 20757 2697 20791
rect 2731 20757 2743 20791
rect 2685 20751 2743 20757
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 5718 20788 5724 20800
rect 3108 20760 5724 20788
rect 3108 20748 3114 20760
rect 5718 20748 5724 20760
rect 5776 20748 5782 20800
rect 8202 20748 8208 20800
rect 8260 20788 8266 20800
rect 8941 20791 8999 20797
rect 8941 20788 8953 20791
rect 8260 20760 8953 20788
rect 8260 20748 8266 20760
rect 8941 20757 8953 20760
rect 8987 20757 8999 20791
rect 9048 20788 9076 20828
rect 9674 20816 9680 20828
rect 9732 20816 9738 20868
rect 10428 20865 10456 21032
rect 14182 21020 14188 21032
rect 14240 21020 14246 21072
rect 15286 21020 15292 21072
rect 15344 21060 15350 21072
rect 15344 21032 16344 21060
rect 15344 21020 15350 21032
rect 10686 20952 10692 21004
rect 10744 20992 10750 21004
rect 10744 20964 11376 20992
rect 10744 20952 10750 20964
rect 10502 20884 10508 20936
rect 10560 20924 10566 20936
rect 11348 20933 11376 20964
rect 12894 20952 12900 21004
rect 12952 20992 12958 21004
rect 14645 20995 14703 21001
rect 14645 20992 14657 20995
rect 12952 20964 14657 20992
rect 12952 20952 12958 20964
rect 14645 20961 14657 20964
rect 14691 20992 14703 20995
rect 14691 20964 15608 20992
rect 14691 20961 14703 20964
rect 14645 20955 14703 20961
rect 11057 20927 11115 20933
rect 11057 20924 11069 20927
rect 10560 20896 11069 20924
rect 10560 20884 10566 20896
rect 11057 20893 11069 20896
rect 11103 20893 11115 20927
rect 11057 20887 11115 20893
rect 11241 20927 11299 20933
rect 11241 20893 11253 20927
rect 11287 20893 11299 20927
rect 11241 20887 11299 20893
rect 11333 20927 11391 20933
rect 11333 20893 11345 20927
rect 11379 20893 11391 20927
rect 11333 20887 11391 20893
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20924 11483 20927
rect 11514 20924 11520 20936
rect 11471 20896 11520 20924
rect 11471 20893 11483 20896
rect 11425 20887 11483 20893
rect 10413 20859 10471 20865
rect 10413 20825 10425 20859
rect 10459 20825 10471 20859
rect 10413 20819 10471 20825
rect 10597 20859 10655 20865
rect 10597 20825 10609 20859
rect 10643 20856 10655 20859
rect 11256 20856 11284 20887
rect 11514 20884 11520 20896
rect 11572 20924 11578 20936
rect 12158 20924 12164 20936
rect 11572 20896 12164 20924
rect 11572 20884 11578 20896
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 12986 20924 12992 20936
rect 12947 20896 12992 20924
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 13265 20927 13323 20933
rect 13265 20924 13277 20927
rect 13096 20896 13277 20924
rect 13096 20856 13124 20896
rect 13265 20893 13277 20896
rect 13311 20893 13323 20927
rect 13265 20887 13323 20893
rect 13357 20927 13415 20933
rect 13357 20893 13369 20927
rect 13403 20924 13415 20927
rect 13446 20924 13452 20936
rect 13403 20896 13452 20924
rect 13403 20893 13415 20896
rect 13357 20887 13415 20893
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 15194 20924 15200 20936
rect 15155 20896 15200 20924
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15378 20924 15384 20936
rect 15339 20896 15384 20924
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 15580 20933 15608 20964
rect 16316 20933 16344 21032
rect 20530 21020 20536 21072
rect 20588 21060 20594 21072
rect 24765 21063 24823 21069
rect 24765 21060 24777 21063
rect 20588 21032 24777 21060
rect 20588 21020 20594 21032
rect 24765 21029 24777 21032
rect 24811 21060 24823 21063
rect 25130 21060 25136 21072
rect 24811 21032 25136 21060
rect 24811 21029 24823 21032
rect 24765 21023 24823 21029
rect 25130 21020 25136 21032
rect 25188 21020 25194 21072
rect 26326 21060 26332 21072
rect 26287 21032 26332 21060
rect 26326 21020 26332 21032
rect 26384 21020 26390 21072
rect 30650 21020 30656 21072
rect 30708 21060 30714 21072
rect 31202 21060 31208 21072
rect 30708 21032 31208 21060
rect 30708 21020 30714 21032
rect 31202 21020 31208 21032
rect 31260 21060 31266 21072
rect 31260 21032 32904 21060
rect 31260 21020 31266 21032
rect 25148 20992 25176 21020
rect 16408 20964 16620 20992
rect 25148 20964 25636 20992
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20893 15623 20927
rect 15565 20887 15623 20893
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 10643 20828 11284 20856
rect 11348 20828 13124 20856
rect 10643 20825 10655 20828
rect 10597 20819 10655 20825
rect 11348 20788 11376 20828
rect 13170 20816 13176 20868
rect 13228 20856 13234 20868
rect 13228 20828 13273 20856
rect 13228 20816 13234 20828
rect 13814 20816 13820 20868
rect 13872 20856 13878 20868
rect 15488 20856 15516 20887
rect 16408 20856 16436 20964
rect 16592 20933 16620 20964
rect 16485 20927 16543 20933
rect 16485 20893 16497 20927
rect 16531 20893 16543 20927
rect 16485 20887 16543 20893
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 13872 20828 16436 20856
rect 16500 20856 16528 20887
rect 16666 20884 16672 20936
rect 16724 20924 16730 20936
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 16724 20896 17417 20924
rect 16724 20884 16730 20896
rect 17405 20893 17417 20896
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 18141 20927 18199 20933
rect 18141 20893 18153 20927
rect 18187 20924 18199 20927
rect 18230 20924 18236 20936
rect 18187 20896 18236 20924
rect 18187 20893 18199 20896
rect 18141 20887 18199 20893
rect 18230 20884 18236 20896
rect 18288 20924 18294 20936
rect 18874 20924 18880 20936
rect 18288 20896 18880 20924
rect 18288 20884 18294 20896
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20924 19763 20927
rect 20162 20924 20168 20936
rect 19751 20896 20168 20924
rect 19751 20893 19763 20896
rect 19705 20887 19763 20893
rect 16850 20856 16856 20868
rect 16500 20828 16856 20856
rect 13872 20816 13878 20828
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 16945 20859 17003 20865
rect 16945 20825 16957 20859
rect 16991 20856 17003 20859
rect 17954 20856 17960 20868
rect 16991 20828 17960 20856
rect 16991 20825 17003 20828
rect 16945 20819 17003 20825
rect 17954 20816 17960 20828
rect 18012 20816 18018 20868
rect 19720 20856 19748 20887
rect 20162 20884 20168 20896
rect 20220 20884 20226 20936
rect 23658 20884 23664 20936
rect 23716 20924 23722 20936
rect 25225 20927 25283 20933
rect 25225 20924 25237 20927
rect 23716 20896 25237 20924
rect 23716 20884 23722 20896
rect 25225 20893 25237 20896
rect 25271 20893 25283 20927
rect 25406 20924 25412 20936
rect 25367 20896 25412 20924
rect 25225 20887 25283 20893
rect 25406 20884 25412 20896
rect 25464 20884 25470 20936
rect 25608 20933 25636 20964
rect 30282 20952 30288 21004
rect 30340 20992 30346 21004
rect 31386 20992 31392 21004
rect 30340 20964 31392 20992
rect 30340 20952 30346 20964
rect 31386 20952 31392 20964
rect 31444 20992 31450 21004
rect 31444 20964 32628 20992
rect 31444 20952 31450 20964
rect 25501 20927 25559 20933
rect 25501 20893 25513 20927
rect 25547 20893 25559 20927
rect 25501 20887 25559 20893
rect 25593 20927 25651 20933
rect 25593 20893 25605 20927
rect 25639 20893 25651 20927
rect 25593 20887 25651 20893
rect 25700 20896 27568 20924
rect 18616 20828 19748 20856
rect 11698 20788 11704 20800
rect 9048 20760 11376 20788
rect 11659 20760 11704 20788
rect 8941 20751 8999 20757
rect 11698 20748 11704 20760
rect 11756 20748 11762 20800
rect 13541 20791 13599 20797
rect 13541 20757 13553 20791
rect 13587 20788 13599 20791
rect 13906 20788 13912 20800
rect 13587 20760 13912 20788
rect 13587 20757 13599 20760
rect 13541 20751 13599 20757
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 18506 20748 18512 20800
rect 18564 20788 18570 20800
rect 18616 20797 18644 20828
rect 19978 20816 19984 20868
rect 20036 20856 20042 20868
rect 20533 20859 20591 20865
rect 20533 20856 20545 20859
rect 20036 20828 20545 20856
rect 20036 20816 20042 20828
rect 20533 20825 20545 20828
rect 20579 20825 20591 20859
rect 20533 20819 20591 20825
rect 20640 20828 22094 20856
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18564 20760 18613 20788
rect 18564 20748 18570 20760
rect 18601 20757 18613 20760
rect 18647 20757 18659 20791
rect 18601 20751 18659 20757
rect 19889 20791 19947 20797
rect 19889 20757 19901 20791
rect 19935 20788 19947 20791
rect 20640 20788 20668 20828
rect 19935 20760 20668 20788
rect 19935 20757 19947 20760
rect 19889 20751 19947 20757
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 21818 20788 21824 20800
rect 20772 20760 21824 20788
rect 20772 20748 20778 20760
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 22066 20788 22094 20828
rect 22186 20816 22192 20868
rect 22244 20856 22250 20868
rect 23382 20856 23388 20868
rect 22244 20828 23388 20856
rect 22244 20816 22250 20828
rect 23382 20816 23388 20828
rect 23440 20856 23446 20868
rect 25516 20856 25544 20887
rect 25700 20856 25728 20896
rect 23440 20828 25728 20856
rect 25869 20859 25927 20865
rect 23440 20816 23446 20828
rect 25869 20825 25881 20859
rect 25915 20856 25927 20859
rect 27442 20859 27500 20865
rect 27442 20856 27454 20859
rect 25915 20828 27454 20856
rect 25915 20825 25927 20828
rect 25869 20819 25927 20825
rect 27442 20825 27454 20828
rect 27488 20825 27500 20859
rect 27540 20856 27568 20896
rect 27614 20884 27620 20936
rect 27672 20924 27678 20936
rect 27709 20927 27767 20933
rect 27709 20924 27721 20927
rect 27672 20896 27721 20924
rect 27672 20884 27678 20896
rect 27709 20893 27721 20896
rect 27755 20893 27767 20927
rect 27709 20887 27767 20893
rect 31110 20884 31116 20936
rect 31168 20924 31174 20936
rect 31662 20924 31668 20936
rect 31168 20896 31668 20924
rect 31168 20884 31174 20896
rect 31662 20884 31668 20896
rect 31720 20924 31726 20936
rect 32600 20933 32628 20964
rect 32876 20933 32904 21032
rect 34072 20992 34100 21088
rect 34422 20992 34428 21004
rect 34072 20964 34428 20992
rect 34422 20952 34428 20964
rect 34480 20992 34486 21004
rect 35897 20995 35955 21001
rect 35897 20992 35909 20995
rect 34480 20964 35909 20992
rect 34480 20952 34486 20964
rect 35897 20961 35909 20964
rect 35943 20961 35955 20995
rect 35897 20955 35955 20961
rect 31757 20927 31815 20933
rect 31757 20924 31769 20927
rect 31720 20896 31769 20924
rect 31720 20884 31726 20896
rect 31757 20893 31769 20896
rect 31803 20893 31815 20927
rect 31757 20887 31815 20893
rect 32585 20927 32643 20933
rect 32585 20893 32597 20927
rect 32631 20893 32643 20927
rect 32585 20887 32643 20893
rect 32769 20927 32827 20933
rect 32769 20893 32781 20927
rect 32815 20893 32827 20927
rect 32769 20887 32827 20893
rect 32861 20927 32919 20933
rect 32861 20893 32873 20927
rect 32907 20893 32919 20927
rect 32861 20887 32919 20893
rect 28442 20856 28448 20868
rect 27540 20828 28448 20856
rect 27442 20819 27500 20825
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 31938 20856 31944 20868
rect 28552 20828 31340 20856
rect 31899 20828 31944 20856
rect 22370 20788 22376 20800
rect 22066 20760 22376 20788
rect 22370 20748 22376 20760
rect 22428 20788 22434 20800
rect 28552 20788 28580 20828
rect 22428 20760 28580 20788
rect 22428 20748 22434 20760
rect 29270 20748 29276 20800
rect 29328 20788 29334 20800
rect 30282 20788 30288 20800
rect 29328 20760 30288 20788
rect 29328 20748 29334 20760
rect 30282 20748 30288 20760
rect 30340 20788 30346 20800
rect 31312 20797 31340 20828
rect 31938 20816 31944 20828
rect 31996 20816 32002 20868
rect 32125 20859 32183 20865
rect 32125 20825 32137 20859
rect 32171 20856 32183 20859
rect 32784 20856 32812 20887
rect 32950 20884 32956 20936
rect 33008 20924 33014 20936
rect 33008 20896 33053 20924
rect 33008 20884 33014 20896
rect 34606 20884 34612 20936
rect 34664 20924 34670 20936
rect 35253 20927 35311 20933
rect 35253 20924 35265 20927
rect 34664 20896 35265 20924
rect 34664 20884 34670 20896
rect 35253 20893 35265 20896
rect 35299 20893 35311 20927
rect 35253 20887 35311 20893
rect 32171 20828 32812 20856
rect 35069 20859 35127 20865
rect 32171 20825 32183 20828
rect 32125 20819 32183 20825
rect 35069 20825 35081 20859
rect 35115 20825 35127 20859
rect 35268 20856 35296 20887
rect 35986 20884 35992 20936
rect 36044 20924 36050 20936
rect 36173 20927 36231 20933
rect 36173 20924 36185 20927
rect 36044 20896 36185 20924
rect 36044 20884 36050 20896
rect 36173 20893 36185 20896
rect 36219 20924 36231 20927
rect 37182 20924 37188 20936
rect 36219 20896 37188 20924
rect 36219 20893 36231 20896
rect 36173 20887 36231 20893
rect 37182 20884 37188 20896
rect 37240 20884 37246 20936
rect 37366 20924 37372 20936
rect 37327 20896 37372 20924
rect 37366 20884 37372 20896
rect 37424 20884 37430 20936
rect 37461 20927 37519 20933
rect 37461 20893 37473 20927
rect 37507 20893 37519 20927
rect 37461 20887 37519 20893
rect 35268 20828 36216 20856
rect 35069 20819 35127 20825
rect 30653 20791 30711 20797
rect 30653 20788 30665 20791
rect 30340 20760 30665 20788
rect 30340 20748 30346 20760
rect 30653 20757 30665 20760
rect 30699 20757 30711 20791
rect 30653 20751 30711 20757
rect 31297 20791 31355 20797
rect 31297 20757 31309 20791
rect 31343 20788 31355 20791
rect 32214 20788 32220 20800
rect 31343 20760 32220 20788
rect 31343 20757 31355 20760
rect 31297 20751 31355 20757
rect 32214 20748 32220 20760
rect 32272 20748 32278 20800
rect 33226 20788 33232 20800
rect 33187 20760 33232 20788
rect 33226 20748 33232 20760
rect 33284 20748 33290 20800
rect 35084 20788 35112 20819
rect 36078 20788 36084 20800
rect 35084 20760 36084 20788
rect 36078 20748 36084 20760
rect 36136 20748 36142 20800
rect 36188 20788 36216 20828
rect 36262 20816 36268 20868
rect 36320 20856 36326 20868
rect 37476 20856 37504 20887
rect 37550 20884 37556 20936
rect 37608 20924 37614 20936
rect 37608 20896 37653 20924
rect 37608 20884 37614 20896
rect 37642 20856 37648 20868
rect 36320 20828 37648 20856
rect 36320 20816 36326 20828
rect 37642 20816 37648 20828
rect 37700 20816 37706 20868
rect 38654 20788 38660 20800
rect 36188 20760 38660 20788
rect 38654 20748 38660 20760
rect 38712 20748 38718 20800
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 2685 20587 2743 20593
rect 2685 20553 2697 20587
rect 2731 20584 2743 20587
rect 3418 20584 3424 20596
rect 2731 20556 3424 20584
rect 2731 20553 2743 20556
rect 2685 20547 2743 20553
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 3789 20587 3847 20593
rect 3789 20553 3801 20587
rect 3835 20584 3847 20587
rect 4614 20584 4620 20596
rect 3835 20556 4620 20584
rect 3835 20553 3847 20556
rect 3789 20547 3847 20553
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 7742 20584 7748 20596
rect 7703 20556 7748 20584
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 7926 20544 7932 20596
rect 7984 20584 7990 20596
rect 8938 20584 8944 20596
rect 7984 20556 8944 20584
rect 7984 20544 7990 20556
rect 8938 20544 8944 20556
rect 8996 20584 9002 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 8996 20556 9965 20584
rect 8996 20544 9002 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 14182 20584 14188 20596
rect 14143 20556 14188 20584
rect 9953 20547 10011 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 16850 20544 16856 20596
rect 16908 20584 16914 20596
rect 17037 20587 17095 20593
rect 17037 20584 17049 20587
rect 16908 20556 17049 20584
rect 16908 20544 16914 20556
rect 17037 20553 17049 20556
rect 17083 20553 17095 20587
rect 19978 20584 19984 20596
rect 19939 20556 19984 20584
rect 17037 20547 17095 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 20438 20544 20444 20596
rect 20496 20584 20502 20596
rect 21913 20587 21971 20593
rect 21913 20584 21925 20587
rect 20496 20556 21925 20584
rect 20496 20544 20502 20556
rect 21913 20553 21925 20556
rect 21959 20584 21971 20587
rect 22002 20584 22008 20596
rect 21959 20556 22008 20584
rect 21959 20553 21971 20556
rect 21913 20547 21971 20553
rect 22002 20544 22008 20556
rect 22060 20584 22066 20596
rect 24302 20584 24308 20596
rect 22060 20556 24308 20584
rect 22060 20544 22066 20556
rect 24302 20544 24308 20556
rect 24360 20544 24366 20596
rect 25406 20544 25412 20596
rect 25464 20584 25470 20596
rect 26053 20587 26111 20593
rect 26053 20584 26065 20587
rect 25464 20556 26065 20584
rect 25464 20544 25470 20556
rect 26053 20553 26065 20556
rect 26099 20553 26111 20587
rect 31938 20584 31944 20596
rect 26053 20547 26111 20553
rect 26160 20556 31944 20584
rect 4798 20516 4804 20528
rect 2746 20488 3280 20516
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 2038 20448 2044 20460
rect 1636 20420 2044 20448
rect 1636 20408 1642 20420
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 2222 20448 2228 20460
rect 2183 20420 2228 20448
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 2314 20408 2320 20460
rect 2372 20448 2378 20460
rect 2455 20451 2513 20457
rect 2372 20420 2417 20448
rect 2372 20408 2378 20420
rect 2455 20417 2467 20451
rect 2501 20448 2513 20451
rect 2746 20448 2774 20488
rect 2501 20420 2774 20448
rect 3145 20451 3203 20457
rect 2501 20417 2513 20420
rect 2455 20411 2513 20417
rect 3145 20417 3157 20451
rect 3191 20417 3203 20451
rect 3145 20411 3203 20417
rect 2130 20340 2136 20392
rect 2188 20380 2194 20392
rect 3160 20380 3188 20411
rect 2188 20352 3188 20380
rect 3252 20380 3280 20488
rect 3344 20488 4804 20516
rect 3344 20457 3372 20488
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 7190 20516 7196 20528
rect 7151 20488 7196 20516
rect 7190 20476 7196 20488
rect 7248 20476 7254 20528
rect 9125 20519 9183 20525
rect 9125 20485 9137 20519
rect 9171 20516 9183 20519
rect 9214 20516 9220 20528
rect 9171 20488 9220 20516
rect 9171 20485 9183 20488
rect 9125 20479 9183 20485
rect 9214 20476 9220 20488
rect 9272 20476 9278 20528
rect 9309 20519 9367 20525
rect 9309 20485 9321 20519
rect 9355 20516 9367 20519
rect 9398 20516 9404 20528
rect 9355 20488 9404 20516
rect 9355 20485 9367 20488
rect 9309 20479 9367 20485
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 11698 20476 11704 20528
rect 11756 20516 11762 20528
rect 13050 20519 13108 20525
rect 13050 20516 13062 20519
rect 11756 20488 13062 20516
rect 11756 20476 11762 20488
rect 13050 20485 13062 20488
rect 13096 20485 13108 20519
rect 18046 20516 18052 20528
rect 13050 20479 13108 20485
rect 17696 20488 18052 20516
rect 3329 20451 3387 20457
rect 3329 20417 3341 20451
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 3418 20408 3424 20460
rect 3476 20448 3482 20460
rect 3559 20451 3617 20457
rect 3476 20420 3521 20448
rect 3476 20408 3482 20420
rect 3559 20417 3571 20451
rect 3605 20448 3617 20451
rect 6546 20448 6552 20460
rect 3605 20420 6552 20448
rect 3605 20417 3617 20420
rect 3559 20411 3617 20417
rect 6546 20408 6552 20420
rect 6604 20408 6610 20460
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 3252 20352 4384 20380
rect 2188 20340 2194 20352
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 4356 20253 4384 20352
rect 5810 20272 5816 20324
rect 5868 20312 5874 20324
rect 7024 20312 7052 20411
rect 7926 20408 7932 20460
rect 7984 20457 7990 20460
rect 7984 20451 8033 20457
rect 7984 20417 7987 20451
rect 8021 20417 8033 20451
rect 8110 20448 8116 20460
rect 8071 20420 8116 20448
rect 7984 20411 8033 20417
rect 7984 20408 7990 20411
rect 8110 20408 8116 20420
rect 8168 20408 8174 20460
rect 8202 20408 8208 20460
rect 8260 20448 8266 20460
rect 8389 20451 8447 20457
rect 8260 20420 8305 20448
rect 8260 20408 8266 20420
rect 8389 20417 8401 20451
rect 8435 20417 8447 20451
rect 8389 20411 8447 20417
rect 8404 20380 8432 20411
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 17696 20457 17724 20488
rect 18046 20476 18052 20488
rect 18104 20516 18110 20528
rect 20714 20516 20720 20528
rect 18104 20488 20720 20516
rect 18104 20476 18110 20488
rect 20714 20476 20720 20488
rect 20772 20476 20778 20528
rect 22738 20525 22744 20528
rect 22732 20516 22744 20525
rect 22699 20488 22744 20516
rect 22732 20479 22744 20488
rect 22738 20476 22744 20479
rect 22796 20476 22802 20528
rect 25225 20519 25283 20525
rect 25225 20485 25237 20519
rect 25271 20516 25283 20519
rect 26160 20516 26188 20556
rect 31938 20544 31944 20556
rect 31996 20584 32002 20596
rect 33137 20587 33195 20593
rect 33137 20584 33149 20587
rect 31996 20556 33149 20584
rect 31996 20544 32002 20556
rect 33137 20553 33149 20556
rect 33183 20553 33195 20587
rect 33137 20547 33195 20553
rect 36265 20587 36323 20593
rect 36265 20553 36277 20587
rect 36311 20553 36323 20587
rect 36265 20547 36323 20553
rect 25271 20488 26188 20516
rect 26229 20519 26287 20525
rect 25271 20485 25283 20488
rect 25225 20479 25283 20485
rect 26229 20485 26241 20519
rect 26275 20485 26287 20519
rect 26229 20479 26287 20485
rect 17954 20457 17960 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 15620 20420 16681 20448
rect 15620 20408 15626 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20417 17739 20451
rect 17948 20448 17960 20457
rect 17915 20420 17960 20448
rect 17681 20411 17739 20417
rect 17948 20411 17960 20420
rect 10502 20380 10508 20392
rect 8404 20352 10508 20380
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 11974 20312 11980 20324
rect 5868 20284 11980 20312
rect 5868 20272 5874 20284
rect 11974 20272 11980 20284
rect 12032 20272 12038 20324
rect 4341 20247 4399 20253
rect 4341 20213 4353 20247
rect 4387 20244 4399 20247
rect 5074 20244 5080 20256
rect 4387 20216 5080 20244
rect 4387 20213 4399 20216
rect 4341 20207 4399 20213
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5718 20244 5724 20256
rect 5631 20216 5724 20244
rect 5718 20204 5724 20216
rect 5776 20244 5782 20256
rect 6454 20244 6460 20256
rect 5776 20216 6460 20244
rect 5776 20204 5782 20216
rect 6454 20204 6460 20216
rect 6512 20204 6518 20256
rect 6730 20204 6736 20256
rect 6788 20244 6794 20256
rect 6825 20247 6883 20253
rect 6825 20244 6837 20247
rect 6788 20216 6837 20244
rect 6788 20204 6794 20216
rect 6825 20213 6837 20216
rect 6871 20213 6883 20247
rect 9490 20244 9496 20256
rect 9451 20216 9496 20244
rect 6825 20207 6883 20213
rect 9490 20204 9496 20216
rect 9548 20204 9554 20256
rect 11514 20244 11520 20256
rect 11475 20216 11520 20244
rect 11514 20204 11520 20216
rect 11572 20204 11578 20256
rect 12820 20244 12848 20343
rect 13170 20244 13176 20256
rect 12820 20216 13176 20244
rect 13170 20204 13176 20216
rect 13228 20244 13234 20256
rect 15746 20244 15752 20256
rect 13228 20216 15752 20244
rect 13228 20204 13234 20216
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 16868 20244 16896 20411
rect 17954 20408 17960 20411
rect 18012 20408 18018 20460
rect 20806 20408 20812 20460
rect 20864 20448 20870 20460
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20864 20420 21005 20448
rect 20864 20408 20870 20420
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 21818 20408 21824 20460
rect 21876 20448 21882 20460
rect 22465 20451 22523 20457
rect 22465 20448 22477 20451
rect 21876 20420 22477 20448
rect 21876 20408 21882 20420
rect 22465 20417 22477 20420
rect 22511 20417 22523 20451
rect 22465 20411 22523 20417
rect 24946 20408 24952 20460
rect 25004 20448 25010 20460
rect 25087 20451 25145 20457
rect 25087 20448 25099 20451
rect 25004 20420 25099 20448
rect 25004 20408 25010 20420
rect 25087 20417 25099 20420
rect 25133 20417 25145 20451
rect 25314 20448 25320 20460
rect 25275 20420 25320 20448
rect 25087 20411 25145 20417
rect 25314 20408 25320 20420
rect 25372 20408 25378 20460
rect 25500 20451 25558 20457
rect 25500 20448 25512 20451
rect 25424 20420 25512 20448
rect 21082 20340 21088 20392
rect 21140 20380 21146 20392
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 21140 20352 21281 20380
rect 21140 20340 21146 20352
rect 21269 20349 21281 20352
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 19061 20315 19119 20321
rect 19061 20281 19073 20315
rect 19107 20312 19119 20315
rect 22462 20312 22468 20324
rect 19107 20284 22468 20312
rect 19107 20281 19119 20284
rect 19061 20275 19119 20281
rect 19076 20244 19104 20275
rect 22462 20272 22468 20284
rect 22520 20272 22526 20324
rect 24949 20315 25007 20321
rect 24949 20312 24961 20315
rect 23400 20284 24961 20312
rect 23400 20256 23428 20284
rect 24949 20281 24961 20284
rect 24995 20281 25007 20315
rect 25424 20312 25452 20420
rect 25500 20417 25512 20420
rect 25546 20417 25558 20451
rect 25500 20411 25558 20417
rect 25590 20408 25596 20460
rect 25648 20448 25654 20460
rect 25648 20420 25693 20448
rect 25648 20408 25654 20420
rect 26252 20380 26280 20479
rect 31386 20476 31392 20528
rect 31444 20516 31450 20528
rect 31481 20519 31539 20525
rect 31481 20516 31493 20519
rect 31444 20488 31493 20516
rect 31444 20476 31450 20488
rect 31481 20485 31493 20488
rect 31527 20485 31539 20519
rect 36280 20516 36308 20547
rect 31481 20479 31539 20485
rect 32416 20488 36308 20516
rect 32416 20460 32444 20488
rect 34532 20460 34560 20488
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20448 26479 20451
rect 26510 20448 26516 20460
rect 26467 20420 26516 20448
rect 26467 20417 26479 20420
rect 26421 20411 26479 20417
rect 26510 20408 26516 20420
rect 26568 20448 26574 20460
rect 27982 20448 27988 20460
rect 26568 20420 27988 20448
rect 26568 20408 26574 20420
rect 27982 20408 27988 20420
rect 28040 20408 28046 20460
rect 28169 20451 28227 20457
rect 28169 20417 28181 20451
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 26326 20380 26332 20392
rect 26252 20352 26332 20380
rect 26326 20340 26332 20352
rect 26384 20340 26390 20392
rect 26418 20312 26424 20324
rect 25424 20284 26424 20312
rect 24949 20275 25007 20281
rect 26418 20272 26424 20284
rect 26476 20272 26482 20324
rect 28184 20312 28212 20411
rect 28994 20408 29000 20460
rect 29052 20448 29058 20460
rect 29926 20451 29984 20457
rect 29926 20448 29938 20451
rect 29052 20420 29938 20448
rect 29052 20408 29058 20420
rect 29926 20417 29938 20420
rect 29972 20417 29984 20451
rect 29926 20411 29984 20417
rect 30193 20451 30251 20457
rect 30193 20417 30205 20451
rect 30239 20448 30251 20451
rect 31754 20448 31760 20460
rect 30239 20420 31760 20448
rect 30239 20417 30251 20420
rect 30193 20411 30251 20417
rect 31754 20408 31760 20420
rect 31812 20448 31818 20460
rect 32398 20448 32404 20460
rect 31812 20420 32404 20448
rect 31812 20408 31818 20420
rect 32398 20408 32404 20420
rect 32456 20408 32462 20460
rect 33226 20408 33232 20460
rect 33284 20448 33290 20460
rect 34250 20451 34308 20457
rect 34250 20448 34262 20451
rect 33284 20420 34262 20448
rect 33284 20408 33290 20420
rect 34250 20417 34262 20420
rect 34296 20417 34308 20451
rect 34514 20448 34520 20460
rect 34427 20420 34520 20448
rect 34250 20411 34308 20417
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 34698 20408 34704 20460
rect 34756 20448 34762 20460
rect 34977 20451 35035 20457
rect 34977 20448 34989 20451
rect 34756 20420 34989 20448
rect 34756 20408 34762 20420
rect 34977 20417 34989 20420
rect 35023 20417 35035 20451
rect 34977 20411 35035 20417
rect 28813 20315 28871 20321
rect 28813 20312 28825 20315
rect 28184 20284 28825 20312
rect 16868 20216 19104 20244
rect 23382 20204 23388 20256
rect 23440 20204 23446 20256
rect 23842 20244 23848 20256
rect 23803 20216 23848 20244
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 26050 20204 26056 20256
rect 26108 20244 26114 20256
rect 28184 20244 28212 20284
rect 28813 20281 28825 20284
rect 28859 20281 28871 20315
rect 28813 20275 28871 20281
rect 26108 20216 28212 20244
rect 28353 20247 28411 20253
rect 26108 20204 26114 20216
rect 28353 20213 28365 20247
rect 28399 20244 28411 20247
rect 28534 20244 28540 20256
rect 28399 20216 28540 20244
rect 28399 20213 28411 20216
rect 28353 20207 28411 20213
rect 28534 20204 28540 20216
rect 28592 20204 28598 20256
rect 31938 20204 31944 20256
rect 31996 20244 32002 20256
rect 32493 20247 32551 20253
rect 32493 20244 32505 20247
rect 31996 20216 32505 20244
rect 31996 20204 32002 20216
rect 32493 20213 32505 20216
rect 32539 20244 32551 20247
rect 32950 20244 32956 20256
rect 32539 20216 32956 20244
rect 32539 20213 32551 20216
rect 32493 20207 32551 20213
rect 32950 20204 32956 20216
rect 33008 20244 33014 20256
rect 37369 20247 37427 20253
rect 37369 20244 37381 20247
rect 33008 20216 37381 20244
rect 33008 20204 33014 20216
rect 37369 20213 37381 20216
rect 37415 20244 37427 20247
rect 37550 20244 37556 20256
rect 37415 20216 37556 20244
rect 37415 20213 37427 20216
rect 37369 20207 37427 20213
rect 37550 20204 37556 20216
rect 37608 20244 37614 20256
rect 40402 20244 40408 20256
rect 37608 20216 40408 20244
rect 37608 20204 37614 20216
rect 40402 20204 40408 20216
rect 40460 20204 40466 20256
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 9033 20043 9091 20049
rect 9033 20009 9045 20043
rect 9079 20040 9091 20043
rect 9398 20040 9404 20052
rect 9079 20012 9404 20040
rect 9079 20009 9091 20012
rect 9033 20003 9091 20009
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 9582 20000 9588 20052
rect 9640 20040 9646 20052
rect 9640 20012 11652 20040
rect 9640 20000 9646 20012
rect 2314 19932 2320 19984
rect 2372 19932 2378 19984
rect 7098 19972 7104 19984
rect 6564 19944 7104 19972
rect 2332 19904 2360 19932
rect 2332 19876 2636 19904
rect 1578 19836 1584 19848
rect 1491 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 2038 19796 2044 19848
rect 2096 19836 2102 19848
rect 2317 19839 2375 19845
rect 2317 19836 2329 19839
rect 2096 19808 2329 19836
rect 2096 19796 2102 19808
rect 2317 19805 2329 19808
rect 2363 19805 2375 19839
rect 2498 19836 2504 19848
rect 2459 19808 2504 19836
rect 2317 19799 2375 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 2608 19845 2636 19876
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19805 2651 19839
rect 2593 19799 2651 19805
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 2731 19808 3801 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 4939 19808 5365 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 5353 19805 5365 19808
rect 5399 19836 5411 19839
rect 5442 19836 5448 19848
rect 5399 19808 5448 19836
rect 5399 19805 5411 19808
rect 5353 19799 5411 19805
rect 1596 19768 1624 19796
rect 2406 19768 2412 19780
rect 1596 19740 2412 19768
rect 2406 19728 2412 19740
rect 2464 19728 2470 19780
rect 3804 19768 3832 19799
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 6454 19836 6460 19848
rect 6415 19808 6460 19836
rect 6454 19796 6460 19808
rect 6512 19796 6518 19848
rect 6564 19845 6592 19944
rect 7098 19932 7104 19944
rect 7156 19972 7162 19984
rect 10042 19972 10048 19984
rect 7156 19944 10048 19972
rect 7156 19932 7162 19944
rect 10042 19932 10048 19944
rect 10100 19972 10106 19984
rect 10686 19972 10692 19984
rect 10100 19944 10692 19972
rect 10100 19932 10106 19944
rect 10686 19932 10692 19944
rect 10744 19932 10750 19984
rect 7466 19904 7472 19916
rect 6840 19876 7472 19904
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19836 6699 19839
rect 6730 19836 6736 19848
rect 6687 19808 6736 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 6840 19845 6868 19876
rect 7466 19864 7472 19876
rect 7524 19904 7530 19916
rect 7561 19907 7619 19913
rect 7561 19904 7573 19907
rect 7524 19876 7573 19904
rect 7524 19864 7530 19876
rect 7561 19873 7573 19876
rect 7607 19873 7619 19907
rect 7561 19867 7619 19873
rect 8110 19864 8116 19916
rect 8168 19904 8174 19916
rect 10704 19904 10732 19932
rect 11624 19913 11652 20012
rect 12710 20000 12716 20052
rect 12768 20040 12774 20052
rect 12989 20043 13047 20049
rect 12989 20040 13001 20043
rect 12768 20012 13001 20040
rect 12768 20000 12774 20012
rect 12989 20009 13001 20012
rect 13035 20040 13047 20043
rect 13722 20040 13728 20052
rect 13035 20012 13728 20040
rect 13035 20009 13047 20012
rect 12989 20003 13047 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 21082 20040 21088 20052
rect 18739 20012 21088 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 24949 20043 25007 20049
rect 24176 20012 24716 20040
rect 24176 20000 24182 20012
rect 13814 19932 13820 19984
rect 13872 19972 13878 19984
rect 13872 19944 14964 19972
rect 13872 19932 13878 19944
rect 11609 19907 11667 19913
rect 8168 19876 9444 19904
rect 10704 19876 10824 19904
rect 8168 19864 8174 19876
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 5258 19768 5264 19780
rect 3804 19740 5264 19768
rect 5258 19728 5264 19740
rect 5316 19728 5322 19780
rect 7300 19768 7328 19799
rect 9122 19796 9128 19848
rect 9180 19836 9186 19848
rect 9416 19845 9444 19876
rect 9309 19839 9367 19845
rect 9309 19836 9321 19839
rect 9180 19808 9321 19836
rect 9180 19796 9186 19808
rect 9309 19805 9321 19808
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 7466 19768 7472 19780
rect 7300 19740 7472 19768
rect 7466 19728 7472 19740
rect 7524 19728 7530 19780
rect 1765 19703 1823 19709
rect 1765 19669 1777 19703
rect 1811 19700 1823 19703
rect 2682 19700 2688 19712
rect 1811 19672 2688 19700
rect 1811 19669 1823 19672
rect 1765 19663 1823 19669
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 2958 19700 2964 19712
rect 2919 19672 2964 19700
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 5534 19700 5540 19712
rect 5495 19672 5540 19700
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 6178 19700 6184 19712
rect 6139 19672 6184 19700
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 9416 19700 9444 19799
rect 9490 19796 9496 19848
rect 9548 19836 9554 19848
rect 9677 19839 9735 19845
rect 9548 19808 9593 19836
rect 9548 19796 9554 19808
rect 9677 19805 9689 19839
rect 9723 19805 9735 19839
rect 10502 19836 10508 19848
rect 10463 19808 10508 19836
rect 9677 19799 9735 19805
rect 9692 19768 9720 19799
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 10686 19836 10692 19848
rect 10647 19808 10692 19836
rect 10686 19796 10692 19808
rect 10744 19796 10750 19848
rect 10796 19845 10824 19876
rect 11609 19873 11621 19907
rect 11655 19873 11667 19907
rect 11609 19867 11667 19873
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 10873 19839 10931 19845
rect 10873 19805 10885 19839
rect 10919 19836 10931 19839
rect 10962 19836 10968 19848
rect 10919 19808 10968 19836
rect 10919 19805 10931 19808
rect 10873 19799 10931 19805
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 14645 19839 14703 19845
rect 14645 19836 14657 19839
rect 11072 19808 14657 19836
rect 11072 19768 11100 19808
rect 14645 19805 14657 19808
rect 14691 19836 14703 19839
rect 14734 19836 14740 19848
rect 14691 19808 14740 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 14936 19845 14964 19944
rect 17770 19932 17776 19984
rect 17828 19972 17834 19984
rect 17865 19975 17923 19981
rect 17865 19972 17877 19975
rect 17828 19944 17877 19972
rect 17828 19932 17834 19944
rect 17865 19941 17877 19944
rect 17911 19941 17923 19975
rect 17865 19935 17923 19941
rect 15746 19904 15752 19916
rect 15707 19876 15752 19904
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 20625 19907 20683 19913
rect 20625 19873 20637 19907
rect 20671 19904 20683 19907
rect 20714 19904 20720 19916
rect 20671 19876 20720 19904
rect 20671 19873 20683 19876
rect 20625 19867 20683 19873
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 21376 19904 21404 20000
rect 21928 19944 22094 19972
rect 21821 19907 21879 19913
rect 21821 19904 21833 19907
rect 21376 19876 21833 19904
rect 21821 19873 21833 19876
rect 21867 19873 21879 19907
rect 21821 19867 21879 19873
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19805 14887 19839
rect 14829 19799 14887 19805
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 9692 19740 11100 19768
rect 11149 19771 11207 19777
rect 11149 19737 11161 19771
rect 11195 19768 11207 19771
rect 11854 19771 11912 19777
rect 11854 19768 11866 19771
rect 11195 19740 11866 19768
rect 11195 19737 11207 19740
rect 11149 19731 11207 19737
rect 11854 19737 11866 19740
rect 11900 19737 11912 19771
rect 11854 19731 11912 19737
rect 13722 19728 13728 19780
rect 13780 19768 13786 19780
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 13780 19740 14105 19768
rect 13780 19728 13786 19740
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14844 19768 14872 19799
rect 15010 19796 15016 19848
rect 15068 19836 15074 19848
rect 15764 19836 15792 19864
rect 17310 19836 17316 19848
rect 15068 19808 15113 19836
rect 15764 19808 17316 19836
rect 15068 19796 15074 19808
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 21928 19836 21956 19944
rect 22066 19904 22094 19944
rect 22462 19932 22468 19984
rect 22520 19972 22526 19984
rect 22520 19944 24532 19972
rect 22520 19932 22526 19944
rect 22066 19876 23612 19904
rect 22094 19836 22100 19848
rect 18156 19808 21956 19836
rect 22055 19808 22100 19836
rect 15194 19768 15200 19780
rect 14844 19740 15200 19768
rect 14093 19731 14151 19737
rect 13814 19700 13820 19712
rect 9416 19672 13820 19700
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 14108 19700 14136 19731
rect 15194 19728 15200 19740
rect 15252 19728 15258 19780
rect 15289 19771 15347 19777
rect 15289 19737 15301 19771
rect 15335 19768 15347 19771
rect 15994 19771 16052 19777
rect 15994 19768 16006 19771
rect 15335 19740 16006 19768
rect 15335 19737 15347 19740
rect 15289 19731 15347 19737
rect 15994 19737 16006 19740
rect 16040 19737 16052 19771
rect 15994 19731 16052 19737
rect 16850 19728 16856 19780
rect 16908 19768 16914 19780
rect 18049 19771 18107 19777
rect 18049 19768 18061 19771
rect 16908 19740 18061 19768
rect 16908 19728 16914 19740
rect 18049 19737 18061 19740
rect 18095 19737 18107 19771
rect 18049 19731 18107 19737
rect 15010 19700 15016 19712
rect 14108 19672 15016 19700
rect 15010 19660 15016 19672
rect 15068 19660 15074 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 17129 19703 17187 19709
rect 17129 19700 17141 19703
rect 15528 19672 17141 19700
rect 15528 19660 15534 19672
rect 17129 19669 17141 19672
rect 17175 19700 17187 19703
rect 18156 19700 18184 19808
rect 22094 19796 22100 19808
rect 22152 19796 22158 19848
rect 23290 19836 23296 19848
rect 23251 19808 23296 19836
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23584 19845 23612 19876
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 23661 19839 23719 19845
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 24118 19836 24124 19848
rect 23707 19808 24124 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 24118 19796 24124 19808
rect 24176 19796 24182 19848
rect 24394 19836 24400 19848
rect 24355 19808 24400 19836
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 24504 19836 24532 19944
rect 24688 19904 24716 20012
rect 24949 20009 24961 20043
rect 24995 20040 25007 20043
rect 25590 20040 25596 20052
rect 24995 20012 25596 20040
rect 24995 20009 25007 20012
rect 24949 20003 25007 20009
rect 25590 20000 25596 20012
rect 25648 20000 25654 20052
rect 27798 20040 27804 20052
rect 27759 20012 27804 20040
rect 27798 20000 27804 20012
rect 27856 20000 27862 20052
rect 28994 20040 29000 20052
rect 28955 20012 29000 20040
rect 28994 20000 29000 20012
rect 29052 20000 29058 20052
rect 32214 20000 32220 20052
rect 32272 20040 32278 20052
rect 32272 20012 34661 20040
rect 32272 20000 32278 20012
rect 27816 19972 27844 20000
rect 31113 19975 31171 19981
rect 31113 19972 31125 19975
rect 27816 19944 28764 19972
rect 24688 19876 24808 19904
rect 24780 19845 24808 19876
rect 25682 19864 25688 19916
rect 25740 19904 25746 19916
rect 25740 19876 26188 19904
rect 25740 19864 25746 19876
rect 24673 19839 24731 19845
rect 24673 19836 24685 19839
rect 24504 19808 24685 19836
rect 24673 19805 24685 19808
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19805 24823 19839
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 24765 19799 24823 19805
rect 24872 19808 25881 19836
rect 20380 19771 20438 19777
rect 20380 19737 20392 19771
rect 20426 19768 20438 19771
rect 20622 19768 20628 19780
rect 20426 19740 20628 19768
rect 20426 19737 20438 19740
rect 20380 19731 20438 19737
rect 20622 19728 20628 19740
rect 20680 19728 20686 19780
rect 23477 19771 23535 19777
rect 23477 19737 23489 19771
rect 23523 19768 23535 19771
rect 23934 19768 23940 19780
rect 23523 19740 23940 19768
rect 23523 19737 23535 19740
rect 23477 19731 23535 19737
rect 23934 19728 23940 19740
rect 23992 19768 23998 19780
rect 24581 19771 24639 19777
rect 24581 19768 24593 19771
rect 23992 19740 24593 19768
rect 23992 19728 23998 19740
rect 24581 19737 24593 19740
rect 24627 19737 24639 19771
rect 24581 19731 24639 19737
rect 17175 19672 18184 19700
rect 19245 19703 19303 19709
rect 17175 19669 17187 19672
rect 17129 19663 17187 19669
rect 19245 19669 19257 19703
rect 19291 19700 19303 19703
rect 20254 19700 20260 19712
rect 19291 19672 20260 19700
rect 19291 19669 19303 19672
rect 19245 19663 19303 19669
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20990 19660 20996 19712
rect 21048 19700 21054 19712
rect 22186 19700 22192 19712
rect 21048 19672 22192 19700
rect 21048 19660 21054 19672
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 23845 19703 23903 19709
rect 23845 19669 23857 19703
rect 23891 19700 23903 19703
rect 24872 19700 24900 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 25958 19796 25964 19848
rect 26016 19836 26022 19848
rect 26160 19836 26188 19876
rect 28442 19864 28448 19916
rect 28500 19904 28506 19916
rect 28500 19876 28672 19904
rect 28500 19864 28506 19876
rect 26334 19839 26392 19845
rect 26334 19836 26346 19839
rect 26016 19808 26061 19836
rect 26160 19808 26346 19836
rect 26016 19796 26022 19808
rect 26334 19805 26346 19808
rect 26380 19805 26392 19839
rect 26334 19799 26392 19805
rect 28166 19796 28172 19848
rect 28224 19836 28230 19848
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 28224 19808 28365 19836
rect 28224 19796 28230 19808
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28534 19836 28540 19848
rect 28495 19808 28540 19836
rect 28353 19799 28411 19805
rect 28534 19796 28540 19808
rect 28592 19796 28598 19848
rect 28644 19845 28672 19876
rect 28736 19845 28764 19944
rect 30484 19944 31125 19972
rect 30484 19845 30512 19944
rect 31113 19941 31125 19944
rect 31159 19941 31171 19975
rect 34633 19972 34661 20012
rect 34698 20000 34704 20052
rect 34756 20040 34762 20052
rect 34793 20043 34851 20049
rect 34793 20040 34805 20043
rect 34756 20012 34805 20040
rect 34756 20000 34762 20012
rect 34793 20009 34805 20012
rect 34839 20009 34851 20043
rect 34793 20003 34851 20009
rect 36449 20043 36507 20049
rect 36449 20009 36461 20043
rect 36495 20040 36507 20043
rect 37366 20040 37372 20052
rect 36495 20012 37372 20040
rect 36495 20009 36507 20012
rect 36449 20003 36507 20009
rect 37366 20000 37372 20012
rect 37424 20000 37430 20052
rect 35526 19972 35532 19984
rect 34633 19944 35532 19972
rect 31113 19935 31171 19941
rect 35526 19932 35532 19944
rect 35584 19932 35590 19984
rect 37458 19864 37464 19916
rect 37516 19904 37522 19916
rect 37645 19907 37703 19913
rect 37645 19904 37657 19907
rect 37516 19876 37657 19904
rect 37516 19864 37522 19876
rect 37645 19873 37657 19876
rect 37691 19873 37703 19907
rect 37645 19867 37703 19873
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19805 28687 19839
rect 28629 19799 28687 19805
rect 28721 19839 28779 19845
rect 28721 19805 28733 19839
rect 28767 19805 28779 19839
rect 30469 19839 30527 19845
rect 30469 19836 30481 19839
rect 28721 19799 28779 19805
rect 29288 19808 30481 19836
rect 26142 19768 26148 19780
rect 26103 19740 26148 19768
rect 26142 19728 26148 19740
rect 26200 19728 26206 19780
rect 26237 19771 26295 19777
rect 26237 19737 26249 19771
rect 26283 19768 26295 19771
rect 29288 19768 29316 19808
rect 30469 19805 30481 19808
rect 30515 19805 30527 19839
rect 30469 19799 30527 19805
rect 32398 19796 32404 19848
rect 32456 19836 32462 19848
rect 32493 19839 32551 19845
rect 32493 19836 32505 19839
rect 32456 19808 32505 19836
rect 32456 19796 32462 19808
rect 32493 19805 32505 19808
rect 32539 19805 32551 19839
rect 36078 19836 36084 19848
rect 36039 19808 36084 19836
rect 32493 19799 32551 19805
rect 36078 19796 36084 19808
rect 36136 19836 36142 19848
rect 37090 19836 37096 19848
rect 36136 19808 37096 19836
rect 36136 19796 36142 19808
rect 37090 19796 37096 19808
rect 37148 19796 37154 19848
rect 37366 19796 37372 19848
rect 37424 19836 37430 19848
rect 68094 19836 68100 19848
rect 37424 19808 39068 19836
rect 68055 19808 68100 19836
rect 37424 19796 37430 19808
rect 26283 19740 29316 19768
rect 30285 19771 30343 19777
rect 26283 19737 26295 19740
rect 26237 19731 26295 19737
rect 30285 19737 30297 19771
rect 30331 19768 30343 19771
rect 31110 19768 31116 19780
rect 30331 19740 31116 19768
rect 30331 19737 30343 19740
rect 30285 19731 30343 19737
rect 31110 19728 31116 19740
rect 31168 19728 31174 19780
rect 31202 19728 31208 19780
rect 31260 19768 31266 19780
rect 32226 19771 32284 19777
rect 32226 19768 32238 19771
rect 31260 19740 32238 19768
rect 31260 19728 31266 19740
rect 32226 19737 32238 19740
rect 32272 19737 32284 19771
rect 32226 19731 32284 19737
rect 36170 19728 36176 19780
rect 36228 19768 36234 19780
rect 36265 19771 36323 19777
rect 36265 19768 36277 19771
rect 36228 19740 36277 19768
rect 36228 19728 36234 19740
rect 36265 19737 36277 19740
rect 36311 19737 36323 19771
rect 36265 19731 36323 19737
rect 37912 19771 37970 19777
rect 37912 19737 37924 19771
rect 37958 19768 37970 19771
rect 38102 19768 38108 19780
rect 37958 19740 38108 19768
rect 37958 19737 37970 19740
rect 37912 19731 37970 19737
rect 38102 19728 38108 19740
rect 38160 19728 38166 19780
rect 26510 19700 26516 19712
rect 23891 19672 24900 19700
rect 26471 19672 26516 19700
rect 23891 19669 23903 19672
rect 23845 19663 23903 19669
rect 26510 19660 26516 19672
rect 26568 19660 26574 19712
rect 30653 19703 30711 19709
rect 30653 19669 30665 19703
rect 30699 19700 30711 19703
rect 30742 19700 30748 19712
rect 30699 19672 30748 19700
rect 30699 19669 30711 19672
rect 30653 19663 30711 19669
rect 30742 19660 30748 19672
rect 30800 19660 30806 19712
rect 36538 19660 36544 19712
rect 36596 19700 36602 19712
rect 37182 19700 37188 19712
rect 36596 19672 37188 19700
rect 36596 19660 36602 19672
rect 37182 19660 37188 19672
rect 37240 19700 37246 19712
rect 38838 19700 38844 19712
rect 37240 19672 38844 19700
rect 37240 19660 37246 19672
rect 38838 19660 38844 19672
rect 38896 19660 38902 19712
rect 39040 19709 39068 19808
rect 68094 19796 68100 19808
rect 68152 19796 68158 19848
rect 39025 19703 39083 19709
rect 39025 19669 39037 19703
rect 39071 19669 39083 19703
rect 39025 19663 39083 19669
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 2133 19499 2191 19505
rect 2133 19465 2145 19499
rect 2179 19496 2191 19499
rect 2498 19496 2504 19508
rect 2179 19468 2504 19496
rect 2179 19465 2191 19468
rect 2133 19459 2191 19465
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 2590 19456 2596 19508
rect 2648 19496 2654 19508
rect 5810 19496 5816 19508
rect 2648 19468 2693 19496
rect 5771 19468 5816 19496
rect 2648 19456 2654 19468
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 11054 19496 11060 19508
rect 8404 19468 11060 19496
rect 1762 19428 1768 19440
rect 1723 19400 1768 19428
rect 1762 19388 1768 19400
rect 1820 19388 1826 19440
rect 1949 19431 2007 19437
rect 1949 19397 1961 19431
rect 1995 19428 2007 19431
rect 2608 19428 2636 19456
rect 1995 19400 2636 19428
rect 1995 19397 2007 19400
rect 1949 19391 2007 19397
rect 2958 19388 2964 19440
rect 3016 19428 3022 19440
rect 3706 19431 3764 19437
rect 3706 19428 3718 19431
rect 3016 19400 3718 19428
rect 3016 19388 3022 19400
rect 3706 19397 3718 19400
rect 3752 19397 3764 19431
rect 3706 19391 3764 19397
rect 4700 19431 4758 19437
rect 4700 19397 4712 19431
rect 4746 19428 4758 19431
rect 6178 19428 6184 19440
rect 4746 19400 6184 19428
rect 4746 19397 4758 19400
rect 4700 19391 4758 19397
rect 6178 19388 6184 19400
rect 6236 19388 6242 19440
rect 6638 19388 6644 19440
rect 6696 19428 6702 19440
rect 6733 19431 6791 19437
rect 6733 19428 6745 19431
rect 6696 19400 6745 19428
rect 6696 19388 6702 19400
rect 6733 19397 6745 19400
rect 6779 19397 6791 19431
rect 6733 19391 6791 19397
rect 3878 19320 3884 19372
rect 3936 19360 3942 19372
rect 4433 19363 4491 19369
rect 3936 19332 4016 19360
rect 3936 19320 3942 19332
rect 3988 19301 4016 19332
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 3973 19295 4031 19301
rect 3973 19261 3985 19295
rect 4019 19292 4031 19295
rect 4448 19292 4476 19323
rect 5074 19320 5080 19372
rect 5132 19360 5138 19372
rect 8404 19360 8432 19468
rect 11054 19456 11060 19468
rect 11112 19496 11118 19508
rect 11514 19496 11520 19508
rect 11112 19468 11520 19496
rect 11112 19456 11118 19468
rect 11514 19456 11520 19468
rect 11572 19496 11578 19508
rect 11790 19496 11796 19508
rect 11572 19468 11796 19496
rect 11572 19456 11578 19468
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 12710 19496 12716 19508
rect 12406 19468 12716 19496
rect 9582 19428 9588 19440
rect 8956 19400 9588 19428
rect 8956 19369 8984 19400
rect 9582 19388 9588 19400
rect 9640 19388 9646 19440
rect 10134 19388 10140 19440
rect 10192 19428 10198 19440
rect 11701 19431 11759 19437
rect 10192 19400 11652 19428
rect 10192 19388 10198 19400
rect 5132 19332 8432 19360
rect 8481 19363 8539 19369
rect 5132 19320 5138 19332
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 8941 19363 8999 19369
rect 8941 19360 8953 19363
rect 8527 19332 8953 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 8941 19329 8953 19332
rect 8987 19329 8999 19363
rect 9197 19363 9255 19369
rect 9197 19360 9209 19363
rect 8941 19323 8999 19329
rect 9048 19332 9209 19360
rect 4019 19264 4476 19292
rect 4019 19261 4031 19264
rect 3973 19255 4031 19261
rect 4448 19156 4476 19264
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 9048 19292 9076 19332
rect 9197 19329 9209 19332
rect 9243 19329 9255 19363
rect 9197 19323 9255 19329
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 10468 19332 11529 19360
rect 10468 19320 10474 19332
rect 11517 19329 11529 19332
rect 11563 19329 11575 19363
rect 11624 19360 11652 19400
rect 11701 19397 11713 19431
rect 11747 19428 11759 19431
rect 12406 19428 12434 19468
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 13446 19496 13452 19508
rect 13403 19468 13452 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 14553 19499 14611 19505
rect 14553 19465 14565 19499
rect 14599 19496 14611 19499
rect 15378 19496 15384 19508
rect 14599 19468 15384 19496
rect 14599 19465 14611 19468
rect 14553 19459 14611 19465
rect 15378 19456 15384 19468
rect 15436 19456 15442 19508
rect 15930 19456 15936 19508
rect 15988 19496 15994 19508
rect 18693 19499 18751 19505
rect 18693 19496 18705 19499
rect 15988 19468 18705 19496
rect 15988 19456 15994 19468
rect 18693 19465 18705 19468
rect 18739 19496 18751 19499
rect 24581 19499 24639 19505
rect 18739 19468 24348 19496
rect 18739 19465 18751 19468
rect 18693 19459 18751 19465
rect 14277 19431 14335 19437
rect 14277 19428 14289 19431
rect 11747 19400 12434 19428
rect 12544 19400 14289 19428
rect 11747 19397 11759 19400
rect 11701 19391 11759 19397
rect 12544 19360 12572 19400
rect 14277 19397 14289 19400
rect 14323 19397 14335 19431
rect 14277 19391 14335 19397
rect 14734 19388 14740 19440
rect 14792 19428 14798 19440
rect 15286 19428 15292 19440
rect 14792 19400 15292 19428
rect 14792 19388 14798 19400
rect 15286 19388 15292 19400
rect 15344 19388 15350 19440
rect 15562 19428 15568 19440
rect 15523 19400 15568 19428
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 20165 19431 20223 19437
rect 20165 19397 20177 19431
rect 20211 19428 20223 19431
rect 22925 19431 22983 19437
rect 22925 19428 22937 19431
rect 20211 19400 21956 19428
rect 20211 19397 20223 19400
rect 20165 19391 20223 19397
rect 11624 19332 12572 19360
rect 12621 19363 12679 19369
rect 11517 19323 11575 19329
rect 12621 19329 12633 19363
rect 12667 19360 12679 19363
rect 13446 19360 13452 19372
rect 12667 19332 13452 19360
rect 12667 19329 12679 19332
rect 12621 19323 12679 19329
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 13906 19360 13912 19372
rect 13867 19332 13912 19360
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 14185 19363 14243 19369
rect 14056 19332 14101 19360
rect 14056 19320 14062 19332
rect 14185 19329 14197 19363
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 6972 19264 9076 19292
rect 6972 19252 6978 19264
rect 10686 19252 10692 19304
rect 10744 19292 10750 19304
rect 11885 19295 11943 19301
rect 11885 19292 11897 19295
rect 10744 19264 11897 19292
rect 10744 19252 10750 19264
rect 11885 19261 11897 19264
rect 11931 19261 11943 19295
rect 14200 19292 14228 19323
rect 14366 19320 14372 19372
rect 14424 19369 14430 19372
rect 14424 19360 14432 19369
rect 15381 19363 15439 19369
rect 14424 19332 14469 19360
rect 14424 19323 14432 19332
rect 15381 19329 15393 19363
rect 15427 19360 15439 19363
rect 15470 19360 15476 19372
rect 15427 19332 15476 19360
rect 15427 19329 15439 19332
rect 15381 19323 15439 19329
rect 14424 19320 14430 19323
rect 15470 19320 15476 19332
rect 15528 19320 15534 19372
rect 17310 19360 17316 19372
rect 17271 19332 17316 19360
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 17402 19320 17408 19372
rect 17460 19360 17466 19372
rect 17569 19363 17627 19369
rect 17569 19360 17581 19363
rect 17460 19332 17581 19360
rect 17460 19320 17466 19332
rect 17569 19329 17581 19332
rect 17615 19329 17627 19363
rect 17569 19323 17627 19329
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19360 20039 19363
rect 20254 19360 20260 19372
rect 20027 19332 20260 19360
rect 20027 19329 20039 19332
rect 19981 19323 20039 19329
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20898 19360 20904 19372
rect 20859 19332 20904 19360
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 20990 19363 21048 19369
rect 20990 19346 21002 19363
rect 21036 19346 21048 19363
rect 21085 19363 21143 19369
rect 14642 19292 14648 19304
rect 11885 19255 11943 19261
rect 14016 19264 14648 19292
rect 14016 19236 14044 19264
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 15194 19292 15200 19304
rect 15155 19264 15200 19292
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 16850 19292 16856 19304
rect 16811 19264 16856 19292
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 19797 19295 19855 19301
rect 19797 19261 19809 19295
rect 19843 19292 19855 19295
rect 20990 19294 20996 19346
rect 21048 19294 21054 19346
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21269 19363 21327 19369
rect 21131 19332 21211 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 19843 19264 20944 19292
rect 19843 19261 19855 19264
rect 19797 19255 19855 19261
rect 12802 19224 12808 19236
rect 9876 19196 12434 19224
rect 12763 19196 12808 19224
rect 5350 19156 5356 19168
rect 4448 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 9876 19156 9904 19196
rect 6512 19128 9904 19156
rect 6512 19116 6518 19128
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10321 19159 10379 19165
rect 10321 19156 10333 19159
rect 10192 19128 10333 19156
rect 10192 19116 10198 19128
rect 10321 19125 10333 19128
rect 10367 19125 10379 19159
rect 12406 19156 12434 19196
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 13998 19184 14004 19236
rect 14056 19184 14062 19236
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 16868 19224 16896 19252
rect 20622 19224 20628 19236
rect 14240 19196 16896 19224
rect 20583 19196 20628 19224
rect 14240 19184 14246 19196
rect 20622 19184 20628 19196
rect 20680 19184 20686 19236
rect 14458 19156 14464 19168
rect 12406 19128 14464 19156
rect 10321 19119 10379 19125
rect 14458 19116 14464 19128
rect 14516 19156 14522 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 14516 19128 16037 19156
rect 14516 19116 14522 19128
rect 16025 19125 16037 19128
rect 16071 19156 16083 19159
rect 16666 19156 16672 19168
rect 16071 19128 16672 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 19337 19159 19395 19165
rect 19337 19125 19349 19159
rect 19383 19156 19395 19159
rect 20070 19156 20076 19168
rect 19383 19128 20076 19156
rect 19383 19125 19395 19128
rect 19337 19119 19395 19125
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 20916 19156 20944 19264
rect 21183 19156 21211 19332
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 21315 19332 21772 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 21744 19224 21772 19332
rect 21928 19292 21956 19400
rect 22388 19400 22937 19428
rect 22002 19320 22008 19372
rect 22060 19369 22066 19372
rect 22060 19363 22109 19369
rect 22060 19329 22063 19363
rect 22097 19329 22109 19363
rect 22183 19360 22189 19372
rect 22144 19332 22189 19360
rect 22060 19323 22109 19329
rect 22060 19320 22066 19323
rect 22183 19320 22189 19332
rect 22241 19320 22247 19372
rect 22281 19363 22339 19369
rect 22281 19329 22293 19363
rect 22327 19360 22339 19363
rect 22388 19360 22416 19400
rect 22925 19397 22937 19400
rect 22971 19397 22983 19431
rect 22925 19391 22983 19397
rect 23934 19388 23940 19440
rect 23992 19428 23998 19440
rect 24320 19437 24348 19468
rect 24581 19465 24593 19499
rect 24627 19465 24639 19499
rect 24581 19459 24639 19465
rect 24213 19431 24271 19437
rect 24213 19428 24225 19431
rect 23992 19400 24225 19428
rect 23992 19388 23998 19400
rect 24213 19397 24225 19400
rect 24259 19397 24271 19431
rect 24213 19391 24271 19397
rect 24305 19431 24363 19437
rect 24305 19397 24317 19431
rect 24351 19397 24363 19431
rect 24596 19428 24624 19459
rect 25590 19456 25596 19508
rect 25648 19496 25654 19508
rect 25777 19499 25835 19505
rect 25777 19496 25789 19499
rect 25648 19468 25789 19496
rect 25648 19456 25654 19468
rect 25777 19465 25789 19468
rect 25823 19465 25835 19499
rect 31202 19496 31208 19508
rect 31163 19468 31208 19496
rect 25777 19459 25835 19465
rect 31202 19456 31208 19468
rect 31260 19456 31266 19508
rect 35897 19499 35955 19505
rect 35897 19465 35909 19499
rect 35943 19496 35955 19499
rect 37274 19496 37280 19508
rect 35943 19468 37280 19496
rect 35943 19465 35955 19468
rect 35897 19459 35955 19465
rect 37274 19456 37280 19468
rect 37332 19456 37338 19508
rect 38102 19496 38108 19508
rect 38063 19468 38108 19496
rect 38102 19456 38108 19468
rect 38160 19456 38166 19508
rect 24596 19400 26464 19428
rect 24305 19391 24363 19397
rect 22327 19332 22416 19360
rect 22465 19363 22523 19369
rect 22327 19329 22339 19332
rect 22281 19323 22339 19329
rect 22465 19329 22477 19363
rect 22511 19334 22523 19363
rect 23109 19363 23167 19369
rect 22554 19334 22560 19346
rect 22511 19329 22560 19334
rect 22465 19323 22560 19329
rect 22480 19306 22560 19323
rect 22554 19294 22560 19306
rect 22612 19294 22618 19346
rect 23109 19329 23121 19363
rect 23155 19329 23167 19363
rect 23293 19363 23351 19369
rect 23293 19360 23305 19363
rect 23109 19323 23167 19329
rect 23216 19332 23305 19360
rect 21928 19264 22140 19292
rect 22112 19224 22140 19264
rect 22922 19252 22928 19304
rect 22980 19292 22986 19304
rect 23124 19292 23152 19323
rect 22980 19264 23152 19292
rect 22980 19252 22986 19264
rect 22646 19224 22652 19236
rect 21744 19196 21951 19224
rect 22112 19196 22652 19224
rect 20916 19128 21211 19156
rect 21450 19116 21456 19168
rect 21508 19156 21514 19168
rect 21821 19159 21879 19165
rect 21821 19156 21833 19159
rect 21508 19128 21833 19156
rect 21508 19116 21514 19128
rect 21821 19125 21833 19128
rect 21867 19125 21879 19159
rect 21923 19156 21951 19196
rect 22646 19184 22652 19196
rect 22704 19224 22710 19236
rect 23216 19224 23244 19332
rect 23293 19329 23305 19332
rect 23339 19329 23351 19363
rect 24026 19360 24032 19372
rect 23987 19332 24032 19360
rect 23293 19323 23351 19329
rect 24026 19320 24032 19332
rect 24084 19320 24090 19372
rect 24118 19320 24124 19372
rect 24176 19360 24182 19372
rect 24397 19363 24455 19369
rect 24397 19360 24409 19363
rect 24176 19332 24409 19360
rect 24176 19320 24182 19332
rect 24397 19329 24409 19332
rect 24443 19329 24455 19363
rect 24397 19323 24455 19329
rect 25682 19320 25688 19372
rect 25740 19360 25746 19372
rect 25915 19363 25973 19369
rect 25915 19360 25927 19363
rect 25740 19332 25927 19360
rect 25740 19320 25746 19332
rect 25915 19329 25927 19332
rect 25961 19329 25973 19363
rect 25915 19323 25973 19329
rect 26053 19363 26111 19369
rect 26053 19329 26065 19363
rect 26099 19329 26111 19363
rect 26053 19323 26111 19329
rect 26068 19292 26096 19323
rect 26142 19320 26148 19372
rect 26200 19360 26206 19372
rect 26326 19360 26332 19372
rect 26200 19332 26245 19360
rect 26287 19332 26332 19360
rect 26200 19320 26206 19332
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 26436 19369 26464 19400
rect 30650 19388 30656 19440
rect 30708 19428 30714 19440
rect 30708 19400 30880 19428
rect 30708 19388 30714 19400
rect 26421 19363 26479 19369
rect 26421 19329 26433 19363
rect 26467 19329 26479 19363
rect 26421 19323 26479 19329
rect 26694 19320 26700 19372
rect 26752 19360 26758 19372
rect 28810 19360 28816 19372
rect 26752 19332 28816 19360
rect 26752 19320 26758 19332
rect 28810 19320 28816 19332
rect 28868 19360 28874 19372
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 28868 19332 29745 19360
rect 28868 19320 28874 19332
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29822 19320 29828 19372
rect 29880 19360 29886 19372
rect 29917 19363 29975 19369
rect 29917 19360 29929 19363
rect 29880 19332 29929 19360
rect 29880 19320 29886 19332
rect 29917 19329 29929 19332
rect 29963 19329 29975 19363
rect 29917 19323 29975 19329
rect 30098 19320 30104 19372
rect 30156 19360 30162 19372
rect 30561 19363 30619 19369
rect 30561 19360 30573 19363
rect 30156 19332 30573 19360
rect 30156 19320 30162 19332
rect 30561 19329 30573 19332
rect 30607 19329 30619 19363
rect 30742 19360 30748 19372
rect 30703 19332 30748 19360
rect 30561 19323 30619 19329
rect 30742 19320 30748 19332
rect 30800 19320 30806 19372
rect 30852 19369 30880 19400
rect 34514 19388 34520 19440
rect 34572 19428 34578 19440
rect 34572 19400 35020 19428
rect 34572 19388 34578 19400
rect 30840 19363 30898 19369
rect 30840 19329 30852 19363
rect 30886 19329 30898 19363
rect 30840 19323 30898 19329
rect 30929 19363 30987 19369
rect 30929 19329 30941 19363
rect 30975 19329 30987 19363
rect 30929 19323 30987 19329
rect 34721 19363 34779 19369
rect 34721 19329 34733 19363
rect 34767 19360 34779 19363
rect 34882 19360 34888 19372
rect 34767 19332 34888 19360
rect 34767 19329 34779 19332
rect 34721 19323 34779 19329
rect 26878 19292 26884 19304
rect 26068 19264 26884 19292
rect 26878 19252 26884 19264
rect 26936 19252 26942 19304
rect 30944 19292 30972 19323
rect 34882 19320 34888 19332
rect 34940 19320 34946 19372
rect 34992 19369 35020 19400
rect 35526 19388 35532 19440
rect 35584 19428 35590 19440
rect 37645 19431 37703 19437
rect 35584 19400 36216 19428
rect 35584 19388 35590 19400
rect 36188 19369 36216 19400
rect 37645 19397 37657 19431
rect 37691 19428 37703 19431
rect 37691 19400 38608 19428
rect 37691 19397 37703 19400
rect 37645 19391 37703 19397
rect 34977 19363 35035 19369
rect 34977 19329 34989 19363
rect 35023 19329 35035 19363
rect 34977 19323 35035 19329
rect 36173 19363 36231 19369
rect 36173 19329 36185 19363
rect 36219 19329 36231 19363
rect 36173 19323 36231 19329
rect 36262 19366 36320 19372
rect 36262 19332 36274 19366
rect 36308 19332 36320 19366
rect 36262 19326 36320 19332
rect 36378 19363 36436 19369
rect 36378 19329 36390 19363
rect 36424 19360 36436 19363
rect 36424 19329 36446 19360
rect 30024 19264 31754 19292
rect 22704 19196 23244 19224
rect 22704 19184 22710 19196
rect 22094 19156 22100 19168
rect 21923 19128 22100 19156
rect 21821 19119 21879 19125
rect 22094 19116 22100 19128
rect 22152 19156 22158 19168
rect 22554 19156 22560 19168
rect 22152 19128 22560 19156
rect 22152 19116 22158 19128
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 26602 19156 26608 19168
rect 24912 19128 26608 19156
rect 24912 19116 24918 19128
rect 26602 19116 26608 19128
rect 26660 19156 26666 19168
rect 30024 19156 30052 19264
rect 31726 19224 31754 19264
rect 36280 19236 36308 19326
rect 36378 19323 36446 19329
rect 36418 19236 36446 19323
rect 36538 19320 36544 19372
rect 36596 19360 36602 19372
rect 36596 19332 36641 19360
rect 36596 19320 36602 19332
rect 37090 19320 37096 19372
rect 37148 19360 37154 19372
rect 37277 19363 37335 19369
rect 37277 19360 37289 19363
rect 37148 19332 37289 19360
rect 37148 19320 37154 19332
rect 37277 19329 37289 19332
rect 37323 19329 37335 19363
rect 37277 19323 37335 19329
rect 37366 19320 37372 19372
rect 37424 19360 37430 19372
rect 37461 19363 37519 19369
rect 37461 19360 37473 19363
rect 37424 19332 37473 19360
rect 37424 19320 37430 19332
rect 37461 19329 37473 19332
rect 37507 19329 37519 19363
rect 37461 19323 37519 19329
rect 37550 19320 37556 19372
rect 37608 19360 37614 19372
rect 38335 19363 38393 19369
rect 38335 19360 38347 19363
rect 37608 19332 38347 19360
rect 37608 19320 37614 19332
rect 38335 19329 38347 19332
rect 38381 19329 38393 19363
rect 38470 19360 38476 19372
rect 38431 19332 38476 19360
rect 38335 19323 38393 19329
rect 38470 19320 38476 19332
rect 38528 19320 38534 19372
rect 38580 19369 38608 19400
rect 38565 19363 38623 19369
rect 38565 19329 38577 19363
rect 38611 19329 38623 19363
rect 38565 19323 38623 19329
rect 38749 19363 38807 19369
rect 38749 19329 38761 19363
rect 38795 19360 38807 19363
rect 38838 19360 38844 19372
rect 38795 19332 38844 19360
rect 38795 19329 38807 19332
rect 38749 19323 38807 19329
rect 38838 19320 38844 19332
rect 38896 19320 38902 19372
rect 32217 19227 32275 19233
rect 32217 19224 32229 19227
rect 31726 19196 32229 19224
rect 32217 19193 32229 19196
rect 32263 19224 32275 19227
rect 32263 19196 34100 19224
rect 32263 19193 32275 19196
rect 32217 19187 32275 19193
rect 26660 19128 30052 19156
rect 30101 19159 30159 19165
rect 26660 19116 26666 19128
rect 30101 19125 30113 19159
rect 30147 19156 30159 19159
rect 30282 19156 30288 19168
rect 30147 19128 30288 19156
rect 30147 19125 30159 19128
rect 30101 19119 30159 19125
rect 30282 19116 30288 19128
rect 30340 19116 30346 19168
rect 33597 19159 33655 19165
rect 33597 19125 33609 19159
rect 33643 19156 33655 19159
rect 33962 19156 33968 19168
rect 33643 19128 33968 19156
rect 33643 19125 33655 19128
rect 33597 19119 33655 19125
rect 33962 19116 33968 19128
rect 34020 19116 34026 19168
rect 34072 19156 34100 19196
rect 36262 19184 36268 19236
rect 36320 19184 36326 19236
rect 36418 19196 36452 19236
rect 36446 19184 36452 19196
rect 36504 19184 36510 19236
rect 37550 19156 37556 19168
rect 34072 19128 37556 19156
rect 37550 19116 37556 19128
rect 37608 19116 37614 19168
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 6914 18952 6920 18964
rect 6503 18924 6920 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 8938 18952 8944 18964
rect 8899 18924 8944 18952
rect 8938 18912 8944 18924
rect 8996 18952 9002 18964
rect 11330 18952 11336 18964
rect 8996 18924 11336 18952
rect 8996 18912 9002 18924
rect 11330 18912 11336 18924
rect 11388 18912 11394 18964
rect 17221 18955 17279 18961
rect 17221 18921 17233 18955
rect 17267 18952 17279 18955
rect 17310 18952 17316 18964
rect 17267 18924 17316 18952
rect 17267 18921 17279 18924
rect 17221 18915 17279 18921
rect 17310 18912 17316 18924
rect 17368 18912 17374 18964
rect 18690 18952 18696 18964
rect 18651 18924 18696 18952
rect 18690 18912 18696 18924
rect 18748 18912 18754 18964
rect 20073 18955 20131 18961
rect 20073 18921 20085 18955
rect 20119 18952 20131 18955
rect 20530 18952 20536 18964
rect 20119 18924 20536 18952
rect 20119 18921 20131 18924
rect 20073 18915 20131 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 24854 18952 24860 18964
rect 20916 18924 24860 18952
rect 7558 18884 7564 18896
rect 6840 18856 7564 18884
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2317 18819 2375 18825
rect 2317 18816 2329 18819
rect 2096 18788 2329 18816
rect 2096 18776 2102 18788
rect 2317 18785 2329 18788
rect 2363 18785 2375 18819
rect 2317 18779 2375 18785
rect 2593 18819 2651 18825
rect 2593 18785 2605 18819
rect 2639 18816 2651 18819
rect 3142 18816 3148 18828
rect 2639 18788 3148 18816
rect 2639 18785 2651 18788
rect 2593 18779 2651 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 6840 18757 6868 18856
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 10502 18844 10508 18896
rect 10560 18844 10566 18896
rect 11698 18844 11704 18896
rect 11756 18884 11762 18896
rect 14093 18887 14151 18893
rect 14093 18884 14105 18887
rect 11756 18856 14105 18884
rect 11756 18844 11762 18856
rect 14093 18853 14105 18856
rect 14139 18884 14151 18887
rect 15838 18884 15844 18896
rect 14139 18856 15844 18884
rect 14139 18853 14151 18856
rect 14093 18847 14151 18853
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 19429 18887 19487 18893
rect 19429 18853 19441 18887
rect 19475 18884 19487 18887
rect 20916 18884 20944 18924
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 29822 18952 29828 18964
rect 25056 18924 29828 18952
rect 19475 18856 20944 18884
rect 19475 18853 19487 18856
rect 19429 18847 19487 18853
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7116 18788 7849 18816
rect 6733 18751 6791 18757
rect 6733 18717 6745 18751
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 6546 18640 6552 18692
rect 6604 18680 6610 18692
rect 6748 18680 6776 18711
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7116 18757 7144 18788
rect 7837 18785 7849 18788
rect 7883 18816 7895 18819
rect 10520 18816 10548 18844
rect 11241 18819 11299 18825
rect 11241 18816 11253 18819
rect 7883 18788 10548 18816
rect 10612 18788 11253 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 7101 18751 7159 18757
rect 6972 18720 7017 18748
rect 6972 18708 6978 18720
rect 7101 18717 7113 18751
rect 7147 18717 7159 18751
rect 7558 18748 7564 18760
rect 7519 18720 7564 18748
rect 7101 18711 7159 18717
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 10152 18757 10180 18788
rect 10137 18751 10195 18757
rect 10137 18717 10149 18751
rect 10183 18717 10195 18751
rect 10318 18748 10324 18760
rect 10279 18720 10324 18748
rect 10137 18711 10195 18717
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 10612 18748 10640 18788
rect 11241 18785 11253 18788
rect 11287 18816 11299 18819
rect 13906 18816 13912 18828
rect 11287 18788 13912 18816
rect 11287 18785 11299 18788
rect 11241 18779 11299 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 15562 18816 15568 18828
rect 15243 18788 15568 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 15562 18776 15568 18788
rect 15620 18776 15626 18828
rect 20714 18776 20720 18828
rect 20772 18816 20778 18828
rect 20901 18819 20959 18825
rect 20901 18816 20913 18819
rect 20772 18788 20913 18816
rect 20772 18776 20778 18788
rect 20901 18785 20913 18788
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 10551 18720 10640 18748
rect 12345 18751 12403 18757
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 12345 18717 12357 18751
rect 12391 18748 12403 18751
rect 12434 18748 12440 18760
rect 12391 18720 12440 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 9674 18680 9680 18692
rect 6604 18652 9680 18680
rect 6604 18640 6610 18652
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 10042 18640 10048 18692
rect 10100 18680 10106 18692
rect 10428 18680 10456 18711
rect 10100 18652 10456 18680
rect 10100 18640 10106 18652
rect 3142 18612 3148 18624
rect 3103 18584 3148 18612
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 3786 18572 3792 18624
rect 3844 18612 3850 18624
rect 4890 18612 4896 18624
rect 3844 18584 4896 18612
rect 3844 18572 3850 18584
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 5258 18572 5264 18624
rect 5316 18612 5322 18624
rect 10520 18612 10548 18711
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 12618 18748 12624 18760
rect 12579 18720 12624 18748
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 12713 18751 12771 18757
rect 12713 18717 12725 18751
rect 12759 18748 12771 18751
rect 13354 18748 13360 18760
rect 12759 18720 13360 18748
rect 12759 18717 12771 18720
rect 12713 18711 12771 18717
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 15470 18748 15476 18760
rect 15431 18720 15476 18748
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 18690 18748 18696 18760
rect 18564 18720 18696 18748
rect 18564 18708 18570 18720
rect 18690 18708 18696 18720
rect 18748 18748 18754 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18748 18720 19257 18748
rect 18748 18708 18754 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 20070 18708 20076 18760
rect 20128 18748 20134 18760
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 20128 18720 20269 18748
rect 20128 18708 20134 18720
rect 20257 18717 20269 18720
rect 20303 18717 20315 18751
rect 20257 18711 20315 18717
rect 21168 18751 21226 18757
rect 21168 18717 21180 18751
rect 21214 18748 21226 18751
rect 21450 18748 21456 18760
rect 21214 18720 21456 18748
rect 21214 18717 21226 18720
rect 21168 18711 21226 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 21726 18708 21732 18760
rect 21784 18748 21790 18760
rect 21910 18748 21916 18760
rect 21784 18720 21916 18748
rect 21784 18708 21790 18720
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22554 18708 22560 18760
rect 22612 18748 22618 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22612 18720 23029 18748
rect 22612 18708 22618 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18748 23351 18751
rect 23934 18748 23940 18760
rect 23339 18720 23940 18748
rect 23339 18717 23351 18720
rect 23293 18711 23351 18717
rect 23934 18708 23940 18720
rect 23992 18708 23998 18760
rect 25056 18757 25084 18924
rect 29822 18912 29828 18924
rect 29880 18952 29886 18964
rect 31573 18955 31631 18961
rect 31573 18952 31585 18955
rect 29880 18924 31585 18952
rect 29880 18912 29886 18924
rect 31573 18921 31585 18924
rect 31619 18921 31631 18955
rect 31573 18915 31631 18921
rect 34701 18955 34759 18961
rect 34701 18921 34713 18955
rect 34747 18952 34759 18955
rect 34790 18952 34796 18964
rect 34747 18924 34796 18952
rect 34747 18921 34759 18924
rect 34701 18915 34759 18921
rect 34790 18912 34796 18924
rect 34848 18912 34854 18964
rect 35066 18912 35072 18964
rect 35124 18952 35130 18964
rect 36262 18952 36268 18964
rect 35124 18924 36268 18952
rect 35124 18912 35130 18924
rect 36262 18912 36268 18924
rect 36320 18952 36326 18964
rect 37642 18952 37648 18964
rect 36320 18924 37648 18952
rect 36320 18912 36326 18924
rect 37642 18912 37648 18924
rect 37700 18952 37706 18964
rect 38470 18952 38476 18964
rect 37700 18924 38476 18952
rect 37700 18912 37706 18924
rect 38470 18912 38476 18924
rect 38528 18912 38534 18964
rect 30650 18884 30656 18896
rect 29840 18856 30656 18884
rect 27430 18816 27436 18828
rect 25332 18788 27436 18816
rect 25332 18757 25360 18788
rect 27430 18776 27436 18788
rect 27488 18776 27494 18828
rect 29840 18825 29868 18856
rect 30650 18844 30656 18856
rect 30708 18844 30714 18896
rect 31021 18887 31079 18893
rect 31021 18853 31033 18887
rect 31067 18884 31079 18887
rect 31110 18884 31116 18896
rect 31067 18856 31116 18884
rect 31067 18853 31079 18856
rect 31021 18847 31079 18853
rect 31110 18844 31116 18856
rect 31168 18844 31174 18896
rect 35081 18856 35204 18884
rect 29825 18819 29883 18825
rect 29825 18785 29837 18819
rect 29871 18785 29883 18819
rect 29825 18779 29883 18785
rect 30374 18776 30380 18828
rect 30432 18816 30438 18828
rect 31938 18816 31944 18828
rect 30432 18788 31944 18816
rect 30432 18776 30438 18788
rect 31938 18776 31944 18788
rect 31996 18776 32002 18828
rect 33781 18819 33839 18825
rect 33781 18785 33793 18819
rect 33827 18816 33839 18819
rect 35081 18816 35109 18856
rect 33827 18788 35109 18816
rect 33827 18785 33839 18788
rect 33781 18779 33839 18785
rect 24944 18751 25002 18757
rect 24944 18717 24956 18751
rect 24990 18717 25002 18751
rect 24944 18711 25002 18717
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18717 25099 18751
rect 25041 18711 25099 18717
rect 25316 18751 25374 18757
rect 25316 18717 25328 18751
rect 25362 18717 25374 18751
rect 25316 18711 25374 18717
rect 12529 18683 12587 18689
rect 12529 18649 12541 18683
rect 12575 18680 12587 18683
rect 13078 18680 13084 18692
rect 12575 18652 13084 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 13078 18640 13084 18652
rect 13136 18640 13142 18692
rect 15010 18640 15016 18692
rect 15068 18680 15074 18692
rect 15933 18683 15991 18689
rect 15933 18680 15945 18683
rect 15068 18652 15945 18680
rect 15068 18640 15074 18652
rect 15933 18649 15945 18652
rect 15979 18680 15991 18683
rect 19978 18680 19984 18692
rect 15979 18652 19984 18680
rect 15979 18649 15991 18652
rect 15933 18643 15991 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 20088 18652 24808 18680
rect 5316 18584 10548 18612
rect 10781 18615 10839 18621
rect 5316 18572 5322 18584
rect 10781 18581 10793 18615
rect 10827 18612 10839 18615
rect 10870 18612 10876 18624
rect 10827 18584 10876 18612
rect 10827 18581 10839 18584
rect 10781 18575 10839 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 12897 18615 12955 18621
rect 12897 18581 12909 18615
rect 12943 18612 12955 18615
rect 13722 18612 13728 18624
rect 12943 18584 13728 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 15562 18572 15568 18624
rect 15620 18612 15626 18624
rect 18138 18612 18144 18624
rect 15620 18584 18144 18612
rect 15620 18572 15626 18584
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 18690 18572 18696 18624
rect 18748 18612 18754 18624
rect 20088 18612 20116 18652
rect 22278 18612 22284 18624
rect 18748 18584 20116 18612
rect 22239 18584 22284 18612
rect 18748 18572 18754 18584
rect 22278 18572 22284 18584
rect 22336 18612 22342 18624
rect 22922 18612 22928 18624
rect 22336 18584 22928 18612
rect 22336 18572 22342 18584
rect 22922 18572 22928 18584
rect 22980 18572 22986 18624
rect 24780 18621 24808 18652
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18581 24823 18615
rect 24964 18612 24992 18711
rect 25406 18708 25412 18760
rect 25464 18748 25470 18760
rect 26694 18748 26700 18760
rect 25464 18720 25509 18748
rect 26655 18720 26700 18748
rect 25464 18708 25470 18720
rect 26694 18708 26700 18720
rect 26752 18708 26758 18760
rect 27525 18751 27583 18757
rect 27525 18717 27537 18751
rect 27571 18748 27583 18751
rect 27614 18748 27620 18760
rect 27571 18720 27620 18748
rect 27571 18717 27583 18720
rect 27525 18711 27583 18717
rect 27614 18708 27620 18720
rect 27672 18708 27678 18760
rect 28534 18708 28540 18760
rect 28592 18748 28598 18760
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 28592 18720 29561 18748
rect 28592 18708 28598 18720
rect 29549 18717 29561 18720
rect 29595 18717 29607 18751
rect 30834 18748 30840 18760
rect 30795 18720 30840 18748
rect 29549 18711 29607 18717
rect 30834 18708 30840 18720
rect 30892 18708 30898 18760
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32398 18748 32404 18760
rect 32272 18720 32404 18748
rect 32272 18708 32278 18720
rect 32398 18708 32404 18720
rect 32456 18748 32462 18760
rect 32953 18751 33011 18757
rect 32953 18748 32965 18751
rect 32456 18720 32965 18748
rect 32456 18708 32462 18720
rect 32953 18717 32965 18720
rect 32999 18717 33011 18751
rect 32953 18711 33011 18717
rect 34238 18708 34244 18760
rect 34296 18748 34302 18760
rect 34931 18751 34989 18757
rect 34931 18748 34943 18751
rect 34296 18720 34943 18748
rect 34296 18708 34302 18720
rect 34931 18717 34943 18720
rect 34977 18717 34989 18751
rect 35063 18748 35069 18760
rect 35024 18720 35069 18748
rect 34931 18711 34989 18717
rect 35063 18708 35069 18720
rect 35121 18708 35127 18760
rect 35176 18757 35204 18856
rect 36078 18816 36084 18828
rect 35268 18788 36084 18816
rect 35166 18751 35224 18757
rect 35166 18717 35178 18751
rect 35212 18717 35224 18751
rect 35166 18711 35224 18717
rect 25130 18680 25136 18692
rect 25091 18652 25136 18680
rect 25130 18640 25136 18652
rect 25188 18680 25194 18692
rect 26142 18680 26148 18692
rect 25188 18652 26148 18680
rect 25188 18640 25194 18652
rect 26142 18640 26148 18652
rect 26200 18640 26206 18692
rect 26878 18640 26884 18692
rect 26936 18680 26942 18692
rect 27798 18689 27804 18692
rect 26936 18652 27476 18680
rect 26936 18640 26942 18652
rect 25682 18612 25688 18624
rect 24964 18584 25688 18612
rect 24765 18575 24823 18581
rect 25682 18572 25688 18584
rect 25740 18572 25746 18624
rect 27065 18615 27123 18621
rect 27065 18581 27077 18615
rect 27111 18612 27123 18615
rect 27338 18612 27344 18624
rect 27111 18584 27344 18612
rect 27111 18581 27123 18584
rect 27065 18575 27123 18581
rect 27338 18572 27344 18584
rect 27396 18572 27402 18624
rect 27448 18612 27476 18652
rect 27792 18643 27804 18689
rect 27856 18680 27862 18692
rect 27856 18652 27892 18680
rect 27798 18640 27804 18643
rect 27856 18640 27862 18652
rect 30742 18640 30748 18692
rect 30800 18680 30806 18692
rect 32686 18683 32744 18689
rect 32686 18680 32698 18683
rect 30800 18652 32698 18680
rect 30800 18640 30806 18652
rect 32686 18649 32698 18652
rect 32732 18649 32744 18683
rect 33962 18680 33968 18692
rect 33923 18652 33968 18680
rect 32686 18643 32744 18649
rect 33962 18640 33968 18652
rect 34020 18640 34026 18692
rect 34149 18683 34207 18689
rect 34149 18649 34161 18683
rect 34195 18680 34207 18683
rect 35268 18680 35296 18788
rect 36078 18776 36084 18788
rect 36136 18776 36142 18828
rect 35345 18751 35403 18757
rect 35345 18717 35357 18751
rect 35391 18717 35403 18751
rect 35345 18711 35403 18717
rect 34195 18652 35296 18680
rect 34195 18649 34207 18652
rect 34149 18643 34207 18649
rect 28905 18615 28963 18621
rect 28905 18612 28917 18615
rect 27448 18584 28917 18612
rect 28905 18581 28917 18584
rect 28951 18581 28963 18615
rect 28905 18575 28963 18581
rect 34054 18572 34060 18624
rect 34112 18612 34118 18624
rect 35360 18612 35388 18711
rect 37274 18708 37280 18760
rect 37332 18757 37338 18760
rect 37332 18748 37344 18757
rect 37332 18720 37377 18748
rect 37332 18711 37344 18720
rect 37332 18708 37338 18711
rect 37458 18708 37464 18760
rect 37516 18748 37522 18760
rect 37553 18751 37611 18757
rect 37553 18748 37565 18751
rect 37516 18720 37565 18748
rect 37516 18708 37522 18720
rect 37553 18717 37565 18720
rect 37599 18717 37611 18751
rect 68094 18748 68100 18760
rect 68055 18720 68100 18748
rect 37553 18711 37611 18717
rect 68094 18708 68100 18720
rect 68152 18708 68158 18760
rect 34112 18584 35388 18612
rect 36173 18615 36231 18621
rect 34112 18572 34118 18584
rect 36173 18581 36185 18615
rect 36219 18612 36231 18615
rect 36262 18612 36268 18624
rect 36219 18584 36268 18612
rect 36219 18581 36231 18584
rect 36173 18575 36231 18581
rect 36262 18572 36268 18584
rect 36320 18572 36326 18624
rect 37274 18572 37280 18624
rect 37332 18612 37338 18624
rect 37550 18612 37556 18624
rect 37332 18584 37556 18612
rect 37332 18572 37338 18584
rect 37550 18572 37556 18584
rect 37608 18612 37614 18624
rect 38013 18615 38071 18621
rect 38013 18612 38025 18615
rect 37608 18584 38025 18612
rect 37608 18572 37614 18584
rect 38013 18581 38025 18584
rect 38059 18581 38071 18615
rect 38013 18575 38071 18581
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 7285 18411 7343 18417
rect 7285 18408 7297 18411
rect 6972 18380 7297 18408
rect 6972 18368 6978 18380
rect 7285 18377 7297 18380
rect 7331 18377 7343 18411
rect 10134 18408 10140 18420
rect 7285 18371 7343 18377
rect 7484 18380 10140 18408
rect 7484 18349 7512 18380
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10318 18408 10324 18420
rect 10279 18380 10324 18408
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 13173 18411 13231 18417
rect 10428 18380 12112 18408
rect 2777 18343 2835 18349
rect 2777 18309 2789 18343
rect 2823 18340 2835 18343
rect 3850 18343 3908 18349
rect 3850 18340 3862 18343
rect 2823 18312 3862 18340
rect 2823 18309 2835 18312
rect 2777 18303 2835 18309
rect 3850 18309 3862 18312
rect 3896 18309 3908 18343
rect 3850 18303 3908 18309
rect 7469 18343 7527 18349
rect 7469 18309 7481 18343
rect 7515 18309 7527 18343
rect 7650 18340 7656 18352
rect 7611 18312 7656 18340
rect 7469 18303 7527 18309
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 8846 18300 8852 18352
rect 8904 18340 8910 18352
rect 10428 18340 10456 18380
rect 8904 18312 10456 18340
rect 10505 18343 10563 18349
rect 8904 18300 8910 18312
rect 10505 18309 10517 18343
rect 10551 18340 10563 18343
rect 11974 18340 11980 18352
rect 10551 18312 11980 18340
rect 10551 18309 10563 18312
rect 10505 18303 10563 18309
rect 11974 18300 11980 18312
rect 12032 18300 12038 18352
rect 2130 18272 2136 18284
rect 2091 18244 2136 18272
rect 2130 18232 2136 18244
rect 2188 18232 2194 18284
rect 2314 18272 2320 18284
rect 2275 18244 2320 18272
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18241 2467 18275
rect 2409 18235 2467 18241
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 3234 18272 3240 18284
rect 2547 18244 3240 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2424 18204 2452 18235
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 7558 18272 7564 18284
rect 6687 18244 7564 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 7668 18272 7696 18300
rect 12084 18284 12112 18380
rect 13173 18377 13185 18411
rect 13219 18408 13231 18411
rect 13814 18408 13820 18420
rect 13219 18380 13820 18408
rect 13219 18377 13231 18380
rect 13173 18371 13231 18377
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 15010 18408 15016 18420
rect 14971 18380 15016 18408
rect 15010 18368 15016 18380
rect 15068 18368 15074 18420
rect 16117 18411 16175 18417
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 17402 18408 17408 18420
rect 16163 18380 17408 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 19981 18411 20039 18417
rect 19981 18408 19993 18411
rect 17604 18380 19993 18408
rect 15562 18340 15568 18352
rect 12544 18312 13584 18340
rect 8110 18272 8116 18284
rect 7668 18244 8116 18272
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 9582 18272 9588 18284
rect 8220 18244 9588 18272
rect 3602 18204 3608 18216
rect 2280 18176 2452 18204
rect 3563 18176 3608 18204
rect 2280 18164 2286 18176
rect 3602 18164 3608 18176
rect 3660 18164 3666 18216
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 6457 18207 6515 18213
rect 6457 18204 6469 18207
rect 5868 18176 6469 18204
rect 5868 18164 5874 18176
rect 6457 18173 6469 18176
rect 6503 18204 6515 18207
rect 7282 18204 7288 18216
rect 6503 18176 7288 18204
rect 6503 18173 6515 18176
rect 6457 18167 6515 18173
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 5350 18096 5356 18148
rect 5408 18136 5414 18148
rect 8220 18136 8248 18244
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 10226 18232 10232 18284
rect 10284 18272 10290 18284
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10284 18244 10701 18272
rect 10284 18232 10290 18244
rect 10689 18241 10701 18244
rect 10735 18241 10747 18275
rect 10689 18235 10747 18241
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 12544 18281 12572 18312
rect 12345 18275 12403 18281
rect 12345 18272 12357 18275
rect 12124 18244 12357 18272
rect 12124 18232 12130 18244
rect 12345 18241 12357 18244
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 12768 18244 13093 18272
rect 12768 18232 12774 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 10244 18204 10272 18232
rect 5408 18108 8248 18136
rect 8312 18176 10272 18204
rect 12437 18207 12495 18213
rect 5408 18096 5414 18108
rect 4985 18071 5043 18077
rect 4985 18037 4997 18071
rect 5031 18068 5043 18071
rect 5442 18068 5448 18080
rect 5031 18040 5448 18068
rect 5031 18037 5043 18040
rect 4985 18031 5043 18037
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 8312 18077 8340 18176
rect 12437 18173 12449 18207
rect 12483 18204 12495 18207
rect 12728 18204 12756 18232
rect 12483 18176 12756 18204
rect 13556 18204 13584 18312
rect 13832 18312 15568 18340
rect 13722 18272 13728 18284
rect 13683 18244 13728 18272
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 13832 18281 13860 18312
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 17221 18343 17279 18349
rect 17221 18309 17233 18343
rect 17267 18340 17279 18343
rect 17604 18340 17632 18380
rect 19981 18377 19993 18380
rect 20027 18408 20039 18411
rect 24305 18411 24363 18417
rect 20027 18380 22094 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 17267 18312 17632 18340
rect 17267 18309 17279 18312
rect 17221 18303 17279 18309
rect 17678 18300 17684 18352
rect 17736 18340 17742 18352
rect 18846 18343 18904 18349
rect 18846 18340 18858 18343
rect 17736 18312 18858 18340
rect 17736 18300 17742 18312
rect 18846 18309 18858 18312
rect 18892 18309 18904 18343
rect 20714 18340 20720 18352
rect 18846 18303 18904 18309
rect 20456 18312 20720 18340
rect 13818 18275 13876 18281
rect 13818 18241 13830 18275
rect 13864 18241 13876 18275
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 13818 18235 13876 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14231 18275 14289 18281
rect 14148 18244 14193 18272
rect 14148 18232 14154 18244
rect 14231 18241 14243 18275
rect 14277 18272 14289 18275
rect 14366 18272 14372 18284
rect 14277 18244 14372 18272
rect 14277 18241 14289 18244
rect 14231 18235 14289 18241
rect 14366 18232 14372 18244
rect 14424 18272 14430 18284
rect 15102 18272 15108 18284
rect 14424 18244 15108 18272
rect 14424 18232 14430 18244
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 15344 18244 15485 18272
rect 15344 18232 15350 18244
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15654 18272 15660 18284
rect 15615 18244 15660 18272
rect 15473 18235 15531 18241
rect 14734 18204 14740 18216
rect 13556 18176 14740 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 15488 18204 15516 18235
rect 15654 18232 15660 18244
rect 15712 18232 15718 18284
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 15562 18204 15568 18216
rect 15488 18176 15568 18204
rect 15562 18164 15568 18176
rect 15620 18164 15626 18216
rect 15764 18204 15792 18235
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 15896 18244 15941 18272
rect 15896 18232 15902 18244
rect 16850 18232 16856 18284
rect 16908 18272 16914 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 16908 18244 17049 18272
rect 16908 18232 16914 18244
rect 17037 18241 17049 18244
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 17310 18232 17316 18284
rect 17368 18272 17374 18284
rect 20456 18281 20484 18312
rect 20714 18300 20720 18312
rect 20772 18300 20778 18352
rect 22066 18340 22094 18380
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 25406 18408 25412 18420
rect 24351 18380 25412 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 27798 18408 27804 18420
rect 27759 18380 27804 18408
rect 27798 18368 27804 18380
rect 27856 18368 27862 18420
rect 30742 18408 30748 18420
rect 30703 18380 30748 18408
rect 30742 18368 30748 18380
rect 30800 18368 30806 18420
rect 32582 18368 32588 18420
rect 32640 18408 32646 18420
rect 34238 18408 34244 18420
rect 32640 18380 34244 18408
rect 32640 18368 32646 18380
rect 34238 18368 34244 18380
rect 34296 18368 34302 18420
rect 36446 18408 36452 18420
rect 36407 18380 36452 18408
rect 36446 18368 36452 18380
rect 36504 18368 36510 18420
rect 24029 18343 24087 18349
rect 24029 18340 24041 18343
rect 22066 18312 24041 18340
rect 24029 18309 24041 18312
rect 24075 18309 24087 18343
rect 24029 18303 24087 18309
rect 24210 18300 24216 18352
rect 24268 18340 24274 18352
rect 25041 18343 25099 18349
rect 25041 18340 25053 18343
rect 24268 18312 25053 18340
rect 24268 18300 24274 18312
rect 25041 18309 25053 18312
rect 25087 18309 25099 18343
rect 32217 18343 32275 18349
rect 25041 18303 25099 18309
rect 27172 18312 28672 18340
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 17368 18244 18613 18272
rect 17368 18232 17374 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 20622 18232 20628 18284
rect 20680 18272 20686 18284
rect 23014 18272 23020 18284
rect 20680 18244 23020 18272
rect 20680 18232 20686 18244
rect 23014 18232 23020 18244
rect 23072 18232 23078 18284
rect 23750 18272 23756 18284
rect 23711 18244 23756 18272
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 23934 18232 23940 18284
rect 23992 18272 23998 18284
rect 23992 18244 24085 18272
rect 23992 18232 23998 18244
rect 24118 18232 24124 18284
rect 24176 18272 24182 18284
rect 24762 18272 24768 18284
rect 24176 18244 24221 18272
rect 24723 18244 24768 18272
rect 24176 18232 24182 18244
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18241 25007 18275
rect 25133 18275 25191 18281
rect 25133 18272 25145 18275
rect 24949 18235 25007 18241
rect 25056 18244 25145 18272
rect 16022 18204 16028 18216
rect 15764 18176 16028 18204
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 20717 18207 20775 18213
rect 20717 18173 20729 18207
rect 20763 18173 20775 18207
rect 20717 18167 20775 18173
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 12802 18136 12808 18148
rect 9732 18108 12808 18136
rect 9732 18096 9738 18108
rect 12802 18096 12808 18108
rect 12860 18096 12866 18148
rect 14752 18136 14780 18164
rect 20732 18136 20760 18167
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 22462 18204 22468 18216
rect 22152 18176 22468 18204
rect 22152 18164 22158 18176
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 22738 18204 22744 18216
rect 22699 18176 22744 18204
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 23952 18204 23980 18232
rect 24964 18204 24992 18235
rect 23952 18176 24992 18204
rect 14752 18108 18644 18136
rect 8297 18071 8355 18077
rect 8297 18037 8309 18071
rect 8343 18037 8355 18071
rect 9214 18068 9220 18080
rect 9175 18040 9220 18068
rect 8297 18031 8355 18037
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18068 9919 18071
rect 10042 18068 10048 18080
rect 9907 18040 10048 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 14090 18068 14096 18080
rect 12032 18040 14096 18068
rect 12032 18028 12038 18040
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 14369 18071 14427 18077
rect 14369 18037 14381 18071
rect 14415 18068 14427 18071
rect 17126 18068 17132 18080
rect 14415 18040 17132 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 17405 18071 17463 18077
rect 17405 18068 17417 18071
rect 17276 18040 17417 18068
rect 17276 18028 17282 18040
rect 17405 18037 17417 18040
rect 17451 18037 17463 18071
rect 17405 18031 17463 18037
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17644 18040 18061 18068
rect 17644 18028 17650 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18616 18068 18644 18108
rect 19536 18108 20760 18136
rect 19536 18080 19564 18108
rect 24118 18096 24124 18148
rect 24176 18136 24182 18148
rect 25056 18136 25084 18244
rect 25133 18241 25145 18244
rect 25179 18241 25191 18275
rect 25133 18235 25191 18241
rect 26970 18232 26976 18284
rect 27028 18272 27034 18284
rect 27172 18281 27200 18312
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 27028 18244 27169 18272
rect 27028 18232 27034 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 27157 18235 27215 18241
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 27433 18275 27491 18281
rect 27433 18241 27445 18275
rect 27479 18241 27491 18275
rect 27433 18235 27491 18241
rect 27571 18275 27629 18281
rect 27571 18241 27583 18275
rect 27617 18272 27629 18275
rect 27982 18272 27988 18284
rect 27617 18244 27988 18272
rect 27617 18241 27629 18244
rect 27571 18235 27629 18241
rect 25774 18204 25780 18216
rect 25735 18176 25780 18204
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 27448 18204 27476 18235
rect 27982 18232 27988 18244
rect 28040 18232 28046 18284
rect 28534 18272 28540 18284
rect 28495 18244 28540 18272
rect 28534 18232 28540 18244
rect 28592 18232 28598 18284
rect 28644 18272 28672 18312
rect 32217 18309 32229 18343
rect 32263 18340 32275 18343
rect 32769 18343 32827 18349
rect 32769 18340 32781 18343
rect 32263 18312 32781 18340
rect 32263 18309 32275 18312
rect 32217 18303 32275 18309
rect 32769 18309 32781 18312
rect 32815 18340 32827 18343
rect 34422 18340 34428 18352
rect 32815 18312 34428 18340
rect 32815 18309 32827 18312
rect 32769 18303 32827 18309
rect 34422 18300 34428 18312
rect 34480 18300 34486 18352
rect 36078 18340 36084 18352
rect 36039 18312 36084 18340
rect 36078 18300 36084 18312
rect 36136 18300 36142 18352
rect 30098 18272 30104 18284
rect 30156 18281 30162 18284
rect 28644 18244 30104 18272
rect 30098 18232 30104 18244
rect 30156 18272 30165 18281
rect 30282 18272 30288 18284
rect 30156 18244 30201 18272
rect 30243 18244 30288 18272
rect 30156 18235 30165 18244
rect 30156 18232 30162 18235
rect 30282 18232 30288 18244
rect 30340 18232 30346 18284
rect 30377 18275 30435 18281
rect 30377 18241 30389 18275
rect 30423 18241 30435 18275
rect 30377 18235 30435 18241
rect 30469 18275 30527 18281
rect 30469 18241 30481 18275
rect 30515 18241 30527 18275
rect 35066 18272 35072 18284
rect 35027 18244 35072 18272
rect 30469 18235 30527 18241
rect 27706 18204 27712 18216
rect 27448 18176 27712 18204
rect 27706 18164 27712 18176
rect 27764 18204 27770 18216
rect 28813 18207 28871 18213
rect 28813 18204 28825 18207
rect 27764 18176 28825 18204
rect 27764 18164 27770 18176
rect 28813 18173 28825 18176
rect 28859 18204 28871 18207
rect 30392 18204 30420 18235
rect 28859 18176 30420 18204
rect 28859 18173 28871 18176
rect 28813 18167 28871 18173
rect 24176 18108 25084 18136
rect 25317 18139 25375 18145
rect 24176 18096 24182 18108
rect 25317 18105 25329 18139
rect 25363 18136 25375 18139
rect 26142 18136 26148 18148
rect 25363 18108 26148 18136
rect 25363 18105 25375 18108
rect 25317 18099 25375 18105
rect 26142 18096 26148 18108
rect 26200 18096 26206 18148
rect 30374 18136 30380 18148
rect 28966 18108 30380 18136
rect 19518 18068 19524 18080
rect 18616 18040 19524 18068
rect 18049 18031 18107 18037
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 20990 18028 20996 18080
rect 21048 18068 21054 18080
rect 21913 18071 21971 18077
rect 21913 18068 21925 18071
rect 21048 18040 21925 18068
rect 21048 18028 21054 18040
rect 21913 18037 21925 18040
rect 21959 18068 21971 18071
rect 22554 18068 22560 18080
rect 21959 18040 22560 18068
rect 21959 18037 21971 18040
rect 21913 18031 21971 18037
rect 22554 18028 22560 18040
rect 22612 18028 22618 18080
rect 22738 18028 22744 18080
rect 22796 18068 22802 18080
rect 25130 18068 25136 18080
rect 22796 18040 25136 18068
rect 22796 18028 22802 18040
rect 25130 18028 25136 18040
rect 25188 18028 25194 18080
rect 25866 18028 25872 18080
rect 25924 18068 25930 18080
rect 28966 18068 28994 18108
rect 30374 18096 30380 18108
rect 30432 18096 30438 18148
rect 25924 18040 28994 18068
rect 25924 18028 25930 18040
rect 30282 18028 30288 18080
rect 30340 18068 30346 18080
rect 30484 18068 30512 18235
rect 35066 18232 35072 18244
rect 35124 18232 35130 18284
rect 36262 18272 36268 18284
rect 36223 18244 36268 18272
rect 36262 18232 36268 18244
rect 36320 18232 36326 18284
rect 37458 18232 37464 18284
rect 37516 18272 37522 18284
rect 38010 18281 38016 18284
rect 37737 18275 37795 18281
rect 37737 18272 37749 18275
rect 37516 18244 37749 18272
rect 37516 18232 37522 18244
rect 37737 18241 37749 18244
rect 37783 18241 37795 18275
rect 37737 18235 37795 18241
rect 38004 18235 38016 18281
rect 38068 18272 38074 18284
rect 38068 18244 38104 18272
rect 38010 18232 38016 18235
rect 38068 18232 38074 18244
rect 34790 18204 34796 18216
rect 34751 18176 34796 18204
rect 34790 18164 34796 18176
rect 34848 18164 34854 18216
rect 32953 18139 33011 18145
rect 32953 18105 32965 18139
rect 32999 18136 33011 18139
rect 34054 18136 34060 18148
rect 32999 18108 34060 18136
rect 32999 18105 33011 18108
rect 32953 18099 33011 18105
rect 34054 18096 34060 18108
rect 34112 18096 34118 18148
rect 31205 18071 31263 18077
rect 31205 18068 31217 18071
rect 30340 18040 31217 18068
rect 30340 18028 30346 18040
rect 31205 18037 31217 18040
rect 31251 18037 31263 18071
rect 31205 18031 31263 18037
rect 38746 18028 38752 18080
rect 38804 18068 38810 18080
rect 39117 18071 39175 18077
rect 39117 18068 39129 18071
rect 38804 18040 39129 18068
rect 38804 18028 38810 18040
rect 39117 18037 39129 18040
rect 39163 18037 39175 18071
rect 39117 18031 39175 18037
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 1489 17867 1547 17873
rect 1489 17833 1501 17867
rect 1535 17864 1547 17867
rect 1535 17836 2360 17864
rect 1535 17833 1547 17836
rect 1489 17827 1547 17833
rect 2222 17756 2228 17808
rect 2280 17756 2286 17808
rect 1949 17663 2007 17669
rect 1949 17629 1961 17663
rect 1995 17660 2007 17663
rect 2038 17660 2044 17672
rect 1995 17632 2044 17660
rect 1995 17629 2007 17632
rect 1949 17623 2007 17629
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 2240 17669 2268 17756
rect 2332 17669 2360 17836
rect 8110 17824 8116 17876
rect 8168 17864 8174 17876
rect 8941 17867 8999 17873
rect 8941 17864 8953 17867
rect 8168 17836 8953 17864
rect 8168 17824 8174 17836
rect 8941 17833 8953 17836
rect 8987 17833 8999 17867
rect 11698 17864 11704 17876
rect 8941 17827 8999 17833
rect 9646 17836 11704 17864
rect 7742 17756 7748 17808
rect 7800 17796 7806 17808
rect 8018 17796 8024 17808
rect 7800 17768 8024 17796
rect 7800 17756 7806 17768
rect 8018 17756 8024 17768
rect 8076 17796 8082 17808
rect 9646 17796 9674 17836
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 11974 17864 11980 17876
rect 11935 17836 11980 17864
rect 11974 17824 11980 17836
rect 12032 17824 12038 17876
rect 12158 17824 12164 17876
rect 12216 17864 12222 17876
rect 14826 17864 14832 17876
rect 12216 17836 14832 17864
rect 12216 17824 12222 17836
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 14921 17867 14979 17873
rect 14921 17833 14933 17867
rect 14967 17864 14979 17867
rect 15470 17864 15476 17876
rect 14967 17836 15476 17864
rect 14967 17833 14979 17836
rect 14921 17827 14979 17833
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 15746 17864 15752 17876
rect 15707 17836 15752 17864
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 17678 17864 17684 17876
rect 17639 17836 17684 17864
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 20898 17824 20904 17876
rect 20956 17864 20962 17876
rect 21450 17864 21456 17876
rect 20956 17836 21456 17864
rect 20956 17824 20962 17836
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 21634 17824 21640 17876
rect 21692 17864 21698 17876
rect 23566 17864 23572 17876
rect 21692 17836 23572 17864
rect 21692 17824 21698 17836
rect 23566 17824 23572 17836
rect 23624 17864 23630 17876
rect 28810 17864 28816 17876
rect 23624 17836 24532 17864
rect 28771 17836 28816 17864
rect 23624 17824 23630 17836
rect 14366 17796 14372 17808
rect 8076 17768 9674 17796
rect 12406 17768 14372 17796
rect 8076 17756 8082 17768
rect 3602 17688 3608 17740
rect 3660 17728 3666 17740
rect 5350 17728 5356 17740
rect 3660 17700 5356 17728
rect 3660 17688 3666 17700
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 7098 17688 7104 17740
rect 7156 17728 7162 17740
rect 9214 17728 9220 17740
rect 7156 17700 9220 17728
rect 7156 17688 7162 17700
rect 9214 17688 9220 17700
rect 9272 17728 9278 17740
rect 9309 17731 9367 17737
rect 9309 17728 9321 17731
rect 9272 17700 9321 17728
rect 9272 17688 9278 17700
rect 9309 17697 9321 17700
rect 9355 17697 9367 17731
rect 9309 17691 9367 17697
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17629 2191 17663
rect 2133 17623 2191 17629
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 2682 17660 2688 17672
rect 2363 17632 2688 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 2148 17592 2176 17623
rect 2682 17620 2688 17632
rect 2740 17660 2746 17672
rect 6822 17660 6828 17672
rect 2740 17632 6828 17660
rect 2740 17620 2746 17632
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 2774 17592 2780 17604
rect 2148 17564 2780 17592
rect 2774 17552 2780 17564
rect 2832 17552 2838 17604
rect 2958 17552 2964 17604
rect 3016 17592 3022 17604
rect 5598 17595 5656 17601
rect 5598 17592 5610 17595
rect 3016 17564 5610 17592
rect 3016 17552 3022 17564
rect 5598 17561 5610 17564
rect 5644 17561 5656 17595
rect 5598 17555 5656 17561
rect 2590 17524 2596 17536
rect 2551 17496 2596 17524
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 2682 17484 2688 17536
rect 2740 17524 2746 17536
rect 5442 17524 5448 17536
rect 2740 17496 5448 17524
rect 2740 17484 2746 17496
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 6730 17524 6736 17536
rect 6691 17496 6736 17524
rect 6730 17484 6736 17496
rect 6788 17484 6794 17536
rect 7208 17524 7236 17623
rect 7282 17620 7288 17672
rect 7340 17660 7346 17672
rect 7469 17663 7527 17669
rect 7469 17660 7481 17663
rect 7340 17632 7481 17660
rect 7340 17620 7346 17632
rect 7469 17629 7481 17632
rect 7515 17629 7527 17663
rect 7469 17623 7527 17629
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17629 9183 17663
rect 9324 17660 9352 17691
rect 9582 17688 9588 17740
rect 9640 17728 9646 17740
rect 10597 17731 10655 17737
rect 10597 17728 10609 17731
rect 9640 17700 10609 17728
rect 9640 17688 9646 17700
rect 10597 17697 10609 17700
rect 10643 17697 10655 17731
rect 10597 17691 10655 17697
rect 9858 17660 9864 17672
rect 9324 17632 9864 17660
rect 9125 17623 9183 17629
rect 9140 17592 9168 17623
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 10042 17660 10048 17672
rect 9999 17632 10048 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 10042 17620 10048 17632
rect 10100 17620 10106 17672
rect 10870 17669 10876 17672
rect 10864 17660 10876 17669
rect 10831 17632 10876 17660
rect 10864 17623 10876 17632
rect 10870 17620 10876 17623
rect 10928 17620 10934 17672
rect 12406 17592 12434 17768
rect 14366 17756 14372 17768
rect 14424 17756 14430 17808
rect 16666 17756 16672 17808
rect 16724 17796 16730 17808
rect 20806 17796 20812 17808
rect 16724 17768 17448 17796
rect 16724 17756 16730 17768
rect 16022 17728 16028 17740
rect 13004 17700 16028 17728
rect 13004 17672 13032 17700
rect 16022 17688 16028 17700
rect 16080 17728 16086 17740
rect 16080 17700 17356 17728
rect 16080 17688 16086 17700
rect 12710 17660 12716 17672
rect 12671 17632 12716 17660
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 12986 17660 12992 17672
rect 12947 17632 12992 17660
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 14553 17663 14611 17669
rect 14553 17629 14565 17663
rect 14599 17629 14611 17663
rect 14734 17660 14740 17672
rect 14695 17632 14740 17660
rect 14553 17623 14611 17629
rect 9140 17564 12434 17592
rect 13446 17552 13452 17604
rect 13504 17592 13510 17604
rect 14568 17592 14596 17623
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 15930 17660 15936 17672
rect 15891 17632 15936 17660
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 17037 17663 17095 17669
rect 17037 17660 17049 17663
rect 17000 17632 17049 17660
rect 17000 17620 17006 17632
rect 17037 17629 17049 17632
rect 17083 17629 17095 17663
rect 17218 17660 17224 17672
rect 17179 17632 17224 17660
rect 17037 17623 17095 17629
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 17328 17669 17356 17700
rect 17420 17669 17448 17768
rect 20640 17768 20812 17796
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 13504 17564 14596 17592
rect 16117 17595 16175 17601
rect 13504 17552 13510 17564
rect 16117 17561 16129 17595
rect 16163 17592 16175 17595
rect 16850 17592 16856 17604
rect 16163 17564 16856 17592
rect 16163 17561 16175 17564
rect 16117 17555 16175 17561
rect 16850 17552 16856 17564
rect 16908 17552 16914 17604
rect 17328 17592 17356 17623
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 17644 17632 19809 17660
rect 17644 17620 17650 17632
rect 19797 17629 19809 17632
rect 19843 17660 19855 17663
rect 20162 17660 20168 17672
rect 19843 17632 20168 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 20162 17620 20168 17632
rect 20220 17620 20226 17672
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 20640 17669 20668 17768
rect 20806 17756 20812 17768
rect 20864 17756 20870 17808
rect 20993 17799 21051 17805
rect 20993 17765 21005 17799
rect 21039 17796 21051 17799
rect 22462 17796 22468 17808
rect 21039 17768 22468 17796
rect 21039 17765 21051 17768
rect 20993 17759 21051 17765
rect 22462 17756 22468 17768
rect 22520 17756 22526 17808
rect 24504 17805 24532 17836
rect 28810 17824 28816 17836
rect 28868 17824 28874 17876
rect 29822 17824 29828 17876
rect 29880 17864 29886 17876
rect 33962 17864 33968 17876
rect 29880 17836 33968 17864
rect 29880 17824 29886 17836
rect 33962 17824 33968 17836
rect 34020 17824 34026 17876
rect 34606 17864 34612 17876
rect 34348 17836 34612 17864
rect 24489 17799 24547 17805
rect 24489 17765 24501 17799
rect 24535 17796 24547 17799
rect 26234 17796 26240 17808
rect 24535 17768 26240 17796
rect 24535 17765 24547 17768
rect 24489 17759 24547 17765
rect 26234 17756 26240 17768
rect 26292 17796 26298 17808
rect 29454 17796 29460 17808
rect 26292 17768 29460 17796
rect 26292 17756 26298 17768
rect 29454 17756 29460 17768
rect 29512 17756 29518 17808
rect 32306 17756 32312 17808
rect 32364 17796 32370 17808
rect 34348 17796 34376 17836
rect 34606 17824 34612 17836
rect 34664 17824 34670 17876
rect 34885 17867 34943 17873
rect 34885 17833 34897 17867
rect 34931 17864 34943 17867
rect 36078 17864 36084 17876
rect 34931 17836 36084 17864
rect 34931 17833 34943 17836
rect 34885 17827 34943 17833
rect 36078 17824 36084 17836
rect 36136 17824 36142 17876
rect 38010 17824 38016 17876
rect 38068 17864 38074 17876
rect 38197 17867 38255 17873
rect 38197 17864 38209 17867
rect 38068 17836 38209 17864
rect 38068 17824 38074 17836
rect 38197 17833 38209 17836
rect 38243 17833 38255 17867
rect 38197 17827 38255 17833
rect 32364 17768 34376 17796
rect 32364 17756 32370 17768
rect 34422 17756 34428 17808
rect 34480 17796 34486 17808
rect 35345 17799 35403 17805
rect 35345 17796 35357 17799
rect 34480 17768 35357 17796
rect 34480 17756 34486 17768
rect 35345 17765 35357 17768
rect 35391 17765 35403 17799
rect 35345 17759 35403 17765
rect 22281 17731 22339 17737
rect 22281 17697 22293 17731
rect 22327 17728 22339 17731
rect 24118 17728 24124 17740
rect 22327 17700 24124 17728
rect 22327 17697 22339 17700
rect 22281 17691 22339 17697
rect 24118 17688 24124 17700
rect 24176 17688 24182 17740
rect 25130 17688 25136 17740
rect 25188 17728 25194 17740
rect 25188 17700 25912 17728
rect 25188 17688 25194 17700
rect 20441 17663 20499 17669
rect 20441 17660 20453 17663
rect 20404 17632 20453 17660
rect 20404 17620 20410 17632
rect 20441 17629 20453 17632
rect 20487 17629 20499 17663
rect 20441 17623 20499 17629
rect 20625 17663 20683 17669
rect 20625 17629 20637 17663
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 22002 17660 22008 17672
rect 20864 17632 22008 17660
rect 20864 17620 20870 17632
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 25682 17669 25688 17672
rect 25639 17663 25688 17669
rect 25639 17660 25651 17663
rect 23308 17632 25651 17660
rect 17770 17592 17776 17604
rect 17328 17564 17776 17592
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 18693 17595 18751 17601
rect 18693 17561 18705 17595
rect 18739 17592 18751 17595
rect 19426 17592 19432 17604
rect 18739 17564 19432 17592
rect 18739 17561 18751 17564
rect 18693 17555 18751 17561
rect 19426 17552 19432 17564
rect 19484 17552 19490 17604
rect 19981 17595 20039 17601
rect 19981 17561 19993 17595
rect 20027 17592 20039 17595
rect 20530 17592 20536 17604
rect 20027 17564 20536 17592
rect 20027 17561 20039 17564
rect 19981 17555 20039 17561
rect 20530 17552 20536 17564
rect 20588 17552 20594 17604
rect 20717 17595 20775 17601
rect 20717 17561 20729 17595
rect 20763 17561 20775 17595
rect 20717 17555 20775 17561
rect 7558 17524 7564 17536
rect 7208 17496 7564 17524
rect 7558 17484 7564 17496
rect 7616 17524 7622 17536
rect 9766 17524 9772 17536
rect 7616 17496 9772 17524
rect 7616 17484 7622 17496
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 13464 17524 13492 17552
rect 9916 17496 13492 17524
rect 9916 17484 9922 17496
rect 15194 17484 15200 17536
rect 15252 17524 15258 17536
rect 20732 17524 20760 17555
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 23308 17592 23336 17632
rect 25639 17629 25651 17632
rect 25685 17629 25688 17663
rect 25639 17623 25688 17629
rect 25682 17620 25688 17623
rect 25740 17660 25746 17672
rect 25884 17669 25912 17700
rect 25958 17688 25964 17740
rect 26016 17728 26022 17740
rect 26016 17700 27614 17728
rect 26016 17688 26022 17700
rect 25869 17663 25927 17669
rect 25740 17632 25787 17660
rect 25740 17620 25746 17632
rect 25869 17629 25881 17663
rect 25915 17629 25927 17663
rect 26050 17660 26056 17672
rect 26011 17632 26056 17660
rect 25869 17623 25927 17629
rect 26050 17620 26056 17632
rect 26108 17620 26114 17672
rect 26142 17620 26148 17672
rect 26200 17660 26206 17672
rect 26605 17663 26663 17669
rect 26200 17632 26245 17660
rect 26200 17620 26206 17632
rect 26605 17629 26617 17663
rect 26651 17660 26663 17663
rect 26694 17660 26700 17672
rect 26651 17632 26700 17660
rect 26651 17629 26663 17632
rect 26605 17623 26663 17629
rect 26694 17620 26700 17632
rect 26752 17620 26758 17672
rect 26786 17620 26792 17672
rect 26844 17660 26850 17672
rect 27586 17660 27614 17700
rect 29362 17688 29368 17740
rect 29420 17728 29426 17740
rect 32214 17728 32220 17740
rect 29420 17700 30144 17728
rect 32175 17700 32220 17728
rect 29420 17688 29426 17700
rect 28997 17663 29055 17669
rect 28997 17660 29009 17663
rect 26844 17632 26889 17660
rect 27586 17632 29009 17660
rect 26844 17620 26850 17632
rect 28997 17629 29009 17632
rect 29043 17660 29055 17663
rect 29086 17660 29092 17672
rect 29043 17632 29092 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 29086 17620 29092 17632
rect 29144 17620 29150 17672
rect 29730 17660 29736 17672
rect 29691 17632 29736 17660
rect 29730 17620 29736 17632
rect 29788 17620 29794 17672
rect 29822 17620 29828 17672
rect 29880 17660 29886 17672
rect 30116 17669 30144 17700
rect 32214 17688 32220 17700
rect 32272 17688 32278 17740
rect 30101 17663 30159 17669
rect 29880 17632 29925 17660
rect 29880 17620 29886 17632
rect 30101 17629 30113 17663
rect 30147 17629 30159 17663
rect 30101 17623 30159 17629
rect 32953 17663 33011 17669
rect 32953 17629 32965 17663
rect 32999 17660 33011 17663
rect 33318 17660 33324 17672
rect 32999 17632 33324 17660
rect 32999 17629 33011 17632
rect 32953 17623 33011 17629
rect 33318 17620 33324 17632
rect 33376 17660 33382 17672
rect 33689 17663 33747 17669
rect 33689 17660 33701 17663
rect 33376 17632 33701 17660
rect 33376 17620 33382 17632
rect 33689 17629 33701 17632
rect 33735 17629 33747 17663
rect 33689 17623 33747 17629
rect 33781 17663 33839 17669
rect 33781 17629 33793 17663
rect 33827 17629 33839 17663
rect 33781 17623 33839 17629
rect 23072 17564 23336 17592
rect 23385 17595 23443 17601
rect 23072 17552 23078 17564
rect 23385 17561 23397 17595
rect 23431 17592 23443 17595
rect 24578 17592 24584 17604
rect 23431 17564 24584 17592
rect 23431 17561 23443 17564
rect 23385 17555 23443 17561
rect 24578 17552 24584 17564
rect 24636 17552 24642 17604
rect 25774 17592 25780 17604
rect 24872 17564 25636 17592
rect 25735 17564 25780 17592
rect 15252 17496 20760 17524
rect 23477 17527 23535 17533
rect 15252 17484 15258 17496
rect 23477 17493 23489 17527
rect 23523 17524 23535 17527
rect 24118 17524 24124 17536
rect 23523 17496 24124 17524
rect 23523 17493 23535 17496
rect 23477 17487 23535 17493
rect 24118 17484 24124 17496
rect 24176 17524 24182 17536
rect 24872 17524 24900 17564
rect 24176 17496 24900 17524
rect 25041 17527 25099 17533
rect 24176 17484 24182 17496
rect 25041 17493 25053 17527
rect 25087 17524 25099 17527
rect 25130 17524 25136 17536
rect 25087 17496 25136 17524
rect 25087 17493 25099 17496
rect 25041 17487 25099 17493
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 25498 17524 25504 17536
rect 25459 17496 25504 17524
rect 25498 17484 25504 17496
rect 25556 17484 25562 17536
rect 25608 17524 25636 17564
rect 25774 17552 25780 17564
rect 25832 17552 25838 17604
rect 29270 17592 29276 17604
rect 26896 17564 29276 17592
rect 26896 17524 26924 17564
rect 29270 17552 29276 17564
rect 29328 17552 29334 17604
rect 29914 17592 29920 17604
rect 29875 17564 29920 17592
rect 29914 17552 29920 17564
rect 29972 17552 29978 17604
rect 31972 17595 32030 17601
rect 31972 17561 31984 17595
rect 32018 17592 32030 17595
rect 33413 17595 33471 17601
rect 33413 17592 33425 17595
rect 32018 17564 33425 17592
rect 32018 17561 32030 17564
rect 31972 17555 32030 17561
rect 33413 17561 33425 17564
rect 33459 17561 33471 17595
rect 33413 17555 33471 17561
rect 25608 17496 26924 17524
rect 26973 17527 27031 17533
rect 26973 17493 26985 17527
rect 27019 17524 27031 17527
rect 27154 17524 27160 17536
rect 27019 17496 27160 17524
rect 27019 17493 27031 17496
rect 26973 17487 27031 17493
rect 27154 17484 27160 17496
rect 27212 17484 27218 17536
rect 27982 17524 27988 17536
rect 27943 17496 27988 17524
rect 27982 17484 27988 17496
rect 28040 17484 28046 17536
rect 29546 17524 29552 17536
rect 29507 17496 29552 17524
rect 29546 17484 29552 17496
rect 29604 17484 29610 17536
rect 30834 17524 30840 17536
rect 30795 17496 30840 17524
rect 30834 17484 30840 17496
rect 30892 17484 30898 17536
rect 32398 17484 32404 17536
rect 32456 17524 32462 17536
rect 33796 17524 33824 17623
rect 33870 17620 33876 17672
rect 33928 17660 33934 17672
rect 34057 17663 34115 17669
rect 33928 17632 33973 17660
rect 33928 17620 33934 17632
rect 34057 17629 34069 17663
rect 34103 17629 34115 17663
rect 34057 17623 34115 17629
rect 34072 17592 34100 17623
rect 34330 17620 34336 17672
rect 34388 17660 34394 17672
rect 34701 17663 34759 17669
rect 34701 17660 34713 17663
rect 34388 17632 34713 17660
rect 34388 17620 34394 17632
rect 34701 17629 34713 17632
rect 34747 17629 34759 17663
rect 35360 17660 35388 17759
rect 36173 17731 36231 17737
rect 36173 17697 36185 17731
rect 36219 17697 36231 17731
rect 36173 17691 36231 17697
rect 35897 17663 35955 17669
rect 35897 17660 35909 17663
rect 35360 17632 35909 17660
rect 34701 17623 34759 17629
rect 35897 17629 35909 17632
rect 35943 17629 35955 17663
rect 35897 17623 35955 17629
rect 35986 17592 35992 17604
rect 34072 17564 35992 17592
rect 35986 17552 35992 17564
rect 36044 17592 36050 17604
rect 36188 17592 36216 17691
rect 38473 17663 38531 17669
rect 38473 17660 38485 17663
rect 37660 17632 38485 17660
rect 36722 17592 36728 17604
rect 36044 17564 36728 17592
rect 36044 17552 36050 17564
rect 36722 17552 36728 17564
rect 36780 17552 36786 17604
rect 34790 17524 34796 17536
rect 32456 17496 34796 17524
rect 32456 17484 32462 17496
rect 34790 17484 34796 17496
rect 34848 17484 34854 17536
rect 35802 17484 35808 17536
rect 35860 17524 35866 17536
rect 37660 17533 37688 17632
rect 38473 17629 38485 17632
rect 38519 17629 38531 17663
rect 38473 17623 38531 17629
rect 38565 17663 38623 17669
rect 38565 17629 38577 17663
rect 38611 17629 38623 17663
rect 38565 17623 38623 17629
rect 37734 17552 37740 17604
rect 37792 17592 37798 17604
rect 38580 17592 38608 17623
rect 38654 17620 38660 17672
rect 38712 17660 38718 17672
rect 38712 17632 38757 17660
rect 38712 17620 38718 17632
rect 38838 17620 38844 17672
rect 38896 17660 38902 17672
rect 38896 17632 38941 17660
rect 38896 17620 38902 17632
rect 37792 17564 38608 17592
rect 37792 17552 37798 17564
rect 37645 17527 37703 17533
rect 37645 17524 37657 17527
rect 35860 17496 37657 17524
rect 35860 17484 35866 17496
rect 37645 17493 37657 17496
rect 37691 17493 37703 17527
rect 37645 17487 37703 17493
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 2314 17320 2320 17332
rect 2275 17292 2320 17320
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 6822 17320 6828 17332
rect 2832 17292 2877 17320
rect 6735 17292 6828 17320
rect 2832 17280 2838 17292
rect 6822 17280 6828 17292
rect 6880 17320 6886 17332
rect 7834 17320 7840 17332
rect 6880 17292 7840 17320
rect 6880 17280 6886 17292
rect 7834 17280 7840 17292
rect 7892 17320 7898 17332
rect 14553 17323 14611 17329
rect 7892 17292 12434 17320
rect 7892 17280 7898 17292
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 3850 17255 3908 17261
rect 3850 17252 3862 17255
rect 2648 17224 3862 17252
rect 2648 17212 2654 17224
rect 3850 17221 3862 17224
rect 3896 17221 3908 17255
rect 3850 17215 3908 17221
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 9738 17255 9796 17261
rect 9738 17252 9750 17255
rect 8168 17224 9750 17252
rect 8168 17212 8174 17224
rect 9738 17221 9750 17224
rect 9784 17221 9796 17255
rect 12406 17252 12434 17292
rect 14553 17289 14565 17323
rect 14599 17289 14611 17323
rect 14553 17283 14611 17289
rect 16025 17323 16083 17329
rect 16025 17289 16037 17323
rect 16071 17289 16083 17323
rect 19153 17323 19211 17329
rect 19153 17320 19165 17323
rect 16025 17283 16083 17289
rect 17052 17292 19165 17320
rect 12894 17252 12900 17264
rect 12406 17224 12900 17252
rect 9738 17215 9796 17221
rect 12894 17212 12900 17224
rect 12952 17212 12958 17264
rect 14568 17252 14596 17283
rect 15194 17252 15200 17264
rect 14568 17224 15200 17252
rect 15194 17212 15200 17224
rect 15252 17212 15258 17264
rect 15381 17255 15439 17261
rect 15381 17221 15393 17255
rect 15427 17252 15439 17255
rect 15470 17252 15476 17264
rect 15427 17224 15476 17252
rect 15427 17221 15439 17224
rect 15381 17215 15439 17221
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 16040 17252 16068 17283
rect 16850 17252 16856 17264
rect 16040 17224 16856 17252
rect 16850 17212 16856 17224
rect 16908 17212 16914 17264
rect 17052 17261 17080 17292
rect 19153 17289 19165 17292
rect 19199 17320 19211 17323
rect 24210 17320 24216 17332
rect 19199 17292 24216 17320
rect 19199 17289 19211 17292
rect 19153 17283 19211 17289
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 25866 17320 25872 17332
rect 24596 17292 25872 17320
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17221 17095 17255
rect 20070 17252 20076 17264
rect 17037 17215 17095 17221
rect 17880 17224 20076 17252
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1949 17187 2007 17193
rect 1949 17184 1961 17187
rect 1636 17156 1961 17184
rect 1636 17144 1642 17156
rect 1949 17153 1961 17156
rect 1995 17153 2007 17187
rect 1949 17147 2007 17153
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2682 17184 2688 17196
rect 2179 17156 2688 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 1964 17116 1992 17147
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 3050 17184 3056 17196
rect 3007 17156 3056 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17153 3203 17187
rect 3602 17184 3608 17196
rect 3563 17156 3608 17184
rect 3145 17147 3203 17153
rect 3160 17116 3188 17147
rect 3602 17144 3608 17156
rect 3660 17144 3666 17196
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 7282 17184 7288 17196
rect 4672 17156 7288 17184
rect 4672 17144 4678 17156
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 7466 17184 7472 17196
rect 7427 17156 7472 17184
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 7558 17144 7564 17196
rect 7616 17184 7622 17196
rect 7699 17187 7757 17193
rect 7616 17156 7661 17184
rect 7616 17144 7622 17156
rect 7699 17153 7711 17187
rect 7745 17184 7757 17187
rect 7834 17184 7840 17196
rect 7745 17156 7840 17184
rect 7745 17153 7757 17156
rect 7699 17147 7757 17153
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 9582 17184 9588 17196
rect 9539 17156 9588 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 13170 17184 13176 17196
rect 13131 17156 13176 17184
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 13262 17144 13268 17196
rect 13320 17184 13326 17196
rect 13429 17187 13487 17193
rect 13429 17184 13441 17187
rect 13320 17156 13441 17184
rect 13320 17144 13326 17156
rect 13429 17153 13441 17156
rect 13475 17153 13487 17187
rect 15488 17184 15516 17212
rect 15841 17187 15899 17193
rect 15841 17184 15853 17187
rect 15488 17156 15853 17184
rect 13429 17147 13487 17153
rect 15841 17153 15853 17156
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17368 17156 17785 17184
rect 17368 17144 17374 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17773 17147 17831 17153
rect 3510 17116 3516 17128
rect 1964 17088 3516 17116
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 17880 17116 17908 17224
rect 20070 17212 20076 17224
rect 20128 17252 20134 17264
rect 20346 17252 20352 17264
rect 20128 17224 20352 17252
rect 20128 17212 20134 17224
rect 20346 17212 20352 17224
rect 20404 17212 20410 17264
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 20993 17255 21051 17261
rect 20993 17252 21005 17255
rect 20864 17224 21005 17252
rect 20864 17212 20870 17224
rect 20993 17221 21005 17224
rect 21039 17221 21051 17255
rect 20993 17215 21051 17221
rect 21174 17212 21180 17264
rect 21232 17252 21238 17264
rect 24596 17252 24624 17292
rect 25866 17280 25872 17292
rect 25924 17280 25930 17332
rect 25958 17280 25964 17332
rect 26016 17320 26022 17332
rect 26053 17323 26111 17329
rect 26053 17320 26065 17323
rect 26016 17292 26065 17320
rect 26016 17280 26022 17292
rect 26053 17289 26065 17292
rect 26099 17289 26111 17323
rect 29641 17323 29699 17329
rect 29641 17320 29653 17323
rect 26053 17283 26111 17289
rect 27356 17292 29653 17320
rect 21232 17224 24624 17252
rect 21232 17212 21238 17224
rect 24670 17212 24676 17264
rect 24728 17252 24734 17264
rect 27356 17252 27384 17292
rect 29641 17289 29653 17292
rect 29687 17289 29699 17323
rect 32306 17320 32312 17332
rect 29641 17283 29699 17289
rect 29932 17292 32312 17320
rect 24728 17224 27384 17252
rect 24728 17212 24734 17224
rect 27614 17212 27620 17264
rect 27672 17252 27678 17264
rect 29932 17261 29960 17292
rect 32306 17280 32312 17292
rect 32364 17280 32370 17332
rect 32398 17280 32404 17332
rect 32456 17320 32462 17332
rect 33229 17323 33287 17329
rect 32456 17292 32501 17320
rect 32456 17280 32462 17292
rect 33229 17289 33241 17323
rect 33275 17320 33287 17323
rect 33870 17320 33876 17332
rect 33275 17292 33876 17320
rect 33275 17289 33287 17292
rect 33229 17283 33287 17289
rect 33870 17280 33876 17292
rect 33928 17280 33934 17332
rect 38654 17280 38660 17332
rect 38712 17320 38718 17332
rect 38841 17323 38899 17329
rect 38841 17320 38853 17323
rect 38712 17292 38853 17320
rect 38712 17280 38718 17292
rect 38841 17289 38853 17292
rect 38887 17289 38899 17323
rect 38841 17283 38899 17289
rect 29917 17255 29975 17261
rect 27672 17224 28672 17252
rect 27672 17212 27678 17224
rect 18046 17193 18052 17196
rect 18040 17147 18052 17193
rect 18104 17184 18110 17196
rect 19978 17184 19984 17196
rect 18104 17156 18140 17184
rect 19939 17156 19984 17184
rect 18046 17144 18052 17147
rect 18104 17144 18110 17156
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17153 20775 17187
rect 20898 17184 20904 17196
rect 20859 17156 20904 17184
rect 20717 17147 20775 17153
rect 14424 17088 17908 17116
rect 20732 17116 20760 17147
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17184 21143 17187
rect 22002 17184 22008 17196
rect 21131 17156 22008 17184
rect 21131 17153 21143 17156
rect 21085 17147 21143 17153
rect 22002 17144 22008 17156
rect 22060 17144 22066 17196
rect 22186 17184 22192 17196
rect 22147 17156 22192 17184
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 25869 17187 25927 17193
rect 25869 17184 25881 17187
rect 25240 17156 25881 17184
rect 21542 17116 21548 17128
rect 20732 17088 21548 17116
rect 14424 17076 14430 17088
rect 21542 17076 21548 17088
rect 21600 17076 21606 17128
rect 24946 17116 24952 17128
rect 24907 17088 24952 17116
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 25130 17076 25136 17128
rect 25188 17116 25194 17128
rect 25240 17125 25268 17156
rect 25869 17153 25881 17156
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 27798 17144 27804 17196
rect 27856 17184 27862 17196
rect 28644 17193 28672 17224
rect 29917 17221 29929 17255
rect 29963 17221 29975 17255
rect 29917 17215 29975 17221
rect 30834 17212 30840 17264
rect 30892 17252 30898 17264
rect 33045 17255 33103 17261
rect 33045 17252 33057 17255
rect 30892 17224 33057 17252
rect 30892 17212 30898 17224
rect 33045 17221 33057 17224
rect 33091 17221 33103 17255
rect 35710 17252 35716 17264
rect 33045 17215 33103 17221
rect 35084 17224 35716 17252
rect 28362 17187 28420 17193
rect 28362 17184 28374 17187
rect 27856 17156 28374 17184
rect 27856 17144 27862 17156
rect 28362 17153 28374 17156
rect 28408 17153 28420 17187
rect 28362 17147 28420 17153
rect 28629 17187 28687 17193
rect 28629 17153 28641 17187
rect 28675 17153 28687 17187
rect 29822 17184 29828 17196
rect 29783 17156 29828 17184
rect 28629 17147 28687 17153
rect 29822 17144 29828 17156
rect 29880 17144 29886 17196
rect 30009 17187 30067 17193
rect 30009 17153 30021 17187
rect 30055 17153 30067 17187
rect 30190 17184 30196 17196
rect 30151 17156 30196 17184
rect 30009 17147 30067 17153
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 25188 17088 25237 17116
rect 25188 17076 25194 17088
rect 25225 17085 25237 17088
rect 25271 17085 25283 17119
rect 25225 17079 25283 17085
rect 25685 17119 25743 17125
rect 25685 17085 25697 17119
rect 25731 17116 25743 17119
rect 26234 17116 26240 17128
rect 25731 17088 26240 17116
rect 25731 17085 25743 17088
rect 25685 17079 25743 17085
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 29914 17076 29920 17128
rect 29972 17116 29978 17128
rect 30024 17116 30052 17147
rect 30190 17144 30196 17156
rect 30248 17144 30254 17196
rect 32030 17184 32036 17196
rect 31312 17156 32036 17184
rect 29972 17088 30052 17116
rect 29972 17076 29978 17088
rect 15746 17008 15752 17060
rect 15804 17048 15810 17060
rect 21634 17048 21640 17060
rect 15804 17020 17632 17048
rect 15804 17008 15810 17020
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 3108 16952 4997 16980
rect 3108 16940 3114 16952
rect 4985 16949 4997 16952
rect 5031 16980 5043 16983
rect 7834 16980 7840 16992
rect 5031 16952 7840 16980
rect 5031 16949 5043 16952
rect 4985 16943 5043 16949
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 7929 16983 7987 16989
rect 7929 16949 7941 16983
rect 7975 16980 7987 16983
rect 8018 16980 8024 16992
rect 7975 16952 8024 16980
rect 7975 16949 7987 16952
rect 7929 16943 7987 16949
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8389 16983 8447 16989
rect 8389 16980 8401 16983
rect 8352 16952 8401 16980
rect 8352 16940 8358 16952
rect 8389 16949 8401 16952
rect 8435 16949 8447 16983
rect 8389 16943 8447 16949
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 10873 16983 10931 16989
rect 10873 16980 10885 16983
rect 9456 16952 10885 16980
rect 9456 16940 9462 16952
rect 10873 16949 10885 16952
rect 10919 16980 10931 16983
rect 11882 16980 11888 16992
rect 10919 16952 11888 16980
rect 10919 16949 10931 16952
rect 10873 16943 10931 16949
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 15013 16983 15071 16989
rect 15013 16980 15025 16983
rect 14700 16952 15025 16980
rect 14700 16940 14706 16952
rect 15013 16949 15025 16952
rect 15059 16949 15071 16983
rect 15013 16943 15071 16949
rect 17221 16983 17279 16989
rect 17221 16949 17233 16983
rect 17267 16980 17279 16983
rect 17494 16980 17500 16992
rect 17267 16952 17500 16980
rect 17267 16949 17279 16952
rect 17221 16943 17279 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 17604 16980 17632 17020
rect 18708 17020 21640 17048
rect 18708 16980 18736 17020
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 25774 17008 25780 17060
rect 25832 17048 25838 17060
rect 26786 17048 26792 17060
rect 25832 17020 26792 17048
rect 25832 17008 25838 17020
rect 26786 17008 26792 17020
rect 26844 17048 26850 17060
rect 27249 17051 27307 17057
rect 27249 17048 27261 17051
rect 26844 17020 27261 17048
rect 26844 17008 26850 17020
rect 27249 17017 27261 17020
rect 27295 17017 27307 17051
rect 31312 17048 31340 17156
rect 32030 17144 32036 17156
rect 32088 17144 32094 17196
rect 32214 17184 32220 17196
rect 32175 17156 32220 17184
rect 32214 17144 32220 17156
rect 32272 17144 32278 17196
rect 32392 17187 32450 17193
rect 32392 17184 32404 17187
rect 32324 17156 32404 17184
rect 32324 17128 32352 17156
rect 32392 17153 32404 17156
rect 32438 17153 32450 17187
rect 32858 17184 32864 17196
rect 32819 17156 32864 17184
rect 32392 17147 32450 17153
rect 32858 17144 32864 17156
rect 32916 17184 32922 17196
rect 34330 17184 34336 17196
rect 32916 17156 34336 17184
rect 32916 17144 32922 17156
rect 34330 17144 34336 17156
rect 34388 17144 34394 17196
rect 34790 17184 34796 17196
rect 34751 17156 34796 17184
rect 34790 17144 34796 17156
rect 34848 17144 34854 17196
rect 35084 17193 35112 17224
rect 35710 17212 35716 17224
rect 35768 17252 35774 17264
rect 37734 17252 37740 17264
rect 35768 17224 37740 17252
rect 35768 17212 35774 17224
rect 36464 17193 36492 17224
rect 37734 17212 37740 17224
rect 37792 17212 37798 17264
rect 35069 17187 35127 17193
rect 35069 17153 35081 17187
rect 35115 17153 35127 17187
rect 35069 17147 35127 17153
rect 36357 17187 36415 17193
rect 36357 17153 36369 17187
rect 36403 17153 36415 17187
rect 36357 17147 36415 17153
rect 36449 17187 36507 17193
rect 36449 17153 36461 17187
rect 36495 17153 36507 17187
rect 36449 17147 36507 17153
rect 32306 17116 32312 17128
rect 27249 17011 27307 17017
rect 29012 17020 31340 17048
rect 31956 17088 32312 17116
rect 17604 16952 18736 16980
rect 20165 16983 20223 16989
rect 20165 16949 20177 16983
rect 20211 16980 20223 16983
rect 21174 16980 21180 16992
rect 20211 16952 21180 16980
rect 20211 16949 20223 16952
rect 20165 16943 20223 16949
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 22370 16980 22376 16992
rect 21315 16952 22376 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 23382 16940 23388 16992
rect 23440 16980 23446 16992
rect 23477 16983 23535 16989
rect 23477 16980 23489 16983
rect 23440 16952 23489 16980
rect 23440 16940 23446 16952
rect 23477 16949 23489 16952
rect 23523 16949 23535 16983
rect 23477 16943 23535 16949
rect 27338 16940 27344 16992
rect 27396 16980 27402 16992
rect 29012 16980 29040 17020
rect 29178 16980 29184 16992
rect 27396 16952 29040 16980
rect 29139 16952 29184 16980
rect 27396 16940 27402 16952
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 29546 16940 29552 16992
rect 29604 16980 29610 16992
rect 31481 16983 31539 16989
rect 31481 16980 31493 16983
rect 29604 16952 31493 16980
rect 29604 16940 29610 16952
rect 31481 16949 31493 16952
rect 31527 16980 31539 16983
rect 31956 16980 31984 17088
rect 32306 17076 32312 17088
rect 32364 17076 32370 17128
rect 32030 17008 32036 17060
rect 32088 17048 32094 17060
rect 36372 17048 36400 17147
rect 36538 17144 36544 17196
rect 36596 17184 36602 17196
rect 36596 17156 36641 17184
rect 36596 17144 36602 17156
rect 36722 17144 36728 17196
rect 36780 17184 36786 17196
rect 38470 17184 38476 17196
rect 36780 17156 36825 17184
rect 38431 17156 38476 17184
rect 36780 17144 36786 17156
rect 38470 17144 38476 17156
rect 38528 17144 38534 17196
rect 38654 17184 38660 17196
rect 38615 17156 38660 17184
rect 38654 17144 38660 17156
rect 38712 17144 38718 17196
rect 37277 17051 37335 17057
rect 37277 17048 37289 17051
rect 32088 17020 37289 17048
rect 32088 17008 32094 17020
rect 37277 17017 37289 17020
rect 37323 17017 37335 17051
rect 67634 17048 67640 17060
rect 67595 17020 67640 17048
rect 37277 17011 37335 17017
rect 67634 17008 67640 17020
rect 67692 17008 67698 17060
rect 34146 16980 34152 16992
rect 31527 16952 31984 16980
rect 34107 16952 34152 16980
rect 31527 16949 31539 16952
rect 31481 16943 31539 16949
rect 34146 16940 34152 16952
rect 34204 16940 34210 16992
rect 36081 16983 36139 16989
rect 36081 16949 36093 16983
rect 36127 16980 36139 16983
rect 36170 16980 36176 16992
rect 36127 16952 36176 16980
rect 36127 16949 36139 16952
rect 36081 16943 36139 16949
rect 36170 16940 36176 16952
rect 36228 16940 36234 16992
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 2608 16748 2774 16776
rect 2038 16600 2044 16652
rect 2096 16640 2102 16652
rect 2608 16649 2636 16748
rect 2746 16708 2774 16748
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 8110 16776 8116 16788
rect 3384 16748 8116 16776
rect 3384 16736 3390 16748
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 11698 16776 11704 16788
rect 10100 16748 11704 16776
rect 10100 16736 10106 16748
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 12805 16779 12863 16785
rect 12805 16745 12817 16779
rect 12851 16776 12863 16779
rect 13262 16776 13268 16788
rect 12851 16748 13268 16776
rect 12851 16745 12863 16748
rect 12805 16739 12863 16745
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 14826 16736 14832 16788
rect 14884 16776 14890 16788
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 14884 16748 15485 16776
rect 14884 16736 14890 16748
rect 15473 16745 15485 16748
rect 15519 16745 15531 16779
rect 15473 16739 15531 16745
rect 2866 16708 2872 16720
rect 2746 16680 2872 16708
rect 2866 16668 2872 16680
rect 2924 16708 2930 16720
rect 3053 16711 3111 16717
rect 3053 16708 3065 16711
rect 2924 16680 3065 16708
rect 2924 16668 2930 16680
rect 3053 16677 3065 16680
rect 3099 16708 3111 16711
rect 3142 16708 3148 16720
rect 3099 16680 3148 16708
rect 3099 16677 3111 16680
rect 3053 16671 3111 16677
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 3234 16668 3240 16720
rect 3292 16708 3298 16720
rect 5350 16708 5356 16720
rect 3292 16680 5356 16708
rect 3292 16668 3298 16680
rect 5350 16668 5356 16680
rect 5408 16708 5414 16720
rect 7653 16711 7711 16717
rect 7653 16708 7665 16711
rect 5408 16680 7665 16708
rect 5408 16668 5414 16680
rect 7653 16677 7665 16680
rect 7699 16708 7711 16711
rect 9122 16708 9128 16720
rect 7699 16680 9128 16708
rect 7699 16677 7711 16680
rect 7653 16671 7711 16677
rect 9122 16668 9128 16680
rect 9180 16668 9186 16720
rect 10318 16708 10324 16720
rect 9508 16680 10324 16708
rect 2317 16643 2375 16649
rect 2317 16640 2329 16643
rect 2096 16612 2329 16640
rect 2096 16600 2102 16612
rect 2317 16609 2329 16612
rect 2363 16609 2375 16643
rect 2317 16603 2375 16609
rect 2593 16643 2651 16649
rect 2593 16609 2605 16643
rect 2639 16609 2651 16643
rect 9398 16640 9404 16652
rect 2593 16603 2651 16609
rect 4264 16612 9404 16640
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 3568 16544 3801 16572
rect 3568 16532 3574 16544
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 3789 16535 3847 16541
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16572 4031 16575
rect 4264 16572 4292 16612
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9508 16649 9536 16680
rect 10318 16668 10324 16680
rect 10376 16668 10382 16720
rect 13446 16668 13452 16720
rect 13504 16708 13510 16720
rect 14369 16711 14427 16717
rect 14369 16708 14381 16711
rect 13504 16680 14381 16708
rect 13504 16668 13510 16680
rect 14369 16677 14381 16680
rect 14415 16677 14427 16711
rect 15488 16708 15516 16739
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 16623 16779 16681 16785
rect 16623 16776 16635 16779
rect 15620 16748 16635 16776
rect 15620 16736 15626 16748
rect 16623 16745 16635 16748
rect 16669 16745 16681 16779
rect 16623 16739 16681 16745
rect 17957 16779 18015 16785
rect 17957 16745 17969 16779
rect 18003 16776 18015 16779
rect 18046 16776 18052 16788
rect 18003 16748 18052 16776
rect 18003 16745 18015 16748
rect 17957 16739 18015 16745
rect 18046 16736 18052 16748
rect 18104 16736 18110 16788
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 21729 16779 21787 16785
rect 21729 16776 21741 16779
rect 18196 16748 21741 16776
rect 18196 16736 18202 16748
rect 21729 16745 21741 16748
rect 21775 16745 21787 16779
rect 21729 16739 21787 16745
rect 22066 16748 23244 16776
rect 17678 16708 17684 16720
rect 15488 16680 17684 16708
rect 14369 16671 14427 16677
rect 17678 16668 17684 16680
rect 17736 16668 17742 16720
rect 18693 16711 18751 16717
rect 18693 16677 18705 16711
rect 18739 16708 18751 16711
rect 19426 16708 19432 16720
rect 18739 16680 19432 16708
rect 18739 16677 18751 16680
rect 18693 16671 18751 16677
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 22066 16708 22094 16748
rect 23014 16708 23020 16720
rect 19812 16680 22094 16708
rect 22664 16680 23020 16708
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 9732 16612 10977 16640
rect 9732 16600 9738 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 12710 16600 12716 16652
rect 12768 16640 12774 16652
rect 12768 16612 13216 16640
rect 12768 16600 12774 16612
rect 8110 16572 8116 16584
rect 4019 16544 4292 16572
rect 8071 16544 8116 16572
rect 4019 16541 4031 16544
rect 3973 16535 4031 16541
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 9766 16572 9772 16584
rect 9727 16544 9772 16572
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10594 16572 10600 16584
rect 10367 16544 10600 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 13188 16581 13216 16612
rect 13556 16612 16712 16640
rect 13556 16584 13584 16612
rect 13081 16575 13139 16581
rect 13081 16572 13093 16575
rect 12860 16544 13093 16572
rect 12860 16532 12866 16544
rect 13081 16541 13093 16544
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16541 13231 16575
rect 13173 16535 13231 16541
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13538 16572 13544 16584
rect 13495 16544 13544 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 6917 16507 6975 16513
rect 6917 16473 6929 16507
rect 6963 16504 6975 16507
rect 7374 16504 7380 16516
rect 6963 16476 7380 16504
rect 6963 16473 6975 16476
rect 6917 16467 6975 16473
rect 7374 16464 7380 16476
rect 7432 16504 7438 16516
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 7432 16476 7481 16504
rect 7432 16464 7438 16476
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 7469 16467 7527 16473
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11210 16507 11268 16513
rect 11210 16504 11222 16507
rect 11020 16476 11222 16504
rect 11020 16464 11026 16476
rect 11210 16473 11222 16476
rect 11256 16473 11268 16507
rect 13280 16504 13308 16535
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 16684 16572 16712 16612
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 19812 16649 19840 16680
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16816 16612 16865 16640
rect 16816 16600 16822 16612
rect 16853 16609 16865 16612
rect 16899 16640 16911 16643
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 16899 16612 19809 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 21542 16640 21548 16652
rect 20588 16612 21548 16640
rect 20588 16600 20594 16612
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 22664 16640 22692 16680
rect 23014 16668 23020 16680
rect 23072 16708 23078 16720
rect 23072 16680 23152 16708
rect 23072 16668 23078 16680
rect 23124 16649 23152 16680
rect 22066 16612 22692 16640
rect 23109 16643 23167 16649
rect 16942 16572 16948 16584
rect 16684 16544 16948 16572
rect 16942 16532 16948 16544
rect 17000 16572 17006 16584
rect 17313 16575 17371 16581
rect 17313 16572 17325 16575
rect 17000 16544 17325 16572
rect 17000 16532 17006 16544
rect 17313 16541 17325 16544
rect 17359 16541 17371 16575
rect 17494 16572 17500 16584
rect 17455 16544 17500 16572
rect 17313 16535 17371 16541
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 14642 16504 14648 16516
rect 13280 16476 14648 16504
rect 11210 16467 11268 16473
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 17604 16504 17632 16535
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 17736 16544 17781 16572
rect 17736 16532 17742 16544
rect 19058 16532 19064 16584
rect 19116 16572 19122 16584
rect 19521 16575 19579 16581
rect 19521 16572 19533 16575
rect 19116 16544 19533 16572
rect 19116 16532 19122 16544
rect 19521 16541 19533 16544
rect 19567 16541 19579 16575
rect 19521 16535 19579 16541
rect 17770 16504 17776 16516
rect 17604 16476 17776 16504
rect 17770 16464 17776 16476
rect 17828 16464 17834 16516
rect 19536 16504 19564 16535
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20809 16575 20867 16581
rect 20809 16572 20821 16575
rect 20772 16544 20821 16572
rect 20772 16532 20778 16544
rect 20809 16541 20821 16544
rect 20855 16541 20867 16575
rect 20809 16535 20867 16541
rect 21908 16575 21966 16581
rect 21908 16541 21920 16575
rect 21954 16572 21966 16575
rect 22066 16572 22094 16612
rect 23109 16609 23121 16643
rect 23155 16609 23167 16643
rect 23216 16640 23244 16748
rect 23382 16736 23388 16788
rect 23440 16776 23446 16788
rect 23440 16748 27568 16776
rect 23440 16736 23446 16748
rect 27540 16708 27568 16748
rect 27614 16736 27620 16788
rect 27672 16776 27678 16788
rect 27709 16779 27767 16785
rect 27709 16776 27721 16779
rect 27672 16748 27721 16776
rect 27672 16736 27678 16748
rect 27709 16745 27721 16748
rect 27755 16745 27767 16779
rect 27709 16739 27767 16745
rect 27982 16736 27988 16788
rect 28040 16776 28046 16788
rect 32677 16779 32735 16785
rect 28040 16748 31754 16776
rect 28040 16736 28046 16748
rect 30374 16708 30380 16720
rect 27540 16680 30380 16708
rect 30374 16668 30380 16680
rect 30432 16668 30438 16720
rect 31726 16708 31754 16748
rect 32677 16745 32689 16779
rect 32723 16776 32735 16779
rect 32858 16776 32864 16788
rect 32723 16748 32864 16776
rect 32723 16745 32735 16748
rect 32677 16739 32735 16745
rect 32858 16736 32864 16748
rect 32916 16736 32922 16788
rect 35069 16779 35127 16785
rect 35069 16745 35081 16779
rect 35115 16776 35127 16779
rect 36538 16776 36544 16788
rect 35115 16748 36544 16776
rect 35115 16745 35127 16748
rect 35069 16739 35127 16745
rect 36538 16736 36544 16748
rect 36596 16736 36602 16788
rect 35802 16708 35808 16720
rect 31726 16680 35808 16708
rect 35802 16668 35808 16680
rect 35860 16668 35866 16720
rect 24578 16640 24584 16652
rect 23216 16612 24584 16640
rect 23109 16603 23167 16609
rect 24578 16600 24584 16612
rect 24636 16600 24642 16652
rect 25777 16643 25835 16649
rect 25777 16609 25789 16643
rect 25823 16640 25835 16643
rect 27522 16640 27528 16652
rect 25823 16612 27528 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 29822 16640 29828 16652
rect 29735 16612 29828 16640
rect 22278 16572 22284 16584
rect 21954 16544 22094 16572
rect 22239 16544 22284 16572
rect 21954 16541 21966 16544
rect 21908 16535 21966 16541
rect 22278 16532 22284 16544
rect 22336 16532 22342 16584
rect 22370 16532 22376 16584
rect 22428 16572 22434 16584
rect 22830 16572 22836 16584
rect 22428 16544 22473 16572
rect 22791 16544 22836 16572
rect 22428 16532 22434 16544
rect 22830 16532 22836 16544
rect 22888 16532 22894 16584
rect 24946 16532 24952 16584
rect 25004 16572 25010 16584
rect 26237 16575 26295 16581
rect 26237 16572 26249 16575
rect 25004 16544 26249 16572
rect 25004 16532 25010 16544
rect 26237 16541 26249 16544
rect 26283 16541 26295 16575
rect 26418 16572 26424 16584
rect 26379 16544 26424 16572
rect 26237 16535 26295 16541
rect 26418 16532 26424 16544
rect 26476 16572 26482 16584
rect 29546 16572 29552 16584
rect 26476 16544 29552 16572
rect 26476 16532 26482 16544
rect 29546 16532 29552 16544
rect 29604 16532 29610 16584
rect 29748 16581 29776 16612
rect 29822 16600 29828 16612
rect 29880 16640 29886 16652
rect 31021 16643 31079 16649
rect 31021 16640 31033 16643
rect 29880 16612 31033 16640
rect 29880 16600 29886 16612
rect 31021 16609 31033 16612
rect 31067 16640 31079 16643
rect 32214 16640 32220 16652
rect 31067 16612 32220 16640
rect 31067 16609 31079 16612
rect 31021 16603 31079 16609
rect 32214 16600 32220 16612
rect 32272 16640 32278 16652
rect 35894 16640 35900 16652
rect 32272 16612 32536 16640
rect 35855 16612 35900 16640
rect 32272 16600 32278 16612
rect 29733 16575 29791 16581
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29914 16572 29920 16584
rect 29875 16544 29920 16572
rect 29733 16535 29791 16541
rect 29914 16532 29920 16544
rect 29972 16532 29978 16584
rect 30006 16532 30012 16584
rect 30064 16572 30070 16584
rect 30101 16575 30159 16581
rect 30101 16572 30113 16575
rect 30064 16544 30113 16572
rect 30064 16532 30070 16544
rect 30101 16541 30113 16544
rect 30147 16541 30159 16575
rect 30101 16535 30159 16541
rect 30745 16575 30803 16581
rect 30745 16541 30757 16575
rect 30791 16572 30803 16575
rect 30926 16572 30932 16584
rect 30791 16544 30932 16572
rect 30791 16541 30803 16544
rect 30745 16535 30803 16541
rect 30926 16532 30932 16544
rect 30984 16532 30990 16584
rect 32306 16572 32312 16584
rect 32267 16544 32312 16572
rect 32306 16532 32312 16544
rect 32364 16532 32370 16584
rect 32508 16581 32536 16612
rect 35894 16600 35900 16612
rect 35952 16600 35958 16652
rect 32493 16575 32551 16581
rect 32493 16541 32505 16575
rect 32539 16541 32551 16575
rect 32493 16535 32551 16541
rect 34146 16532 34152 16584
rect 34204 16572 34210 16584
rect 36170 16581 36176 16584
rect 34701 16575 34759 16581
rect 34701 16572 34713 16575
rect 34204 16544 34713 16572
rect 34204 16532 34210 16544
rect 34701 16541 34713 16544
rect 34747 16572 34759 16575
rect 36164 16572 36176 16581
rect 34747 16544 35940 16572
rect 36131 16544 36176 16572
rect 34747 16541 34759 16544
rect 34701 16535 34759 16541
rect 21634 16504 21640 16516
rect 19536 16476 21640 16504
rect 21634 16464 21640 16476
rect 21692 16464 21698 16516
rect 22005 16507 22063 16513
rect 22005 16473 22017 16507
rect 22051 16473 22063 16507
rect 22005 16467 22063 16473
rect 22097 16507 22155 16513
rect 22097 16473 22109 16507
rect 22143 16504 22155 16507
rect 22738 16504 22744 16516
rect 22143 16476 22744 16504
rect 22143 16473 22155 16476
rect 22097 16467 22155 16473
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 4157 16439 4215 16445
rect 4157 16436 4169 16439
rect 2832 16408 4169 16436
rect 2832 16396 2838 16408
rect 4157 16405 4169 16408
rect 4203 16405 4215 16439
rect 8294 16436 8300 16448
rect 8255 16408 8300 16436
rect 4157 16399 4215 16405
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 11606 16396 11612 16448
rect 11664 16436 11670 16448
rect 12345 16439 12403 16445
rect 12345 16436 12357 16439
rect 11664 16408 12357 16436
rect 11664 16396 11670 16408
rect 12345 16405 12357 16408
rect 12391 16405 12403 16439
rect 12345 16399 12403 16405
rect 18966 16396 18972 16448
rect 19024 16436 19030 16448
rect 20714 16436 20720 16448
rect 19024 16408 20720 16436
rect 19024 16396 19030 16408
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 20990 16436 20996 16448
rect 20951 16408 20996 16436
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 22020 16436 22048 16467
rect 22738 16464 22744 16476
rect 22796 16464 22802 16516
rect 25532 16507 25590 16513
rect 25532 16473 25544 16507
rect 25578 16504 25590 16507
rect 28074 16504 28080 16516
rect 25578 16476 28080 16504
rect 25578 16473 25590 16476
rect 25532 16467 25590 16473
rect 28074 16464 28080 16476
rect 28132 16464 28138 16516
rect 28997 16507 29055 16513
rect 28997 16473 29009 16507
rect 29043 16504 29055 16507
rect 29178 16504 29184 16516
rect 29043 16476 29184 16504
rect 29043 16473 29055 16476
rect 28997 16467 29055 16473
rect 29178 16464 29184 16476
rect 29236 16504 29242 16516
rect 29822 16504 29828 16516
rect 29236 16476 29684 16504
rect 29783 16476 29828 16504
rect 29236 16464 29242 16476
rect 24210 16436 24216 16448
rect 22020 16408 24216 16436
rect 24210 16396 24216 16408
rect 24268 16396 24274 16448
rect 24394 16436 24400 16448
rect 24355 16408 24400 16436
rect 24394 16396 24400 16408
rect 24452 16396 24458 16448
rect 26421 16439 26479 16445
rect 26421 16405 26433 16439
rect 26467 16436 26479 16439
rect 28442 16436 28448 16448
rect 26467 16408 28448 16436
rect 26467 16405 26479 16408
rect 26421 16399 26479 16405
rect 28442 16396 28448 16408
rect 28500 16396 28506 16448
rect 28534 16396 28540 16448
rect 28592 16436 28598 16448
rect 29549 16439 29607 16445
rect 29549 16436 29561 16439
rect 28592 16408 29561 16436
rect 28592 16396 28598 16408
rect 29549 16405 29561 16408
rect 29595 16405 29607 16439
rect 29656 16436 29684 16476
rect 29822 16464 29828 16476
rect 29880 16464 29886 16516
rect 32324 16504 32352 16532
rect 33137 16507 33195 16513
rect 33137 16504 33149 16507
rect 32324 16476 33149 16504
rect 33137 16473 33149 16476
rect 33183 16473 33195 16507
rect 33137 16467 33195 16473
rect 33226 16464 33232 16516
rect 33284 16504 33290 16516
rect 34885 16507 34943 16513
rect 34885 16504 34897 16507
rect 33284 16476 34897 16504
rect 33284 16464 33290 16476
rect 34885 16473 34897 16476
rect 34931 16473 34943 16507
rect 35912 16504 35940 16544
rect 36164 16535 36176 16544
rect 36170 16532 36176 16535
rect 36228 16532 36234 16584
rect 37642 16572 37648 16584
rect 36280 16544 37648 16572
rect 36280 16504 36308 16544
rect 37642 16532 37648 16544
rect 37700 16532 37706 16584
rect 39114 16572 39120 16584
rect 39075 16544 39120 16572
rect 39114 16532 39120 16544
rect 39172 16532 39178 16584
rect 35912 16476 36308 16504
rect 34885 16467 34943 16473
rect 30190 16436 30196 16448
rect 29656 16408 30196 16436
rect 29549 16399 29607 16405
rect 30190 16396 30196 16408
rect 30248 16396 30254 16448
rect 33962 16436 33968 16448
rect 33923 16408 33968 16436
rect 33962 16396 33968 16408
rect 34020 16396 34026 16448
rect 34900 16436 34928 16467
rect 36538 16464 36544 16516
rect 36596 16504 36602 16516
rect 38850 16507 38908 16513
rect 38850 16504 38862 16507
rect 36596 16476 38862 16504
rect 36596 16464 36602 16476
rect 38850 16473 38862 16476
rect 38896 16473 38908 16507
rect 38850 16467 38908 16473
rect 37277 16439 37335 16445
rect 37277 16436 37289 16439
rect 34900 16408 37289 16436
rect 37277 16405 37289 16408
rect 37323 16405 37335 16439
rect 37277 16399 37335 16405
rect 37458 16396 37464 16448
rect 37516 16436 37522 16448
rect 37737 16439 37795 16445
rect 37737 16436 37749 16439
rect 37516 16408 37749 16436
rect 37516 16396 37522 16408
rect 37737 16405 37749 16408
rect 37783 16405 37795 16439
rect 37737 16399 37795 16405
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3326 16232 3332 16244
rect 3283 16204 3332 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 7926 16232 7932 16244
rect 5224 16204 7932 16232
rect 5224 16192 5230 16204
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 9766 16232 9772 16244
rect 9727 16204 9772 16232
rect 9766 16192 9772 16204
rect 9824 16232 9830 16244
rect 10962 16232 10968 16244
rect 9824 16204 10732 16232
rect 10923 16204 10968 16232
rect 9824 16192 9830 16204
rect 3786 16164 3792 16176
rect 2976 16136 3792 16164
rect 2038 16056 2044 16108
rect 2096 16096 2102 16108
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 2096 16068 2605 16096
rect 2096 16056 2102 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2774 16096 2780 16108
rect 2735 16068 2780 16096
rect 2593 16059 2651 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 2976 16105 3004 16136
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 9674 16164 9680 16176
rect 7760 16136 9680 16164
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 2222 15988 2228 16040
rect 2280 16028 2286 16040
rect 2884 16028 2912 16059
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 4522 16096 4528 16108
rect 3752 16068 4528 16096
rect 3752 16056 3758 16068
rect 4522 16056 4528 16068
rect 4580 16056 4586 16108
rect 4704 16099 4762 16105
rect 4704 16065 4716 16099
rect 4750 16065 4762 16099
rect 4704 16059 4762 16065
rect 2280 16000 2912 16028
rect 4724 16028 4752 16059
rect 4801 16056 4807 16108
rect 4859 16096 4865 16108
rect 4939 16099 4997 16105
rect 4859 16068 4904 16096
rect 4859 16056 4865 16068
rect 4939 16065 4951 16099
rect 4985 16096 4997 16099
rect 5350 16096 5356 16108
rect 4985 16068 5356 16096
rect 4985 16065 4997 16068
rect 4939 16059 4997 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 6638 16096 6644 16108
rect 6599 16068 6644 16096
rect 6638 16056 6644 16068
rect 6696 16056 6702 16108
rect 6822 16096 6828 16108
rect 6783 16068 6828 16096
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7760 16105 7788 16136
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 8018 16105 8024 16108
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16065 7803 16099
rect 8012 16096 8024 16105
rect 7979 16068 8024 16096
rect 7745 16059 7803 16065
rect 8012 16059 8024 16068
rect 8018 16056 8024 16059
rect 8076 16056 8082 16108
rect 10318 16096 10324 16108
rect 10279 16068 10324 16096
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 10704 16105 10732 16204
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11388 16204 11897 16232
rect 11388 16192 11394 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 18417 16235 18475 16241
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 19242 16232 19248 16244
rect 18463 16204 19248 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10468 16068 10517 16096
rect 10468 16056 10474 16068
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 10689 16099 10747 16105
rect 10689 16065 10701 16099
rect 10735 16065 10747 16099
rect 10689 16059 10747 16065
rect 6457 16031 6515 16037
rect 6457 16028 6469 16031
rect 4724 16000 6469 16028
rect 2280 15988 2286 16000
rect 2608 15972 2636 16000
rect 6457 15997 6469 16000
rect 6503 15997 6515 16031
rect 10612 16028 10640 16059
rect 6457 15991 6515 15997
rect 10520 16000 10640 16028
rect 11900 16028 11928 16195
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 20898 16232 20904 16244
rect 19484 16204 20904 16232
rect 19484 16192 19490 16204
rect 12066 16124 12072 16176
rect 12124 16164 12130 16176
rect 12437 16167 12495 16173
rect 12437 16164 12449 16167
rect 12124 16136 12449 16164
rect 12124 16124 12130 16136
rect 12437 16133 12449 16136
rect 12483 16133 12495 16167
rect 15473 16167 15531 16173
rect 15473 16164 15485 16167
rect 12437 16127 12495 16133
rect 13740 16136 15485 16164
rect 12618 16096 12624 16108
rect 12579 16068 12624 16096
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 13538 16096 13544 16108
rect 13499 16068 13544 16096
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 13740 16105 13768 16136
rect 15473 16133 15485 16136
rect 15519 16133 15531 16167
rect 15473 16127 15531 16133
rect 15841 16167 15899 16173
rect 15841 16133 15853 16167
rect 15887 16164 15899 16167
rect 16666 16164 16672 16176
rect 15887 16136 16672 16164
rect 15887 16133 15899 16136
rect 15841 16127 15899 16133
rect 16666 16124 16672 16136
rect 16724 16164 16730 16176
rect 16850 16164 16856 16176
rect 16724 16136 16856 16164
rect 16724 16124 16730 16136
rect 16850 16124 16856 16136
rect 16908 16124 16914 16176
rect 19812 16173 19840 16204
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 21085 16235 21143 16241
rect 21085 16201 21097 16235
rect 21131 16232 21143 16235
rect 21818 16232 21824 16244
rect 21131 16204 21824 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 22830 16232 22836 16244
rect 21974 16204 22836 16232
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 17144 16136 19717 16164
rect 13704 16099 13768 16105
rect 13704 16065 13716 16099
rect 13750 16068 13768 16099
rect 13820 16099 13878 16105
rect 13750 16065 13762 16068
rect 13704 16059 13762 16065
rect 13820 16065 13832 16099
rect 13866 16065 13878 16099
rect 13820 16059 13878 16065
rect 11900 16000 12434 16028
rect 10520 15972 10548 16000
rect 2590 15920 2596 15972
rect 2648 15920 2654 15972
rect 10502 15920 10508 15972
rect 10560 15920 10566 15972
rect 12406 15960 12434 16000
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 13835 16028 13863 16059
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14642 16096 14648 16108
rect 13964 16068 14648 16096
rect 13964 16056 13970 16068
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 16114 16096 16120 16108
rect 15703 16068 16120 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 16114 16056 16120 16068
rect 16172 16096 16178 16108
rect 17144 16096 17172 16136
rect 19705 16133 19717 16136
rect 19751 16133 19763 16167
rect 19705 16127 19763 16133
rect 19797 16167 19855 16173
rect 19797 16133 19809 16167
rect 19843 16133 19855 16167
rect 21726 16164 21732 16176
rect 19797 16127 19855 16133
rect 19996 16136 21732 16164
rect 19996 16105 20024 16136
rect 21726 16124 21732 16136
rect 21784 16124 21790 16176
rect 16172 16068 17172 16096
rect 19613 16099 19671 16105
rect 16172 16056 16178 16068
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 13044 16000 13863 16028
rect 14185 16031 14243 16037
rect 13044 15988 13050 16000
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 14826 16028 14832 16040
rect 14231 16000 14832 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 16669 16031 16727 16037
rect 16669 15997 16681 16031
rect 16715 16028 16727 16031
rect 16758 16028 16764 16040
rect 16715 16000 16764 16028
rect 16715 15997 16727 16000
rect 16669 15991 16727 15997
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 16942 16028 16948 16040
rect 16903 16000 16948 16028
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 19628 16028 19656 16059
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21974 16105 22002 16204
rect 22830 16192 22836 16204
rect 22888 16232 22894 16244
rect 24213 16235 24271 16241
rect 24213 16232 24225 16235
rect 22888 16204 24225 16232
rect 22888 16192 22894 16204
rect 24213 16201 24225 16204
rect 24259 16232 24271 16235
rect 25130 16232 25136 16244
rect 24259 16204 25136 16232
rect 24259 16201 24271 16204
rect 24213 16195 24271 16201
rect 25130 16192 25136 16204
rect 25188 16192 25194 16244
rect 27617 16235 27675 16241
rect 27617 16201 27629 16235
rect 27663 16232 27675 16235
rect 27798 16232 27804 16244
rect 27663 16204 27804 16232
rect 27663 16201 27675 16204
rect 27617 16195 27675 16201
rect 27798 16192 27804 16204
rect 27856 16192 27862 16244
rect 28074 16232 28080 16244
rect 28035 16204 28080 16232
rect 28074 16192 28080 16204
rect 28132 16192 28138 16244
rect 28166 16192 28172 16244
rect 28224 16232 28230 16244
rect 33962 16232 33968 16244
rect 28224 16204 33968 16232
rect 28224 16192 28230 16204
rect 33962 16192 33968 16204
rect 34020 16232 34026 16244
rect 36538 16232 36544 16244
rect 34020 16204 34468 16232
rect 36499 16204 36544 16232
rect 34020 16192 34026 16204
rect 22097 16167 22155 16173
rect 22097 16133 22109 16167
rect 22143 16164 22155 16167
rect 24394 16164 24400 16176
rect 22143 16136 24400 16164
rect 22143 16133 22155 16136
rect 22097 16127 22155 16133
rect 24394 16124 24400 16136
rect 24452 16164 24458 16176
rect 25961 16167 26019 16173
rect 25961 16164 25973 16167
rect 24452 16136 25973 16164
rect 24452 16124 24458 16136
rect 25961 16133 25973 16136
rect 26007 16133 26019 16167
rect 27706 16164 27712 16176
rect 25961 16127 26019 16133
rect 27264 16136 27712 16164
rect 21177 16099 21235 16105
rect 21177 16096 21189 16099
rect 20956 16068 21189 16096
rect 20956 16056 20962 16068
rect 21177 16065 21189 16068
rect 21223 16065 21235 16099
rect 21177 16059 21235 16065
rect 21959 16099 22017 16105
rect 21959 16065 21971 16099
rect 22005 16065 22017 16099
rect 22186 16096 22192 16108
rect 22147 16068 22192 16096
rect 21959 16059 22017 16065
rect 20438 16028 20444 16040
rect 19628 16000 20444 16028
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 21082 15988 21088 16040
rect 21140 16028 21146 16040
rect 21974 16028 22002 16059
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22372 16099 22430 16105
rect 22372 16065 22384 16099
rect 22418 16065 22430 16099
rect 22372 16059 22430 16065
rect 21140 16000 22002 16028
rect 22388 16028 22416 16059
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 23014 16096 23020 16108
rect 22520 16068 22565 16096
rect 22927 16068 23020 16096
rect 22520 16056 22526 16068
rect 23014 16056 23020 16068
rect 23072 16096 23078 16108
rect 23474 16096 23480 16108
rect 23072 16068 23480 16096
rect 23072 16056 23078 16068
rect 23474 16056 23480 16068
rect 23532 16096 23538 16108
rect 23569 16099 23627 16105
rect 23569 16096 23581 16099
rect 23532 16068 23581 16096
rect 23532 16056 23538 16068
rect 23569 16065 23581 16068
rect 23615 16065 23627 16099
rect 23569 16059 23627 16065
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16096 25835 16099
rect 25866 16096 25872 16108
rect 25823 16068 25872 16096
rect 25823 16065 25835 16068
rect 25777 16059 25835 16065
rect 25866 16056 25872 16068
rect 25924 16056 25930 16108
rect 26970 16096 26976 16108
rect 26931 16068 26976 16096
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 27154 16096 27160 16108
rect 27115 16068 27160 16096
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27264 16105 27292 16136
rect 27706 16124 27712 16136
rect 27764 16124 27770 16176
rect 28626 16164 28632 16176
rect 28276 16136 28632 16164
rect 27252 16099 27310 16105
rect 27252 16065 27264 16099
rect 27298 16065 27310 16099
rect 27252 16059 27310 16065
rect 27338 16056 27344 16108
rect 27396 16096 27402 16108
rect 28276 16096 28304 16136
rect 28626 16124 28632 16136
rect 28684 16124 28690 16176
rect 30834 16124 30840 16176
rect 30892 16164 30898 16176
rect 31021 16167 31079 16173
rect 31021 16164 31033 16167
rect 30892 16136 31033 16164
rect 30892 16124 30898 16136
rect 31021 16133 31033 16136
rect 31067 16133 31079 16167
rect 31021 16127 31079 16133
rect 33444 16167 33502 16173
rect 33444 16133 33456 16167
rect 33490 16164 33502 16167
rect 34149 16167 34207 16173
rect 34149 16164 34161 16167
rect 33490 16136 34161 16164
rect 33490 16133 33502 16136
rect 33444 16127 33502 16133
rect 34149 16133 34161 16136
rect 34195 16133 34207 16167
rect 34149 16127 34207 16133
rect 28353 16099 28411 16105
rect 28353 16096 28365 16099
rect 27396 16068 27441 16096
rect 28276 16068 28365 16096
rect 27396 16056 27402 16068
rect 28353 16065 28365 16068
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 28445 16099 28503 16105
rect 28445 16065 28457 16099
rect 28491 16065 28503 16099
rect 28445 16059 28503 16065
rect 28537 16099 28595 16105
rect 28537 16065 28549 16099
rect 28583 16065 28595 16099
rect 28718 16096 28724 16108
rect 28679 16068 28724 16096
rect 28537 16059 28595 16065
rect 23842 16028 23848 16040
rect 22388 16000 23848 16028
rect 21140 15988 21146 16000
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 26145 16031 26203 16037
rect 26145 15997 26157 16031
rect 26191 15997 26203 16031
rect 26145 15991 26203 15997
rect 13722 15960 13728 15972
rect 12406 15932 13728 15960
rect 12406 15904 12434 15932
rect 13722 15920 13728 15932
rect 13780 15960 13786 15972
rect 15010 15960 15016 15972
rect 13780 15932 15016 15960
rect 13780 15920 13786 15932
rect 15010 15920 15016 15932
rect 15068 15920 15074 15972
rect 19610 15920 19616 15972
rect 19668 15960 19674 15972
rect 21821 15963 21879 15969
rect 21821 15960 21833 15963
rect 19668 15932 21833 15960
rect 19668 15920 19674 15932
rect 21821 15929 21833 15932
rect 21867 15929 21879 15963
rect 21821 15923 21879 15929
rect 22462 15920 22468 15972
rect 22520 15960 22526 15972
rect 23014 15960 23020 15972
rect 22520 15932 23020 15960
rect 22520 15920 22526 15932
rect 23014 15920 23020 15932
rect 23072 15920 23078 15972
rect 26160 15960 26188 15991
rect 28460 15972 28488 16059
rect 26160 15932 26924 15960
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5258 15892 5264 15904
rect 5215 15864 5264 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5442 15852 5448 15904
rect 5500 15892 5506 15904
rect 7374 15892 7380 15904
rect 5500 15864 7380 15892
rect 5500 15852 5506 15864
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8996 15864 9137 15892
rect 8996 15852 9002 15864
rect 9125 15861 9137 15864
rect 9171 15861 9183 15895
rect 12406 15864 12440 15904
rect 9125 15855 9183 15861
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 16206 15892 16212 15904
rect 14976 15864 16212 15892
rect 14976 15852 14982 15864
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 17586 15892 17592 15904
rect 16816 15864 17592 15892
rect 16816 15852 16822 15864
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 18966 15892 18972 15904
rect 18927 15864 18972 15892
rect 18966 15852 18972 15864
rect 19024 15852 19030 15904
rect 19429 15895 19487 15901
rect 19429 15861 19441 15895
rect 19475 15892 19487 15895
rect 20346 15892 20352 15904
rect 19475 15864 20352 15892
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 20346 15852 20352 15864
rect 20404 15852 20410 15904
rect 20530 15892 20536 15904
rect 20491 15864 20536 15892
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 23566 15852 23572 15904
rect 23624 15892 23630 15904
rect 23661 15895 23719 15901
rect 23661 15892 23673 15895
rect 23624 15864 23673 15892
rect 23624 15852 23630 15864
rect 23661 15861 23673 15864
rect 23707 15892 23719 15895
rect 25225 15895 25283 15901
rect 25225 15892 25237 15895
rect 23707 15864 25237 15892
rect 23707 15861 23719 15864
rect 23661 15855 23719 15861
rect 25225 15861 25237 15864
rect 25271 15892 25283 15895
rect 26418 15892 26424 15904
rect 25271 15864 26424 15892
rect 25271 15861 25283 15864
rect 25225 15855 25283 15861
rect 26418 15852 26424 15864
rect 26476 15852 26482 15904
rect 26896 15892 26924 15932
rect 28442 15920 28448 15972
rect 28500 15920 28506 15972
rect 28552 15892 28580 16059
rect 28718 16056 28724 16068
rect 28776 16056 28782 16108
rect 29914 16096 29920 16108
rect 29875 16068 29920 16096
rect 29914 16056 29920 16068
rect 29972 16056 29978 16108
rect 30926 16096 30932 16108
rect 30887 16068 30932 16096
rect 30926 16056 30932 16068
rect 30984 16056 30990 16108
rect 31113 16099 31171 16105
rect 31113 16065 31125 16099
rect 31159 16096 31171 16099
rect 31294 16096 31300 16108
rect 31159 16068 31193 16096
rect 31255 16068 31300 16096
rect 31159 16065 31171 16068
rect 31113 16059 31171 16065
rect 30193 16031 30251 16037
rect 30193 15997 30205 16031
rect 30239 16028 30251 16031
rect 31128 16028 31156 16059
rect 31294 16056 31300 16068
rect 31352 16056 31358 16108
rect 32674 16056 32680 16108
rect 32732 16096 32738 16108
rect 34440 16105 34468 16204
rect 36538 16192 36544 16204
rect 36596 16192 36602 16244
rect 37277 16167 37335 16173
rect 37277 16164 37289 16167
rect 36096 16136 37289 16164
rect 33689 16099 33747 16105
rect 33689 16096 33701 16099
rect 32732 16068 33701 16096
rect 32732 16056 32738 16068
rect 33689 16065 33701 16068
rect 33735 16065 33747 16099
rect 33689 16059 33747 16065
rect 34425 16099 34483 16105
rect 34425 16065 34437 16099
rect 34471 16065 34483 16099
rect 34425 16059 34483 16065
rect 34517 16099 34575 16105
rect 34517 16065 34529 16099
rect 34563 16065 34575 16099
rect 34517 16059 34575 16065
rect 31202 16028 31208 16040
rect 30239 16000 31208 16028
rect 30239 15997 30251 16000
rect 30193 15991 30251 15997
rect 31202 15988 31208 16000
rect 31260 15988 31266 16040
rect 34532 16028 34560 16059
rect 34606 16056 34612 16108
rect 34664 16096 34670 16108
rect 34793 16099 34851 16105
rect 34664 16068 34709 16096
rect 34664 16056 34670 16068
rect 34793 16065 34805 16099
rect 34839 16096 34851 16099
rect 35897 16099 35955 16105
rect 35897 16096 35909 16099
rect 34839 16068 35909 16096
rect 34839 16065 34851 16068
rect 34793 16059 34851 16065
rect 35897 16065 35909 16068
rect 35943 16096 35955 16099
rect 35986 16096 35992 16108
rect 35943 16068 35992 16096
rect 35943 16065 35955 16068
rect 35897 16059 35955 16065
rect 35986 16056 35992 16068
rect 36044 16056 36050 16108
rect 36096 16105 36124 16136
rect 37277 16133 37289 16136
rect 37323 16133 37335 16167
rect 37642 16164 37648 16176
rect 37555 16136 37648 16164
rect 37277 16127 37335 16133
rect 37642 16124 37648 16136
rect 37700 16164 37706 16176
rect 38470 16164 38476 16176
rect 37700 16136 38476 16164
rect 37700 16124 37706 16136
rect 38470 16124 38476 16136
rect 38528 16124 38534 16176
rect 36081 16099 36139 16105
rect 36081 16065 36093 16099
rect 36127 16065 36139 16099
rect 36081 16059 36139 16065
rect 36173 16099 36231 16105
rect 36173 16065 36185 16099
rect 36219 16065 36231 16099
rect 36173 16059 36231 16065
rect 36265 16099 36323 16105
rect 36265 16065 36277 16099
rect 36311 16065 36323 16099
rect 37458 16096 37464 16108
rect 37419 16068 37464 16096
rect 36265 16059 36323 16065
rect 35710 16028 35716 16040
rect 34532 16000 35716 16028
rect 35710 15988 35716 16000
rect 35768 16028 35774 16040
rect 36188 16028 36216 16059
rect 35768 16000 36216 16028
rect 35768 15988 35774 16000
rect 29086 15920 29092 15972
rect 29144 15960 29150 15972
rect 30282 15960 30288 15972
rect 29144 15932 30288 15960
rect 29144 15920 29150 15932
rect 30282 15920 30288 15932
rect 30340 15960 30346 15972
rect 36280 15960 36308 16059
rect 37458 16056 37464 16068
rect 37516 16056 37522 16108
rect 30340 15932 32812 15960
rect 30340 15920 30346 15932
rect 30742 15892 30748 15904
rect 26896 15864 28580 15892
rect 30703 15864 30748 15892
rect 30742 15852 30748 15864
rect 30800 15852 30806 15904
rect 32306 15892 32312 15904
rect 32267 15864 32312 15892
rect 32306 15852 32312 15864
rect 32364 15852 32370 15904
rect 32784 15892 32812 15932
rect 35360 15932 36308 15960
rect 35360 15901 35388 15932
rect 35345 15895 35403 15901
rect 35345 15892 35357 15895
rect 32784 15864 35357 15892
rect 35345 15861 35357 15864
rect 35391 15861 35403 15895
rect 67634 15892 67640 15904
rect 67595 15864 67640 15892
rect 35345 15855 35403 15861
rect 67634 15852 67640 15864
rect 67692 15852 67698 15904
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 2958 15688 2964 15700
rect 2919 15660 2964 15688
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 4525 15691 4583 15697
rect 4525 15657 4537 15691
rect 4571 15688 4583 15691
rect 5166 15688 5172 15700
rect 4571 15660 5172 15688
rect 4571 15657 4583 15660
rect 4525 15651 4583 15657
rect 4540 15552 4568 15651
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 6365 15691 6423 15697
rect 6365 15657 6377 15691
rect 6411 15688 6423 15691
rect 6638 15688 6644 15700
rect 6411 15660 6644 15688
rect 6411 15657 6423 15660
rect 6365 15651 6423 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 7650 15688 7656 15700
rect 7611 15660 7656 15688
rect 7650 15648 7656 15660
rect 7708 15648 7714 15700
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 7984 15660 8309 15688
rect 7984 15648 7990 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 8297 15651 8355 15657
rect 9398 15648 9404 15700
rect 9456 15688 9462 15700
rect 10873 15691 10931 15697
rect 10873 15688 10885 15691
rect 9456 15660 10885 15688
rect 9456 15648 9462 15660
rect 10873 15657 10885 15660
rect 10919 15688 10931 15691
rect 11330 15688 11336 15700
rect 10919 15660 11336 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 14182 15688 14188 15700
rect 14143 15660 14188 15688
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 15378 15688 15384 15700
rect 15339 15660 15384 15688
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 17236 15660 19334 15688
rect 2746 15524 4568 15552
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2317 15487 2375 15493
rect 2317 15484 2329 15487
rect 2096 15456 2329 15484
rect 2096 15444 2102 15456
rect 2317 15453 2329 15456
rect 2363 15453 2375 15487
rect 2317 15447 2375 15453
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 1489 15419 1547 15425
rect 1489 15385 1501 15419
rect 1535 15416 1547 15419
rect 1578 15416 1584 15428
rect 1535 15388 1584 15416
rect 1535 15385 1547 15388
rect 1489 15379 1547 15385
rect 1578 15376 1584 15388
rect 1636 15376 1642 15428
rect 1670 15376 1676 15428
rect 1728 15416 1734 15428
rect 1857 15419 1915 15425
rect 1728 15388 1773 15416
rect 1728 15376 1734 15388
rect 1857 15385 1869 15419
rect 1903 15416 1915 15419
rect 2516 15416 2544 15447
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 2746 15493 2774 15524
rect 2731 15487 2789 15493
rect 2648 15456 2693 15484
rect 2648 15444 2654 15456
rect 2731 15453 2743 15487
rect 2777 15453 2789 15487
rect 3786 15484 3792 15496
rect 3747 15456 3792 15484
rect 2731 15447 2789 15453
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4062 15444 4068 15496
rect 4120 15484 4126 15496
rect 5258 15493 5264 15496
rect 4985 15487 5043 15493
rect 4985 15484 4997 15487
rect 4120 15456 4997 15484
rect 4120 15444 4126 15456
rect 4985 15453 4997 15456
rect 5031 15453 5043 15487
rect 5252 15484 5264 15493
rect 5219 15456 5264 15484
rect 4985 15447 5043 15453
rect 5252 15447 5264 15456
rect 5258 15444 5264 15447
rect 5316 15444 5322 15496
rect 6656 15484 6684 15648
rect 9490 15620 9496 15632
rect 7484 15592 9352 15620
rect 9451 15592 9496 15620
rect 7006 15512 7012 15564
rect 7064 15552 7070 15564
rect 7484 15552 7512 15592
rect 7064 15524 7512 15552
rect 7064 15512 7070 15524
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 6656 15456 7113 15484
rect 7101 15453 7113 15456
rect 7147 15453 7159 15487
rect 7374 15484 7380 15496
rect 7335 15456 7380 15484
rect 7101 15447 7159 15453
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7484 15493 7512 15524
rect 7834 15512 7840 15564
rect 7892 15552 7898 15564
rect 7892 15524 9260 15552
rect 7892 15512 7898 15524
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 8018 15444 8024 15496
rect 8076 15484 8082 15496
rect 8938 15484 8944 15496
rect 8076 15456 8944 15484
rect 8076 15444 8082 15456
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9232 15493 9260 15524
rect 9324 15496 9352 15592
rect 9490 15580 9496 15592
rect 9548 15580 9554 15632
rect 17236 15620 17264 15660
rect 17770 15620 17776 15632
rect 15488 15592 17264 15620
rect 17328 15592 17776 15620
rect 15488 15561 15516 15592
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15521 15531 15555
rect 15473 15515 15531 15521
rect 17034 15512 17040 15564
rect 17092 15512 17098 15564
rect 17328 15552 17356 15592
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 19306 15620 19334 15660
rect 19702 15648 19708 15700
rect 19760 15688 19766 15700
rect 20162 15688 20168 15700
rect 19760 15660 20168 15688
rect 19760 15648 19766 15660
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 20254 15648 20260 15700
rect 20312 15648 20318 15700
rect 21450 15688 21456 15700
rect 21411 15660 21456 15688
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 22370 15688 22376 15700
rect 22331 15660 22376 15688
rect 22370 15648 22376 15660
rect 22428 15648 22434 15700
rect 22830 15648 22836 15700
rect 22888 15688 22894 15700
rect 23753 15691 23811 15697
rect 23753 15688 23765 15691
rect 22888 15660 23765 15688
rect 22888 15648 22894 15660
rect 23753 15657 23765 15660
rect 23799 15657 23811 15691
rect 23753 15651 23811 15657
rect 26329 15691 26387 15697
rect 26329 15657 26341 15691
rect 26375 15688 26387 15691
rect 27338 15688 27344 15700
rect 26375 15660 27344 15688
rect 26375 15657 26387 15660
rect 26329 15651 26387 15657
rect 27338 15648 27344 15660
rect 27396 15648 27402 15700
rect 33781 15691 33839 15697
rect 33781 15657 33793 15691
rect 33827 15688 33839 15691
rect 34606 15688 34612 15700
rect 33827 15660 34612 15688
rect 33827 15657 33839 15660
rect 33781 15651 33839 15657
rect 34606 15648 34612 15660
rect 34664 15648 34670 15700
rect 38654 15688 38660 15700
rect 35176 15660 38660 15688
rect 19978 15620 19984 15632
rect 19306 15592 19984 15620
rect 19978 15580 19984 15592
rect 20036 15580 20042 15632
rect 17236 15524 17356 15552
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 9306 15444 9312 15496
rect 9364 15484 9370 15496
rect 9364 15456 9457 15484
rect 9364 15444 9370 15456
rect 11790 15444 11796 15496
rect 11848 15484 11854 15496
rect 15565 15487 15623 15493
rect 11848 15456 15332 15484
rect 11848 15444 11854 15456
rect 1903 15388 2544 15416
rect 3804 15416 3832 15444
rect 7006 15416 7012 15428
rect 3804 15388 7012 15416
rect 1903 15385 1915 15388
rect 1857 15379 1915 15385
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 7282 15416 7288 15428
rect 7243 15388 7288 15416
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 7834 15376 7840 15428
rect 7892 15416 7898 15428
rect 8202 15416 8208 15428
rect 7892 15388 8208 15416
rect 7892 15376 7898 15388
rect 8202 15376 8208 15388
rect 8260 15376 8266 15428
rect 9122 15416 9128 15428
rect 9083 15388 9128 15416
rect 9122 15376 9128 15388
rect 9180 15376 9186 15428
rect 12161 15419 12219 15425
rect 12161 15385 12173 15419
rect 12207 15416 12219 15419
rect 13446 15416 13452 15428
rect 12207 15388 13452 15416
rect 12207 15385 12219 15388
rect 12161 15379 12219 15385
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 15304 15416 15332 15456
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 16758 15484 16764 15496
rect 15611 15456 16764 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 16758 15444 16764 15456
rect 16816 15444 16822 15496
rect 16942 15484 16948 15496
rect 16903 15456 16948 15484
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17052 15478 17080 15512
rect 17236 15493 17264 15524
rect 17586 15512 17592 15564
rect 17644 15552 17650 15564
rect 19610 15552 19616 15564
rect 17644 15524 19616 15552
rect 17644 15512 17650 15524
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 17129 15487 17187 15493
rect 17129 15478 17141 15487
rect 17052 15453 17141 15478
rect 17175 15453 17187 15487
rect 17052 15450 17187 15453
rect 17129 15447 17187 15450
rect 17224 15487 17282 15493
rect 17224 15453 17236 15487
rect 17270 15453 17282 15487
rect 17224 15447 17282 15453
rect 17333 15487 17391 15493
rect 17333 15453 17345 15487
rect 17379 15484 17391 15487
rect 17379 15481 17448 15484
rect 17379 15456 17540 15481
rect 17379 15453 17391 15456
rect 17420 15453 17540 15456
rect 17333 15447 17391 15453
rect 15470 15416 15476 15428
rect 15304 15388 15476 15416
rect 15470 15376 15476 15388
rect 15528 15416 15534 15428
rect 16393 15419 16451 15425
rect 16393 15416 16405 15419
rect 15528 15388 16405 15416
rect 15528 15376 15534 15388
rect 16393 15385 16405 15388
rect 16439 15416 16451 15419
rect 17512 15416 17540 15453
rect 17862 15444 17868 15496
rect 17920 15484 17926 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 17920 15456 18613 15484
rect 17920 15444 17926 15456
rect 18601 15453 18613 15456
rect 18647 15484 18659 15487
rect 19058 15484 19064 15496
rect 18647 15456 19064 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19334 15484 19340 15496
rect 19208 15456 19340 15484
rect 19208 15444 19214 15456
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 19702 15444 19708 15496
rect 19760 15484 19766 15496
rect 19843 15487 19901 15493
rect 19843 15484 19855 15487
rect 19760 15456 19855 15484
rect 19760 15444 19766 15456
rect 19843 15453 19855 15456
rect 19889 15453 19901 15487
rect 19843 15447 19901 15453
rect 19984 15487 20042 15493
rect 19984 15453 19996 15487
rect 20030 15481 20042 15487
rect 20162 15481 20168 15496
rect 20030 15453 20168 15481
rect 19984 15447 20042 15453
rect 20162 15444 20168 15453
rect 20220 15444 20226 15496
rect 20271 15493 20299 15648
rect 29546 15620 29552 15632
rect 26988 15592 29552 15620
rect 20438 15512 20444 15564
rect 20496 15552 20502 15564
rect 21450 15552 21456 15564
rect 20496 15524 21456 15552
rect 20496 15512 20502 15524
rect 21450 15512 21456 15524
rect 21508 15552 21514 15564
rect 22002 15552 22008 15564
rect 21508 15524 22008 15552
rect 21508 15512 21514 15524
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 24210 15512 24216 15564
rect 24268 15552 24274 15564
rect 26988 15552 27016 15592
rect 29546 15580 29552 15592
rect 29604 15580 29610 15632
rect 35176 15620 35204 15660
rect 38654 15648 38660 15660
rect 38712 15648 38718 15700
rect 35986 15620 35992 15632
rect 30116 15592 35204 15620
rect 35268 15592 35992 15620
rect 24268 15524 27016 15552
rect 24268 15512 24274 15524
rect 20256 15487 20314 15493
rect 20256 15453 20268 15487
rect 20302 15453 20314 15487
rect 20256 15447 20314 15453
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 20404 15456 20449 15484
rect 20404 15444 20410 15456
rect 21726 15444 21732 15496
rect 21784 15484 21790 15496
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 21784 15456 22293 15484
rect 21784 15444 21790 15456
rect 22281 15453 22293 15456
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 22373 15487 22431 15493
rect 22373 15453 22385 15487
rect 22419 15484 22431 15487
rect 22922 15484 22928 15496
rect 22419 15456 22928 15484
rect 22419 15453 22431 15456
rect 22373 15447 22431 15453
rect 22922 15444 22928 15456
rect 22980 15444 22986 15496
rect 23106 15484 23112 15496
rect 23067 15456 23112 15484
rect 23106 15444 23112 15456
rect 23164 15484 23170 15496
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 23164 15456 24409 15484
rect 23164 15444 23170 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 24397 15447 24455 15453
rect 26326 15444 26332 15496
rect 26384 15484 26390 15496
rect 26694 15484 26700 15496
rect 26384 15456 26700 15484
rect 26384 15444 26390 15456
rect 26694 15444 26700 15456
rect 26752 15484 26758 15496
rect 26988 15493 27016 15524
rect 27157 15555 27215 15561
rect 27157 15521 27169 15555
rect 27203 15552 27215 15555
rect 27203 15524 27844 15552
rect 27203 15521 27215 15524
rect 27157 15515 27215 15521
rect 26789 15487 26847 15493
rect 26789 15484 26801 15487
rect 26752 15456 26801 15484
rect 26752 15444 26758 15456
rect 26789 15453 26801 15456
rect 26835 15453 26847 15487
rect 26789 15447 26847 15453
rect 26973 15487 27031 15493
rect 26973 15453 26985 15487
rect 27019 15453 27031 15487
rect 26973 15447 27031 15453
rect 27062 15444 27068 15496
rect 27120 15484 27126 15496
rect 27816 15493 27844 15524
rect 27617 15487 27675 15493
rect 27617 15484 27629 15487
rect 27120 15456 27629 15484
rect 27120 15444 27126 15456
rect 27617 15453 27629 15456
rect 27663 15453 27675 15487
rect 27617 15447 27675 15453
rect 27801 15487 27859 15493
rect 27801 15453 27813 15487
rect 27847 15453 27859 15487
rect 27801 15447 27859 15453
rect 27893 15487 27951 15493
rect 27893 15453 27905 15487
rect 27939 15453 27951 15487
rect 27893 15447 27951 15453
rect 27985 15487 28043 15493
rect 27985 15453 27997 15487
rect 28031 15484 28043 15487
rect 28166 15484 28172 15496
rect 28031 15456 28172 15484
rect 28031 15453 28043 15456
rect 27985 15447 28043 15453
rect 16439 15388 17540 15416
rect 16439 15385 16451 15388
rect 16393 15379 16451 15385
rect 17678 15376 17684 15428
rect 17736 15416 17742 15428
rect 18049 15419 18107 15425
rect 18049 15416 18061 15419
rect 17736 15388 18061 15416
rect 17736 15376 17742 15388
rect 18049 15385 18061 15388
rect 18095 15416 18107 15419
rect 20073 15419 20131 15425
rect 20073 15416 20085 15419
rect 18095 15388 19840 15416
rect 18095 15385 18107 15388
rect 18049 15379 18107 15385
rect 3142 15308 3148 15360
rect 3200 15348 3206 15360
rect 3881 15351 3939 15357
rect 3881 15348 3893 15351
rect 3200 15320 3893 15348
rect 3200 15308 3206 15320
rect 3881 15317 3893 15320
rect 3927 15317 3939 15351
rect 3881 15311 3939 15317
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 8938 15348 8944 15360
rect 4028 15320 8944 15348
rect 4028 15308 4034 15320
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12676 15320 12817 15348
rect 12676 15308 12682 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 14550 15308 14556 15360
rect 14608 15348 14614 15360
rect 14645 15351 14703 15357
rect 14645 15348 14657 15351
rect 14608 15320 14657 15348
rect 14608 15308 14614 15320
rect 14645 15317 14657 15320
rect 14691 15317 14703 15351
rect 15194 15348 15200 15360
rect 15155 15320 15200 15348
rect 14645 15311 14703 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 17589 15351 17647 15357
rect 17589 15317 17601 15351
rect 17635 15348 17647 15351
rect 17954 15348 17960 15360
rect 17635 15320 17960 15348
rect 17635 15317 17647 15320
rect 17589 15311 17647 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 19705 15351 19763 15357
rect 19705 15348 19717 15351
rect 19392 15320 19717 15348
rect 19392 15308 19398 15320
rect 19705 15317 19717 15320
rect 19751 15317 19763 15351
rect 19812 15348 19840 15388
rect 19904 15388 20085 15416
rect 19904 15348 19932 15388
rect 20073 15385 20085 15388
rect 20119 15416 20131 15419
rect 20530 15416 20536 15428
rect 20119 15388 20536 15416
rect 20119 15385 20131 15388
rect 20073 15379 20131 15385
rect 20530 15376 20536 15388
rect 20588 15376 20594 15428
rect 21545 15419 21603 15425
rect 21545 15385 21557 15419
rect 21591 15385 21603 15419
rect 21545 15379 21603 15385
rect 19812 15320 19932 15348
rect 19705 15311 19763 15317
rect 20254 15308 20260 15360
rect 20312 15348 20318 15360
rect 20809 15351 20867 15357
rect 20809 15348 20821 15351
rect 20312 15320 20821 15348
rect 20312 15308 20318 15320
rect 20809 15317 20821 15320
rect 20855 15348 20867 15351
rect 21082 15348 21088 15360
rect 20855 15320 21088 15348
rect 20855 15317 20867 15320
rect 20809 15311 20867 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21560 15348 21588 15379
rect 22094 15376 22100 15428
rect 22152 15416 22158 15428
rect 22152 15388 22197 15416
rect 22152 15376 22158 15388
rect 22738 15376 22744 15428
rect 22796 15416 22802 15428
rect 23124 15416 23152 15444
rect 22796 15388 23152 15416
rect 23293 15419 23351 15425
rect 22796 15376 22802 15388
rect 23293 15385 23305 15419
rect 23339 15416 23351 15419
rect 23474 15416 23480 15428
rect 23339 15388 23480 15416
rect 23339 15385 23351 15388
rect 23293 15379 23351 15385
rect 23474 15376 23480 15388
rect 23532 15376 23538 15428
rect 27706 15376 27712 15428
rect 27764 15416 27770 15428
rect 27908 15416 27936 15447
rect 28166 15444 28172 15456
rect 28224 15444 28230 15496
rect 29822 15444 29828 15496
rect 29880 15484 29886 15496
rect 30116 15493 30144 15592
rect 30190 15512 30196 15564
rect 30248 15552 30254 15564
rect 32953 15555 33011 15561
rect 32953 15552 32965 15555
rect 30248 15524 32965 15552
rect 30248 15512 30254 15524
rect 32953 15521 32965 15524
rect 32999 15552 33011 15555
rect 34698 15552 34704 15564
rect 32999 15524 34704 15552
rect 32999 15521 33011 15524
rect 32953 15515 33011 15521
rect 34698 15512 34704 15524
rect 34756 15512 34762 15564
rect 30009 15487 30067 15493
rect 30009 15484 30021 15487
rect 29880 15456 30021 15484
rect 29880 15444 29886 15456
rect 30009 15453 30021 15456
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 30101 15487 30159 15493
rect 30101 15453 30113 15487
rect 30147 15453 30159 15487
rect 30101 15447 30159 15453
rect 30377 15487 30435 15493
rect 30377 15453 30389 15487
rect 30423 15453 30435 15487
rect 30377 15447 30435 15453
rect 27764 15388 27936 15416
rect 30193 15419 30251 15425
rect 27764 15376 27770 15388
rect 30193 15385 30205 15419
rect 30239 15385 30251 15419
rect 30392 15416 30420 15447
rect 30466 15444 30472 15496
rect 30524 15484 30530 15496
rect 31205 15487 31263 15493
rect 31205 15484 31217 15487
rect 30524 15456 31217 15484
rect 30524 15444 30530 15456
rect 31205 15453 31217 15456
rect 31251 15453 31263 15487
rect 31205 15447 31263 15453
rect 32306 15444 32312 15496
rect 32364 15484 32370 15496
rect 33965 15487 34023 15493
rect 33965 15484 33977 15487
rect 32364 15456 33977 15484
rect 32364 15444 32370 15456
rect 33965 15453 33977 15456
rect 34011 15453 34023 15487
rect 34146 15484 34152 15496
rect 34107 15456 34152 15484
rect 33965 15447 34023 15453
rect 34146 15444 34152 15456
rect 34204 15444 34210 15496
rect 35268 15493 35296 15592
rect 35986 15580 35992 15592
rect 36044 15580 36050 15632
rect 38933 15555 38991 15561
rect 35360 15524 35664 15552
rect 35253 15487 35311 15493
rect 35253 15453 35265 15487
rect 35299 15453 35311 15487
rect 35253 15447 35311 15453
rect 32766 15416 32772 15428
rect 30392 15388 32772 15416
rect 30193 15379 30251 15385
rect 22186 15348 22192 15360
rect 21560 15320 22192 15348
rect 22186 15308 22192 15320
rect 22244 15308 22250 15360
rect 22370 15308 22376 15360
rect 22428 15348 22434 15360
rect 22557 15351 22615 15357
rect 22557 15348 22569 15351
rect 22428 15320 22569 15348
rect 22428 15308 22434 15320
rect 22557 15317 22569 15320
rect 22603 15317 22615 15351
rect 28258 15348 28264 15360
rect 28219 15320 28264 15348
rect 22557 15311 22615 15317
rect 28258 15308 28264 15320
rect 28316 15308 28322 15360
rect 28626 15308 28632 15360
rect 28684 15348 28690 15360
rect 28721 15351 28779 15357
rect 28721 15348 28733 15351
rect 28684 15320 28733 15348
rect 28684 15308 28690 15320
rect 28721 15317 28733 15320
rect 28767 15317 28779 15351
rect 28721 15311 28779 15317
rect 29825 15351 29883 15357
rect 29825 15317 29837 15351
rect 29871 15348 29883 15351
rect 29914 15348 29920 15360
rect 29871 15320 29920 15348
rect 29871 15317 29883 15320
rect 29825 15311 29883 15317
rect 29914 15308 29920 15320
rect 29972 15308 29978 15360
rect 30208 15348 30236 15379
rect 32766 15376 32772 15388
rect 32824 15376 32830 15428
rect 35360 15416 35388 15524
rect 35636 15493 35664 15524
rect 38933 15521 38945 15555
rect 38979 15552 38991 15555
rect 39114 15552 39120 15564
rect 38979 15524 39120 15552
rect 38979 15521 38991 15524
rect 38933 15515 38991 15521
rect 39114 15512 39120 15524
rect 39172 15512 39178 15564
rect 35437 15487 35495 15493
rect 35437 15453 35449 15487
rect 35483 15453 35495 15487
rect 35437 15447 35495 15453
rect 35529 15487 35587 15493
rect 35529 15453 35541 15487
rect 35575 15453 35587 15487
rect 35529 15447 35587 15453
rect 35621 15487 35679 15493
rect 35621 15453 35633 15487
rect 35667 15453 35679 15487
rect 35621 15447 35679 15453
rect 34716 15388 35388 15416
rect 30466 15348 30472 15360
rect 30208 15320 30472 15348
rect 30466 15308 30472 15320
rect 30524 15308 30530 15360
rect 34606 15308 34612 15360
rect 34664 15348 34670 15360
rect 34716 15357 34744 15388
rect 34701 15351 34759 15357
rect 34701 15348 34713 15351
rect 34664 15320 34713 15348
rect 34664 15308 34670 15320
rect 34701 15317 34713 15320
rect 34747 15317 34759 15351
rect 35452 15348 35480 15447
rect 35544 15416 35572 15447
rect 35710 15416 35716 15428
rect 35544 15388 35716 15416
rect 35710 15376 35716 15388
rect 35768 15376 35774 15428
rect 35897 15419 35955 15425
rect 35897 15385 35909 15419
rect 35943 15416 35955 15419
rect 38666 15419 38724 15425
rect 38666 15416 38678 15419
rect 35943 15388 38678 15416
rect 35943 15385 35955 15388
rect 35897 15379 35955 15385
rect 38666 15385 38678 15388
rect 38712 15385 38724 15419
rect 38666 15379 38724 15385
rect 36170 15348 36176 15360
rect 35452 15320 36176 15348
rect 34701 15311 34759 15317
rect 36170 15308 36176 15320
rect 36228 15308 36234 15360
rect 37550 15348 37556 15360
rect 37511 15320 37556 15348
rect 37550 15308 37556 15320
rect 37608 15308 37614 15360
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7524 15116 7849 15144
rect 7524 15104 7530 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 9861 15147 9919 15153
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 10410 15144 10416 15156
rect 9907 15116 10416 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10502 15104 10508 15156
rect 10560 15104 10566 15156
rect 11698 15144 11704 15156
rect 11659 15116 11704 15144
rect 11698 15104 11704 15116
rect 11756 15144 11762 15156
rect 11756 15116 12848 15144
rect 11756 15104 11762 15116
rect 4798 15076 4804 15088
rect 3988 15048 4804 15076
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 15008 2467 15011
rect 2774 15008 2780 15020
rect 2455 14980 2780 15008
rect 2455 14977 2467 14980
rect 2409 14971 2467 14977
rect 2774 14968 2780 14980
rect 2832 15008 2838 15020
rect 3142 15008 3148 15020
rect 2832 14980 3148 15008
rect 2832 14968 2838 14980
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 3694 15008 3700 15020
rect 3607 14980 3700 15008
rect 3694 14968 3700 14980
rect 3752 14968 3758 15020
rect 3878 15008 3884 15020
rect 3839 14980 3884 15008
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 3988 15017 4016 15048
rect 4798 15036 4804 15048
rect 4856 15036 4862 15088
rect 4893 15079 4951 15085
rect 4893 15045 4905 15079
rect 4939 15076 4951 15079
rect 5166 15076 5172 15088
rect 4939 15048 5172 15076
rect 4939 15045 4951 15048
rect 4893 15039 4951 15045
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 15008 4123 15011
rect 4908 15008 4936 15039
rect 5166 15036 5172 15048
rect 5224 15036 5230 15088
rect 6825 15079 6883 15085
rect 6825 15045 6837 15079
rect 6871 15076 6883 15079
rect 7282 15076 7288 15088
rect 6871 15048 7288 15076
rect 6871 15045 6883 15048
rect 6825 15039 6883 15045
rect 7282 15036 7288 15048
rect 7340 15036 7346 15088
rect 8018 15076 8024 15088
rect 7979 15048 8024 15076
rect 8018 15036 8024 15048
rect 8076 15036 8082 15088
rect 9033 15079 9091 15085
rect 8680 15048 8984 15076
rect 4111 14980 4936 15008
rect 4111 14977 4123 14980
rect 4065 14971 4123 14977
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6236 14980 6653 15008
rect 6236 14968 6242 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 6917 15011 6975 15017
rect 6917 15008 6929 15011
rect 6788 14980 6929 15008
rect 6788 14968 6794 14980
rect 6917 14977 6929 14980
rect 6963 14977 6975 15011
rect 6917 14971 6975 14977
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 8205 15011 8263 15017
rect 7064 14980 7109 15008
rect 7064 14968 7070 14980
rect 8205 14977 8217 15011
rect 8251 15008 8263 15011
rect 8294 15008 8300 15020
rect 8251 14980 8300 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2590 14940 2596 14952
rect 2280 14912 2596 14940
rect 2280 14900 2286 14912
rect 2590 14900 2596 14912
rect 2648 14940 2654 14952
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 2648 14912 2697 14940
rect 2648 14900 2654 14912
rect 2685 14909 2697 14912
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 2958 14900 2964 14952
rect 3016 14940 3022 14952
rect 3712 14940 3740 14968
rect 3016 14912 3740 14940
rect 3016 14900 3022 14912
rect 1670 14832 1676 14884
rect 1728 14872 1734 14884
rect 6748 14872 6776 14968
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 8220 14940 8248 14971
rect 8294 14968 8300 14980
rect 8352 15008 8358 15020
rect 8680 15017 8708 15048
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 8352 14980 8677 15008
rect 8352 14968 8358 14980
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8956 15008 8984 15048
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 10520 15076 10548 15104
rect 9079 15048 10456 15076
rect 10520 15048 10640 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 8956 14980 9505 15008
rect 8849 14971 8907 14977
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 6880 14912 8248 14940
rect 6880 14900 6886 14912
rect 1728 14844 6776 14872
rect 7193 14875 7251 14881
rect 1728 14832 1734 14844
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 8202 14872 8208 14884
rect 7239 14844 8208 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 8202 14832 8208 14844
rect 8260 14832 8266 14884
rect 4341 14807 4399 14813
rect 4341 14773 4353 14807
rect 4387 14804 4399 14807
rect 4614 14804 4620 14816
rect 4387 14776 4620 14804
rect 4387 14773 4399 14776
rect 4341 14767 4399 14773
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 8864 14804 8892 14971
rect 9692 14940 9720 14971
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 10318 15008 10324 15020
rect 9824 14980 10324 15008
rect 9824 14968 9830 14980
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 10428 15011 10456 15048
rect 10484 15014 10542 15020
rect 10612 15017 10640 15048
rect 12434 15036 12440 15088
rect 12492 15076 12498 15088
rect 12529 15079 12587 15085
rect 12529 15076 12541 15079
rect 12492 15048 12541 15076
rect 12492 15036 12498 15048
rect 12529 15045 12541 15048
rect 12575 15045 12587 15079
rect 12529 15039 12587 15045
rect 10484 15011 10496 15014
rect 10428 14983 10496 15011
rect 10484 14980 10496 14983
rect 10530 14980 10542 15014
rect 10484 14974 10542 14980
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 14977 10655 15011
rect 10597 14971 10655 14977
rect 10686 14968 10692 15020
rect 10744 15017 10750 15020
rect 10744 15011 10767 15017
rect 10755 14977 10767 15011
rect 10744 14971 10767 14977
rect 10744 14968 10750 14971
rect 10962 14968 10968 15020
rect 11020 15008 11026 15020
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 11020 14980 11529 15008
rect 11020 14968 11026 14980
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 12820 15008 12848 15116
rect 15010 15104 15016 15156
rect 15068 15144 15074 15156
rect 18966 15144 18972 15156
rect 15068 15116 18972 15144
rect 15068 15104 15074 15116
rect 18966 15104 18972 15116
rect 19024 15104 19030 15156
rect 19245 15147 19303 15153
rect 19245 15113 19257 15147
rect 19291 15113 19303 15147
rect 19245 15107 19303 15113
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20346 15144 20352 15156
rect 19935 15116 20352 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 12894 15036 12900 15088
rect 12952 15076 12958 15088
rect 14185 15079 14243 15085
rect 14185 15076 14197 15079
rect 12952 15048 14197 15076
rect 12952 15036 12958 15048
rect 14185 15045 14197 15048
rect 14231 15076 14243 15079
rect 15378 15076 15384 15088
rect 14231 15048 15384 15076
rect 14231 15045 14243 15048
rect 14185 15039 14243 15045
rect 14752 15017 14780 15048
rect 15378 15036 15384 15048
rect 15436 15076 15442 15088
rect 15436 15048 17908 15076
rect 15436 15036 15442 15048
rect 14737 15011 14795 15017
rect 12820 14980 14596 15008
rect 11517 14971 11575 14977
rect 11606 14940 11612 14952
rect 9692 14912 11612 14940
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 14366 14940 14372 14952
rect 11756 14912 14372 14940
rect 11756 14900 11762 14912
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 10965 14875 11023 14881
rect 10965 14841 10977 14875
rect 11011 14872 11023 14875
rect 12526 14872 12532 14884
rect 11011 14844 12532 14872
rect 11011 14841 11023 14844
rect 10965 14835 11023 14841
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 11514 14804 11520 14816
rect 8864 14776 11520 14804
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 14568 14804 14596 14980
rect 14737 14977 14749 15011
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 14993 15011 15051 15017
rect 14993 15008 15005 15011
rect 14884 14980 15005 15008
rect 14884 14968 14890 14980
rect 14993 14977 15005 14980
rect 15039 14977 15051 15011
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 14993 14971 15051 14977
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 17034 15008 17040 15020
rect 16995 14980 17040 15008
rect 16853 14971 16911 14977
rect 16868 14940 16896 14971
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 17880 15017 17908 15048
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 18110 15079 18168 15085
rect 18110 15076 18122 15079
rect 18012 15048 18122 15076
rect 18012 15036 18018 15048
rect 18110 15045 18122 15048
rect 18156 15045 18168 15079
rect 18110 15039 18168 15045
rect 19260 15076 19288 15107
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 20772 15116 21312 15144
rect 20772 15104 20778 15116
rect 20806 15076 20812 15088
rect 19260 15048 20812 15076
rect 17865 15011 17923 15017
rect 17865 14977 17877 15011
rect 17911 14977 17923 15011
rect 19260 15008 19288 15048
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 21284 15085 21312 15116
rect 22646 15104 22652 15156
rect 22704 15144 22710 15156
rect 28534 15144 28540 15156
rect 22704 15116 28540 15144
rect 22704 15104 22710 15116
rect 28534 15104 28540 15116
rect 28592 15104 28598 15156
rect 29546 15144 29552 15156
rect 29507 15116 29552 15144
rect 29546 15104 29552 15116
rect 29604 15104 29610 15156
rect 30374 15144 30380 15156
rect 30335 15116 30380 15144
rect 30374 15104 30380 15116
rect 30432 15104 30438 15156
rect 36170 15144 36176 15156
rect 36131 15116 36176 15144
rect 36170 15104 36176 15116
rect 36228 15104 36234 15156
rect 39298 15104 39304 15156
rect 39356 15144 39362 15156
rect 39669 15147 39727 15153
rect 39669 15144 39681 15147
rect 39356 15116 39681 15144
rect 39356 15104 39362 15116
rect 39669 15113 39681 15116
rect 39715 15144 39727 15147
rect 40218 15144 40224 15156
rect 39715 15116 40224 15144
rect 39715 15113 39727 15116
rect 39669 15107 39727 15113
rect 40218 15104 40224 15116
rect 40276 15104 40282 15156
rect 21269 15079 21327 15085
rect 21269 15045 21281 15079
rect 21315 15045 21327 15079
rect 21269 15039 21327 15045
rect 21358 15036 21364 15088
rect 21416 15076 21422 15088
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 21416 15048 21833 15076
rect 21416 15036 21422 15048
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 24302 15076 24308 15088
rect 21821 15039 21879 15045
rect 22020 15048 24308 15076
rect 17865 14971 17923 14977
rect 17972 14980 19288 15008
rect 20257 15011 20315 15017
rect 17972 14940 18000 14980
rect 20257 14977 20269 15011
rect 20303 15008 20315 15011
rect 20622 15008 20628 15020
rect 20303 14980 20628 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 15008 21051 15011
rect 22020 15008 22048 15048
rect 24302 15036 24308 15048
rect 24360 15036 24366 15088
rect 25900 15079 25958 15085
rect 25900 15045 25912 15079
rect 25946 15076 25958 15079
rect 26973 15079 27031 15085
rect 26973 15076 26985 15079
rect 25946 15048 26985 15076
rect 25946 15045 25958 15048
rect 25900 15039 25958 15045
rect 26973 15045 26985 15048
rect 27019 15045 27031 15079
rect 26973 15039 27031 15045
rect 27080 15048 27476 15076
rect 21039 14980 22048 15008
rect 22097 15011 22155 15017
rect 21039 14977 21051 14980
rect 20993 14971 21051 14977
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22830 15008 22836 15020
rect 22143 14980 22836 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22830 14968 22836 14980
rect 22888 14968 22894 15020
rect 23014 15017 23020 15020
rect 23008 14971 23020 15017
rect 23072 15008 23078 15020
rect 23072 14980 23108 15008
rect 23014 14968 23020 14971
rect 23072 14968 23078 14980
rect 26694 14968 26700 15020
rect 26752 15008 26758 15020
rect 27080 15008 27108 15048
rect 27448 15017 27476 15048
rect 28258 15036 28264 15088
rect 28316 15076 28322 15088
rect 28414 15079 28472 15085
rect 28414 15076 28426 15079
rect 28316 15048 28426 15076
rect 28316 15036 28322 15048
rect 28414 15045 28426 15048
rect 28460 15045 28472 15079
rect 28414 15039 28472 15045
rect 31113 15079 31171 15085
rect 31113 15045 31125 15079
rect 31159 15076 31171 15079
rect 32306 15076 32312 15088
rect 31159 15048 32312 15076
rect 31159 15045 31171 15048
rect 31113 15039 31171 15045
rect 32306 15036 32312 15048
rect 32364 15036 32370 15088
rect 33505 15079 33563 15085
rect 33505 15045 33517 15079
rect 33551 15076 33563 15079
rect 33965 15079 34023 15085
rect 33965 15076 33977 15079
rect 33551 15048 33977 15076
rect 33551 15045 33563 15048
rect 33505 15039 33563 15045
rect 33965 15045 33977 15048
rect 34011 15076 34023 15079
rect 34698 15076 34704 15088
rect 34011 15048 34704 15076
rect 34011 15045 34023 15048
rect 33965 15039 34023 15045
rect 34698 15036 34704 15048
rect 34756 15076 34762 15088
rect 35342 15076 35348 15088
rect 34756 15048 35348 15076
rect 34756 15036 34762 15048
rect 35342 15036 35348 15048
rect 35400 15036 35406 15088
rect 37550 15076 37556 15088
rect 36372 15048 37556 15076
rect 26752 14980 27108 15008
rect 27249 15011 27307 15017
rect 26752 14968 26758 14980
rect 27249 14977 27261 15011
rect 27295 14977 27307 15011
rect 27249 14971 27307 14977
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 27433 15011 27491 15017
rect 27433 14977 27445 15011
rect 27479 14977 27491 15011
rect 27433 14971 27491 14977
rect 27617 15011 27675 15017
rect 27617 14977 27629 15011
rect 27663 15008 27675 15011
rect 28718 15008 28724 15020
rect 27663 14980 28724 15008
rect 27663 14977 27675 14980
rect 27617 14971 27675 14977
rect 16868 14912 18000 14940
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 21177 14943 21235 14949
rect 21177 14909 21189 14943
rect 21223 14909 21235 14943
rect 21910 14940 21916 14952
rect 21871 14912 21916 14940
rect 21177 14903 21235 14909
rect 16114 14872 16120 14884
rect 16075 14844 16120 14872
rect 16114 14832 16120 14844
rect 16172 14832 16178 14884
rect 17862 14872 17868 14884
rect 16592 14844 17868 14872
rect 16592 14804 16620 14844
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 20180 14872 20208 14903
rect 20809 14875 20867 14881
rect 20809 14872 20821 14875
rect 20180 14844 20821 14872
rect 20809 14841 20821 14844
rect 20855 14841 20867 14875
rect 20809 14835 20867 14841
rect 21192 14816 21220 14903
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 22002 14900 22008 14952
rect 22060 14940 22066 14952
rect 22741 14943 22799 14949
rect 22741 14940 22753 14943
rect 22060 14912 22753 14940
rect 22060 14900 22066 14912
rect 22741 14909 22753 14912
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 26145 14943 26203 14949
rect 26145 14909 26157 14943
rect 26191 14940 26203 14943
rect 26786 14940 26792 14952
rect 26191 14912 26792 14940
rect 26191 14909 26203 14912
rect 26145 14903 26203 14909
rect 26786 14900 26792 14912
rect 26844 14900 26850 14952
rect 22646 14872 22652 14884
rect 21284 14844 22652 14872
rect 14568 14776 16620 14804
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 18138 14804 18144 14816
rect 16724 14776 18144 14804
rect 16724 14764 16730 14776
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 18598 14764 18604 14816
rect 18656 14804 18662 14816
rect 20073 14807 20131 14813
rect 20073 14804 20085 14807
rect 18656 14776 20085 14804
rect 18656 14764 18662 14776
rect 20073 14773 20085 14776
rect 20119 14773 20131 14807
rect 20073 14767 20131 14773
rect 21174 14764 21180 14816
rect 21232 14764 21238 14816
rect 21284 14813 21312 14844
rect 22646 14832 22652 14844
rect 22704 14832 22710 14884
rect 24762 14872 24768 14884
rect 24723 14844 24768 14872
rect 24762 14832 24768 14844
rect 24820 14832 24826 14884
rect 21269 14807 21327 14813
rect 21269 14773 21281 14807
rect 21315 14773 21327 14807
rect 21818 14804 21824 14816
rect 21779 14776 21824 14804
rect 21269 14767 21327 14773
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 22278 14804 22284 14816
rect 22239 14776 22284 14804
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 24121 14807 24179 14813
rect 24121 14804 24133 14807
rect 23992 14776 24133 14804
rect 23992 14764 23998 14776
rect 24121 14773 24133 14776
rect 24167 14773 24179 14807
rect 24121 14767 24179 14773
rect 26418 14764 26424 14816
rect 26476 14804 26482 14816
rect 27264 14804 27292 14971
rect 27356 14872 27384 14971
rect 28718 14968 28724 14980
rect 28776 14968 28782 15020
rect 30742 14968 30748 15020
rect 30800 15008 30806 15020
rect 30926 15008 30932 15020
rect 30800 14980 30932 15008
rect 30800 14968 30806 14980
rect 30926 14968 30932 14980
rect 30984 15008 30990 15020
rect 31021 15011 31079 15017
rect 31021 15008 31033 15011
rect 30984 14980 31033 15008
rect 30984 14968 30990 14980
rect 31021 14977 31033 14980
rect 31067 14977 31079 15011
rect 31202 15008 31208 15020
rect 31163 14980 31208 15008
rect 31021 14971 31079 14977
rect 31202 14968 31208 14980
rect 31260 14968 31266 15020
rect 31389 15011 31447 15017
rect 31389 14977 31401 15011
rect 31435 15008 31447 15011
rect 31478 15008 31484 15020
rect 31435 14980 31484 15008
rect 31435 14977 31447 14980
rect 31389 14971 31447 14977
rect 31478 14968 31484 14980
rect 31536 14968 31542 15020
rect 32950 14968 32956 15020
rect 33008 15008 33014 15020
rect 36372 15017 36400 15048
rect 37550 15036 37556 15048
rect 37608 15036 37614 15088
rect 36357 15011 36415 15017
rect 36357 15008 36369 15011
rect 33008 14980 36369 15008
rect 33008 14968 33014 14980
rect 36357 14977 36369 14980
rect 36403 14977 36415 15011
rect 36357 14971 36415 14977
rect 36541 15011 36599 15017
rect 36541 14977 36553 15011
rect 36587 15008 36599 15011
rect 37642 15008 37648 15020
rect 36587 14980 37648 15008
rect 36587 14977 36599 14980
rect 36541 14971 36599 14977
rect 37642 14968 37648 14980
rect 37700 14968 37706 15020
rect 27522 14900 27528 14952
rect 27580 14940 27586 14952
rect 28169 14943 28227 14949
rect 28169 14940 28181 14943
rect 27580 14912 28181 14940
rect 27580 14900 27586 14912
rect 28169 14909 28181 14912
rect 28215 14909 28227 14943
rect 28169 14903 28227 14909
rect 27706 14872 27712 14884
rect 27356 14844 27712 14872
rect 27706 14832 27712 14844
rect 27764 14832 27770 14884
rect 30926 14872 30932 14884
rect 29104 14844 30932 14872
rect 29104 14804 29132 14844
rect 30926 14832 30932 14844
rect 30984 14872 30990 14884
rect 34606 14872 34612 14884
rect 30984 14844 34612 14872
rect 30984 14832 30990 14844
rect 34606 14832 34612 14844
rect 34664 14832 34670 14884
rect 30834 14804 30840 14816
rect 26476 14776 29132 14804
rect 30795 14776 30840 14804
rect 26476 14764 26482 14776
rect 30834 14764 30840 14776
rect 30892 14764 30898 14816
rect 32674 14764 32680 14816
rect 32732 14804 32738 14816
rect 35253 14807 35311 14813
rect 35253 14804 35265 14807
rect 32732 14776 35265 14804
rect 32732 14764 32738 14776
rect 35253 14773 35265 14776
rect 35299 14804 35311 14807
rect 35894 14804 35900 14816
rect 35299 14776 35900 14804
rect 35299 14773 35311 14776
rect 35253 14767 35311 14773
rect 35894 14764 35900 14776
rect 35952 14764 35958 14816
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 3936 14572 6009 14600
rect 3936 14560 3942 14572
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 8110 14600 8116 14612
rect 7515 14572 8116 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 11057 14603 11115 14609
rect 8996 14572 11008 14600
rect 8996 14560 9002 14572
rect 5353 14535 5411 14541
rect 5353 14501 5365 14535
rect 5399 14532 5411 14535
rect 6178 14532 6184 14544
rect 5399 14504 6184 14532
rect 5399 14501 5411 14504
rect 5353 14495 5411 14501
rect 6178 14492 6184 14504
rect 6236 14492 6242 14544
rect 7558 14532 7564 14544
rect 6564 14504 7564 14532
rect 3786 14464 3792 14476
rect 2516 14436 3792 14464
rect 2516 14405 2544 14436
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 6564 14464 6592 14504
rect 7558 14492 7564 14504
rect 7616 14532 7622 14544
rect 7929 14535 7987 14541
rect 7929 14532 7941 14535
rect 7616 14504 7941 14532
rect 7616 14492 7622 14504
rect 7929 14501 7941 14504
rect 7975 14532 7987 14535
rect 10502 14532 10508 14544
rect 7975 14504 10508 14532
rect 7975 14501 7987 14504
rect 7929 14495 7987 14501
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 9585 14467 9643 14473
rect 6012 14436 6592 14464
rect 7392 14436 9168 14464
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 2501 14399 2559 14405
rect 1903 14368 2360 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 2332 14272 2360 14368
rect 2501 14365 2513 14399
rect 2547 14365 2559 14399
rect 2501 14359 2559 14365
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14396 2743 14399
rect 3145 14399 3203 14405
rect 3145 14396 3157 14399
rect 2731 14368 3157 14396
rect 2731 14365 2743 14368
rect 2685 14359 2743 14365
rect 3145 14365 3157 14368
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4062 14396 4068 14408
rect 4019 14368 4068 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 3160 14328 3188 14359
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4240 14399 4298 14405
rect 4240 14365 4252 14399
rect 4286 14396 4298 14399
rect 4614 14396 4620 14408
rect 4286 14368 4620 14396
rect 4286 14365 4298 14368
rect 4240 14359 4298 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 6012 14396 6040 14436
rect 6178 14396 6184 14408
rect 4856 14368 6040 14396
rect 6139 14368 6184 14396
rect 4856 14356 4862 14368
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 6822 14396 6828 14408
rect 6411 14368 6828 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 7098 14396 7104 14408
rect 7011 14368 7104 14396
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7282 14356 7288 14408
rect 7340 14405 7346 14408
rect 7340 14399 7363 14405
rect 7351 14396 7363 14399
rect 7392 14396 7420 14436
rect 9140 14408 9168 14436
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 10778 14464 10784 14476
rect 9631 14436 10784 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 8938 14396 8944 14408
rect 7351 14368 7433 14396
rect 8899 14368 8944 14396
rect 7351 14365 7363 14368
rect 7340 14359 7363 14365
rect 7340 14356 7346 14359
rect 8938 14356 8944 14368
rect 8996 14356 9002 14408
rect 9122 14396 9128 14408
rect 9083 14368 9128 14396
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9364 14368 9873 14396
rect 9364 14356 9370 14368
rect 9861 14365 9873 14368
rect 9907 14365 9919 14399
rect 10980 14396 11008 14572
rect 11057 14569 11069 14603
rect 11103 14600 11115 14603
rect 14274 14600 14280 14612
rect 11103 14572 12940 14600
rect 14235 14572 14280 14600
rect 11103 14569 11115 14572
rect 11057 14563 11115 14569
rect 11514 14532 11520 14544
rect 11475 14504 11520 14532
rect 11514 14492 11520 14504
rect 11572 14532 11578 14544
rect 11790 14532 11796 14544
rect 11572 14504 11796 14532
rect 11572 14492 11578 14504
rect 11790 14492 11796 14504
rect 11848 14492 11854 14544
rect 12912 14532 12940 14572
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 14918 14600 14924 14612
rect 14384 14572 14924 14600
rect 12986 14532 12992 14544
rect 12912 14504 12992 14532
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 14384 14532 14412 14572
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 16574 14600 16580 14612
rect 16535 14572 16580 14600
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17126 14560 17132 14612
rect 17184 14600 17190 14612
rect 17405 14603 17463 14609
rect 17405 14600 17417 14603
rect 17184 14572 17417 14600
rect 17184 14560 17190 14572
rect 17405 14569 17417 14572
rect 17451 14569 17463 14603
rect 18598 14600 18604 14612
rect 18559 14572 18604 14600
rect 17405 14563 17463 14569
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 20530 14560 20536 14612
rect 20588 14600 20594 14612
rect 21545 14603 21603 14609
rect 21545 14600 21557 14603
rect 20588 14572 21557 14600
rect 20588 14560 20594 14572
rect 21545 14569 21557 14572
rect 21591 14600 21603 14603
rect 22370 14600 22376 14612
rect 21591 14572 22376 14600
rect 21591 14569 21603 14572
rect 21545 14563 21603 14569
rect 22370 14560 22376 14572
rect 22428 14560 22434 14612
rect 24670 14600 24676 14612
rect 24631 14572 24676 14600
rect 24670 14560 24676 14572
rect 24728 14560 24734 14612
rect 26694 14600 26700 14612
rect 26655 14572 26700 14600
rect 26694 14560 26700 14572
rect 26752 14560 26758 14612
rect 26786 14560 26792 14612
rect 26844 14600 26850 14612
rect 27430 14600 27436 14612
rect 26844 14572 27436 14600
rect 26844 14560 26850 14572
rect 27430 14560 27436 14572
rect 27488 14560 27494 14612
rect 27525 14603 27583 14609
rect 27525 14569 27537 14603
rect 27571 14600 27583 14603
rect 28166 14600 28172 14612
rect 27571 14572 28172 14600
rect 27571 14569 27583 14572
rect 27525 14563 27583 14569
rect 28166 14560 28172 14572
rect 28224 14560 28230 14612
rect 28718 14560 28724 14612
rect 28776 14600 28782 14612
rect 33042 14600 33048 14612
rect 28776 14572 33048 14600
rect 28776 14560 28782 14572
rect 33042 14560 33048 14572
rect 33100 14560 33106 14612
rect 37737 14603 37795 14609
rect 37737 14600 37749 14603
rect 33244 14572 37749 14600
rect 16298 14532 16304 14544
rect 13587 14504 14412 14532
rect 14476 14504 16304 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 12894 14464 12900 14476
rect 12855 14436 12900 14464
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 12066 14396 12072 14408
rect 10980 14368 12072 14396
rect 9861 14359 9919 14365
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 12912 14396 12940 14424
rect 14476 14405 14504 14504
rect 16298 14492 16304 14504
rect 16356 14492 16362 14544
rect 24857 14535 24915 14541
rect 24857 14532 24869 14535
rect 16500 14504 24869 14532
rect 12406 14368 12940 14396
rect 14369 14399 14427 14405
rect 6454 14328 6460 14340
rect 3160 14300 6460 14328
rect 6454 14288 6460 14300
rect 6512 14328 6518 14340
rect 7116 14328 7144 14356
rect 6512 14300 7144 14328
rect 8113 14331 8171 14337
rect 6512 14288 6518 14300
rect 8113 14297 8125 14331
rect 8159 14328 8171 14331
rect 8294 14328 8300 14340
rect 8159 14300 8300 14328
rect 8159 14297 8171 14300
rect 8113 14291 8171 14297
rect 8294 14288 8300 14300
rect 8352 14328 8358 14340
rect 9033 14331 9091 14337
rect 9033 14328 9045 14331
rect 8352 14300 9045 14328
rect 8352 14288 8358 14300
rect 9033 14297 9045 14300
rect 9079 14297 9091 14331
rect 9033 14291 9091 14297
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 12406 14328 12434 14368
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14918 14396 14924 14408
rect 14879 14368 14924 14396
rect 14461 14359 14519 14365
rect 9732 14300 12434 14328
rect 9732 14288 9738 14300
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 12630 14331 12688 14337
rect 12630 14328 12642 14331
rect 12584 14300 12642 14328
rect 12584 14288 12590 14300
rect 12630 14297 12642 14300
rect 12676 14297 12688 14331
rect 14384 14328 14412 14359
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 16500 14328 16528 14504
rect 24857 14501 24869 14504
rect 24903 14501 24915 14535
rect 28184 14532 28212 14560
rect 28902 14532 28908 14544
rect 28184 14504 28908 14532
rect 24857 14495 24915 14501
rect 28902 14492 28908 14504
rect 28960 14492 28966 14544
rect 33134 14532 33140 14544
rect 32140 14504 33140 14532
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14464 16635 14467
rect 16623 14436 19380 14464
rect 16623 14433 16635 14436
rect 16577 14427 16635 14433
rect 16666 14396 16672 14408
rect 16627 14368 16672 14396
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17586 14396 17592 14408
rect 17547 14368 17592 14396
rect 17405 14359 17463 14365
rect 14384 14300 16528 14328
rect 17420 14328 17448 14359
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 19352 14396 19380 14436
rect 19978 14424 19984 14476
rect 20036 14464 20042 14476
rect 20898 14464 20904 14476
rect 20036 14436 20904 14464
rect 20036 14424 20042 14436
rect 20898 14424 20904 14436
rect 20956 14424 20962 14476
rect 21634 14424 21640 14476
rect 21692 14464 21698 14476
rect 24486 14464 24492 14476
rect 21692 14436 24256 14464
rect 24447 14436 24492 14464
rect 21692 14424 21698 14436
rect 22738 14396 22744 14408
rect 19352 14368 22744 14396
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 19334 14328 19340 14340
rect 17420 14300 19340 14328
rect 12630 14291 12688 14297
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 20714 14328 20720 14340
rect 19812 14300 20720 14328
rect 1578 14220 1584 14272
rect 1636 14260 1642 14272
rect 1673 14263 1731 14269
rect 1673 14260 1685 14263
rect 1636 14232 1685 14260
rect 1636 14220 1642 14232
rect 1673 14229 1685 14232
rect 1719 14229 1731 14263
rect 2314 14260 2320 14272
rect 2275 14232 2320 14260
rect 1673 14223 1731 14229
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 7650 14260 7656 14272
rect 7156 14232 7656 14260
rect 7156 14220 7162 14232
rect 7650 14220 7656 14232
rect 7708 14260 7714 14272
rect 11698 14260 11704 14272
rect 7708 14232 11704 14260
rect 7708 14220 7714 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 12768 14232 14105 14260
rect 12768 14220 12774 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14516 14232 15117 14260
rect 14516 14220 14522 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15838 14260 15844 14272
rect 15799 14232 15844 14260
rect 15105 14223 15163 14229
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 16298 14260 16304 14272
rect 16259 14232 16304 14260
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 17770 14260 17776 14272
rect 17731 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 19245 14263 19303 14269
rect 19245 14229 19257 14263
rect 19291 14260 19303 14263
rect 19426 14260 19432 14272
rect 19291 14232 19432 14260
rect 19291 14229 19303 14232
rect 19245 14223 19303 14229
rect 19426 14220 19432 14232
rect 19484 14260 19490 14272
rect 19812 14260 19840 14300
rect 20714 14288 20720 14300
rect 20772 14288 20778 14340
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 23109 14331 23167 14337
rect 23109 14328 23121 14331
rect 21048 14300 23121 14328
rect 21048 14288 21054 14300
rect 23109 14297 23121 14300
rect 23155 14297 23167 14331
rect 23109 14291 23167 14297
rect 23293 14331 23351 14337
rect 23293 14297 23305 14331
rect 23339 14328 23351 14331
rect 24118 14328 24124 14340
rect 23339 14300 24124 14328
rect 23339 14297 23351 14300
rect 23293 14291 23351 14297
rect 24118 14288 24124 14300
rect 24176 14288 24182 14340
rect 24228 14328 24256 14436
rect 24486 14424 24492 14436
rect 24544 14424 24550 14476
rect 28442 14464 28448 14476
rect 24596 14436 28448 14464
rect 24394 14396 24400 14408
rect 24355 14368 24400 14396
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 24596 14328 24624 14436
rect 28442 14424 28448 14436
rect 28500 14464 28506 14476
rect 28813 14467 28871 14473
rect 28813 14464 28825 14467
rect 28500 14436 28825 14464
rect 28500 14424 28506 14436
rect 28813 14433 28825 14436
rect 28859 14433 28871 14467
rect 28813 14427 28871 14433
rect 30377 14467 30435 14473
rect 30377 14433 30389 14467
rect 30423 14464 30435 14467
rect 30466 14464 30472 14476
rect 30423 14436 30472 14464
rect 30423 14433 30435 14436
rect 30377 14427 30435 14433
rect 30466 14424 30472 14436
rect 30524 14464 30530 14476
rect 30524 14436 32076 14464
rect 30524 14424 30530 14436
rect 24673 14399 24731 14405
rect 24673 14365 24685 14399
rect 24719 14396 24731 14399
rect 24719 14368 28028 14396
rect 24719 14365 24731 14368
rect 24673 14359 24731 14365
rect 26326 14328 26332 14340
rect 24228 14300 24624 14328
rect 26287 14300 26332 14328
rect 26326 14288 26332 14300
rect 26384 14288 26390 14340
rect 26513 14331 26571 14337
rect 26513 14297 26525 14331
rect 26559 14297 26571 14331
rect 28000 14328 28028 14368
rect 28074 14356 28080 14408
rect 28132 14396 28138 14408
rect 28132 14368 28177 14396
rect 28132 14356 28138 14368
rect 28258 14356 28264 14408
rect 28316 14396 28322 14408
rect 30101 14399 30159 14405
rect 30101 14396 30113 14399
rect 28316 14368 30113 14396
rect 28316 14356 28322 14368
rect 30101 14365 30113 14368
rect 30147 14396 30159 14399
rect 31202 14396 31208 14408
rect 30147 14368 31208 14396
rect 30147 14365 30159 14368
rect 30101 14359 30159 14365
rect 31202 14356 31208 14368
rect 31260 14396 31266 14408
rect 31386 14396 31392 14408
rect 31260 14368 31392 14396
rect 31260 14356 31266 14368
rect 31386 14356 31392 14368
rect 31444 14356 31450 14408
rect 31846 14396 31852 14408
rect 31807 14368 31852 14396
rect 31846 14356 31852 14368
rect 31904 14356 31910 14408
rect 32048 14405 32076 14436
rect 32033 14399 32091 14405
rect 32033 14365 32045 14399
rect 32079 14365 32091 14399
rect 32033 14359 32091 14365
rect 31941 14331 31999 14337
rect 28000 14300 31892 14328
rect 26513 14291 26571 14297
rect 19484 14232 19840 14260
rect 19889 14263 19947 14269
rect 19484 14220 19490 14232
rect 19889 14229 19901 14263
rect 19935 14260 19947 14263
rect 20070 14260 20076 14272
rect 19935 14232 20076 14260
rect 19935 14229 19947 14232
rect 19889 14223 19947 14229
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 22097 14263 22155 14269
rect 22097 14229 22109 14263
rect 22143 14260 22155 14263
rect 22186 14260 22192 14272
rect 22143 14232 22192 14260
rect 22143 14229 22155 14232
rect 22097 14223 22155 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22925 14263 22983 14269
rect 22925 14229 22937 14263
rect 22971 14260 22983 14263
rect 23382 14260 23388 14272
rect 22971 14232 23388 14260
rect 22971 14229 22983 14232
rect 22925 14223 22983 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 24762 14220 24768 14272
rect 24820 14260 24826 14272
rect 26528 14260 26556 14291
rect 24820 14232 26556 14260
rect 24820 14220 24826 14232
rect 27982 14220 27988 14272
rect 28040 14260 28046 14272
rect 28261 14263 28319 14269
rect 28261 14260 28273 14263
rect 28040 14232 28273 14260
rect 28040 14220 28046 14232
rect 28261 14229 28273 14232
rect 28307 14229 28319 14263
rect 28261 14223 28319 14229
rect 30558 14220 30564 14272
rect 30616 14260 30622 14272
rect 31665 14263 31723 14269
rect 31665 14260 31677 14263
rect 30616 14232 31677 14260
rect 30616 14220 30622 14232
rect 31665 14229 31677 14232
rect 31711 14229 31723 14263
rect 31864 14260 31892 14300
rect 31941 14297 31953 14331
rect 31987 14328 31999 14331
rect 32140 14328 32168 14504
rect 33134 14492 33140 14504
rect 33192 14492 33198 14544
rect 32217 14399 32275 14405
rect 32217 14365 32229 14399
rect 32263 14365 32275 14399
rect 33134 14396 33140 14408
rect 33095 14368 33140 14396
rect 32217 14359 32275 14365
rect 31987 14300 32168 14328
rect 32232 14328 32260 14359
rect 33134 14356 33140 14368
rect 33192 14356 33198 14408
rect 33244 14405 33272 14572
rect 37737 14569 37749 14572
rect 37783 14600 37795 14603
rect 39942 14600 39948 14612
rect 37783 14572 39948 14600
rect 37783 14569 37795 14572
rect 37737 14563 37795 14569
rect 39942 14560 39948 14572
rect 40000 14560 40006 14612
rect 33229 14399 33287 14405
rect 33229 14365 33241 14399
rect 33275 14365 33287 14399
rect 33229 14359 33287 14365
rect 33505 14399 33563 14405
rect 33505 14365 33517 14399
rect 33551 14396 33563 14399
rect 35802 14396 35808 14408
rect 33551 14368 35808 14396
rect 33551 14365 33563 14368
rect 33505 14359 33563 14365
rect 35802 14356 35808 14368
rect 35860 14356 35866 14408
rect 37090 14396 37096 14408
rect 37051 14368 37096 14396
rect 37090 14356 37096 14368
rect 37148 14356 37154 14408
rect 38838 14356 38844 14408
rect 38896 14405 38902 14408
rect 38896 14399 38919 14405
rect 38907 14365 38919 14399
rect 38896 14359 38919 14365
rect 38896 14356 38902 14359
rect 39022 14356 39028 14408
rect 39080 14396 39086 14408
rect 39128 14399 39186 14405
rect 39128 14396 39140 14399
rect 39080 14368 39140 14396
rect 39080 14356 39086 14368
rect 39128 14365 39140 14368
rect 39174 14365 39186 14399
rect 39128 14359 39186 14365
rect 39390 14356 39396 14408
rect 39448 14396 39454 14408
rect 39853 14399 39911 14405
rect 39853 14396 39865 14399
rect 39448 14368 39865 14396
rect 39448 14356 39454 14368
rect 39853 14365 39865 14368
rect 39899 14365 39911 14399
rect 40016 14399 40074 14405
rect 40016 14396 40028 14399
rect 39853 14359 39911 14365
rect 39960 14368 40028 14396
rect 32232 14300 33272 14328
rect 31987 14297 31999 14300
rect 31941 14291 31999 14297
rect 32953 14263 33011 14269
rect 32953 14260 32965 14263
rect 31864 14232 32965 14260
rect 31665 14223 31723 14229
rect 32953 14229 32965 14232
rect 32999 14229 33011 14263
rect 33244 14260 33272 14300
rect 33318 14288 33324 14340
rect 33376 14328 33382 14340
rect 33376 14300 33421 14328
rect 33376 14288 33382 14300
rect 34606 14288 34612 14340
rect 34664 14328 34670 14340
rect 34885 14331 34943 14337
rect 34885 14328 34897 14331
rect 34664 14300 34897 14328
rect 34664 14288 34670 14300
rect 34885 14297 34897 14300
rect 34931 14297 34943 14331
rect 34885 14291 34943 14297
rect 35069 14331 35127 14337
rect 35069 14297 35081 14331
rect 35115 14328 35127 14331
rect 35158 14328 35164 14340
rect 35115 14300 35164 14328
rect 35115 14297 35127 14300
rect 35069 14291 35127 14297
rect 33410 14260 33416 14272
rect 33244 14232 33416 14260
rect 32953 14223 33011 14229
rect 33410 14220 33416 14232
rect 33468 14220 33474 14272
rect 34701 14263 34759 14269
rect 34701 14229 34713 14263
rect 34747 14260 34759 14263
rect 34790 14260 34796 14272
rect 34747 14232 34796 14260
rect 34747 14229 34759 14232
rect 34701 14223 34759 14229
rect 34790 14220 34796 14232
rect 34848 14220 34854 14272
rect 34900 14260 34928 14291
rect 35158 14288 35164 14300
rect 35216 14288 35222 14340
rect 35434 14288 35440 14340
rect 35492 14328 35498 14340
rect 36826 14331 36884 14337
rect 36826 14328 36838 14331
rect 35492 14300 36838 14328
rect 35492 14288 35498 14300
rect 36826 14297 36838 14300
rect 36872 14297 36884 14331
rect 36826 14291 36884 14297
rect 39758 14288 39764 14340
rect 39816 14328 39822 14340
rect 39960 14328 39988 14368
rect 40016 14365 40028 14368
rect 40062 14365 40074 14399
rect 40016 14359 40074 14365
rect 40129 14399 40187 14405
rect 40129 14365 40141 14399
rect 40175 14365 40187 14399
rect 40129 14359 40187 14365
rect 39816 14300 39988 14328
rect 40144 14328 40172 14359
rect 40218 14356 40224 14408
rect 40276 14405 40282 14408
rect 40276 14399 40299 14405
rect 40287 14365 40299 14399
rect 68094 14396 68100 14408
rect 68055 14368 68100 14396
rect 40276 14359 40299 14365
rect 40276 14356 40282 14359
rect 68094 14356 68100 14368
rect 68152 14356 68158 14408
rect 40494 14328 40500 14340
rect 40144 14300 40264 14328
rect 40455 14300 40500 14328
rect 39816 14288 39822 14300
rect 35713 14263 35771 14269
rect 35713 14260 35725 14263
rect 34900 14232 35725 14260
rect 35713 14229 35725 14232
rect 35759 14229 35771 14263
rect 35713 14223 35771 14229
rect 36446 14220 36452 14272
rect 36504 14260 36510 14272
rect 40236 14260 40264 14300
rect 40494 14288 40500 14300
rect 40552 14288 40558 14340
rect 40310 14260 40316 14272
rect 36504 14232 40316 14260
rect 36504 14220 36510 14232
rect 40310 14220 40316 14232
rect 40368 14220 40374 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 2148 14028 4077 14056
rect 1762 13920 1768 13932
rect 1723 13892 1768 13920
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2148 13929 2176 14028
rect 4065 14025 4077 14028
rect 4111 14056 4123 14059
rect 5534 14056 5540 14068
rect 4111 14028 5540 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 5810 14056 5816 14068
rect 5771 14028 5816 14056
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6512 14028 6561 14056
rect 6512 14016 6518 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 7282 14056 7288 14068
rect 7195 14028 7288 14056
rect 6549 14019 6607 14025
rect 7282 14016 7288 14028
rect 7340 14056 7346 14068
rect 7742 14056 7748 14068
rect 7340 14028 7748 14056
rect 7340 14016 7346 14028
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 10870 14056 10876 14068
rect 10831 14028 10876 14056
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 12161 14059 12219 14065
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 12207 14028 15424 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 2774 13948 2780 14000
rect 2832 13988 2838 14000
rect 5828 13988 5856 14016
rect 7190 13988 7196 14000
rect 2832 13960 3188 13988
rect 5828 13960 7196 13988
rect 2832 13948 2838 13960
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13889 2099 13923
rect 2041 13883 2099 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13889 2191 13923
rect 2869 13923 2927 13929
rect 2869 13920 2881 13923
rect 2133 13883 2191 13889
rect 2792 13892 2881 13920
rect 2056 13852 2084 13883
rect 2222 13852 2228 13864
rect 2056 13824 2228 13852
rect 2222 13812 2228 13824
rect 2280 13812 2286 13864
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2792 13852 2820 13892
rect 2869 13889 2881 13892
rect 2915 13889 2927 13923
rect 3050 13920 3056 13932
rect 3011 13892 3056 13920
rect 2869 13883 2927 13889
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 3160 13929 3188 13960
rect 7190 13948 7196 13960
rect 7248 13988 7254 14000
rect 8294 13988 8300 14000
rect 7248 13960 7880 13988
rect 7248 13948 7254 13960
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13920 3295 13923
rect 5261 13923 5319 13929
rect 3283 13892 5212 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 2958 13852 2964 13864
rect 2455 13824 2728 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2700 13716 2728 13824
rect 2792 13824 2964 13852
rect 2792 13796 2820 13824
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 4614 13852 4620 13864
rect 3068 13824 4620 13852
rect 2774 13744 2780 13796
rect 2832 13744 2838 13796
rect 3068 13716 3096 13824
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5184 13852 5212 13892
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 7098 13920 7104 13932
rect 5307 13892 7104 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 7852 13929 7880 13960
rect 8128 13960 8300 13988
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13889 7895 13923
rect 8018 13920 8024 13932
rect 7979 13892 8024 13920
rect 7837 13883 7895 13889
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8128 13929 8156 13960
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 10505 13991 10563 13997
rect 10505 13988 10517 13991
rect 8956 13960 10517 13988
rect 8956 13929 8984 13960
rect 10505 13957 10517 13960
rect 10551 13988 10563 13991
rect 11514 13988 11520 14000
rect 10551 13960 11520 13988
rect 10551 13957 10563 13960
rect 10505 13951 10563 13957
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 11882 13988 11888 14000
rect 11843 13960 11888 13988
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 14458 13988 14464 14000
rect 12406 13960 14464 13988
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13889 8171 13923
rect 8113 13883 8171 13889
rect 8205 13923 8263 13929
rect 8205 13889 8217 13923
rect 8251 13889 8263 13923
rect 8205 13883 8263 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 6546 13852 6552 13864
rect 5184 13824 6552 13852
rect 6546 13812 6552 13824
rect 6604 13852 6610 13864
rect 8220 13852 8248 13883
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 9180 13892 9229 13920
rect 9180 13880 9186 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 9916 13892 10333 13920
rect 9916 13880 9922 13892
rect 10321 13889 10333 13892
rect 10367 13889 10379 13923
rect 10594 13920 10600 13932
rect 10555 13892 10600 13920
rect 10321 13883 10379 13889
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 10778 13920 10784 13932
rect 10735 13892 10784 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 11606 13920 11612 13932
rect 11567 13892 11612 13920
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11756 13892 11805 13920
rect 11756 13880 11762 13892
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12032 13892 12077 13920
rect 12032 13880 12038 13892
rect 12406 13852 12434 13960
rect 14458 13948 14464 13960
rect 14516 13948 14522 14000
rect 14642 13988 14648 14000
rect 14603 13960 14648 13988
rect 14642 13948 14648 13960
rect 14700 13948 14706 14000
rect 15396 13988 15424 14028
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 15528 14028 15577 14056
rect 15528 14016 15534 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 19886 14056 19892 14068
rect 15896 14028 19892 14056
rect 15896 14016 15902 14028
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 19981 14059 20039 14065
rect 19981 14025 19993 14059
rect 20027 14056 20039 14059
rect 20990 14056 20996 14068
rect 20027 14028 20996 14056
rect 20027 14025 20039 14028
rect 19981 14019 20039 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21269 14059 21327 14065
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 21910 14056 21916 14068
rect 21315 14028 21916 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22830 14016 22836 14068
rect 22888 14056 22894 14068
rect 32861 14059 32919 14065
rect 32861 14056 32873 14059
rect 22888 14028 32873 14056
rect 22888 14016 22894 14028
rect 32861 14025 32873 14028
rect 32907 14025 32919 14059
rect 32861 14019 32919 14025
rect 33042 14016 33048 14068
rect 33100 14056 33106 14068
rect 34057 14059 34115 14065
rect 34057 14056 34069 14059
rect 33100 14028 34069 14056
rect 33100 14016 33106 14028
rect 34057 14025 34069 14028
rect 34103 14056 34115 14059
rect 35345 14059 35403 14065
rect 34103 14028 34744 14056
rect 34103 14025 34115 14028
rect 34057 14019 34115 14025
rect 17402 13988 17408 14000
rect 15396 13960 17408 13988
rect 17402 13948 17408 13960
rect 17460 13948 17466 14000
rect 18868 13991 18926 13997
rect 18868 13957 18880 13991
rect 18914 13988 18926 13991
rect 22925 13991 22983 13997
rect 22925 13988 22937 13991
rect 18914 13960 22937 13988
rect 18914 13957 18926 13960
rect 18868 13951 18926 13957
rect 22925 13957 22937 13960
rect 22971 13957 22983 13991
rect 22925 13951 22983 13957
rect 23934 13948 23940 14000
rect 23992 13988 23998 14000
rect 24213 13991 24271 13997
rect 24213 13988 24225 13991
rect 23992 13960 24225 13988
rect 23992 13948 23998 13960
rect 24213 13957 24225 13960
rect 24259 13957 24271 13991
rect 24213 13951 24271 13957
rect 24949 13991 25007 13997
rect 24949 13957 24961 13991
rect 24995 13988 25007 13991
rect 25406 13988 25412 14000
rect 24995 13960 25412 13988
rect 24995 13957 25007 13960
rect 24949 13951 25007 13957
rect 25406 13948 25412 13960
rect 25464 13948 25470 14000
rect 26418 13988 26424 14000
rect 26379 13960 26424 13988
rect 26418 13948 26424 13960
rect 26476 13948 26482 14000
rect 31297 13991 31355 13997
rect 31297 13957 31309 13991
rect 31343 13988 31355 13991
rect 32950 13988 32956 14000
rect 31343 13960 32956 13988
rect 31343 13957 31355 13960
rect 31297 13951 31355 13957
rect 32950 13948 32956 13960
rect 33008 13948 33014 14000
rect 33137 13991 33195 13997
rect 33137 13957 33149 13991
rect 33183 13988 33195 13991
rect 34606 13988 34612 14000
rect 33183 13960 34612 13988
rect 33183 13957 33195 13960
rect 33137 13951 33195 13957
rect 34606 13948 34612 13960
rect 34664 13948 34670 14000
rect 34716 13988 34744 14028
rect 35345 14025 35357 14059
rect 35391 14056 35403 14059
rect 35434 14056 35440 14068
rect 35391 14028 35440 14056
rect 35391 14025 35403 14028
rect 35345 14019 35403 14025
rect 35434 14016 35440 14028
rect 35492 14016 35498 14068
rect 39298 14056 39304 14068
rect 35544 14028 36584 14056
rect 39259 14028 39304 14056
rect 35544 13988 35572 14028
rect 36446 13988 36452 14000
rect 34716 13960 35572 13988
rect 36277 13960 36452 13988
rect 12986 13920 12992 13932
rect 12947 13892 12992 13920
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13906 13920 13912 13932
rect 13819 13892 13912 13920
rect 13906 13880 13912 13892
rect 13964 13920 13970 13932
rect 14182 13920 14188 13932
rect 13964 13892 14188 13920
rect 13964 13880 13970 13892
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15286 13920 15292 13932
rect 14875 13892 15292 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 15838 13920 15844 13932
rect 15427 13892 15844 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 20530 13920 20536 13932
rect 18064 13892 20536 13920
rect 12894 13852 12900 13864
rect 6604 13824 8248 13852
rect 10888 13824 12434 13852
rect 12855 13824 12900 13852
rect 6604 13812 6610 13824
rect 10888 13728 10916 13824
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 14734 13852 14740 13864
rect 14108 13824 14740 13852
rect 14108 13796 14136 13824
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 18064 13861 18092 13892
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 20717 13923 20775 13929
rect 20717 13889 20729 13923
rect 20763 13889 20775 13923
rect 20898 13920 20904 13932
rect 20859 13892 20904 13920
rect 20717 13883 20775 13889
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 15528 13824 17141 13852
rect 15528 13812 15534 13824
rect 17129 13821 17141 13824
rect 17175 13852 17187 13855
rect 17589 13855 17647 13861
rect 17589 13852 17601 13855
rect 17175 13824 17601 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17589 13821 17601 13824
rect 17635 13821 17647 13855
rect 17589 13815 17647 13821
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18598 13852 18604 13864
rect 18559 13824 18604 13852
rect 18049 13815 18107 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 19610 13812 19616 13864
rect 19668 13852 19674 13864
rect 20732 13852 20760 13883
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 20990 13880 20996 13932
rect 21048 13920 21054 13932
rect 21131 13923 21189 13929
rect 21048 13892 21093 13920
rect 21048 13880 21054 13892
rect 21131 13889 21143 13923
rect 21177 13920 21189 13923
rect 21266 13920 21272 13932
rect 21177 13892 21272 13920
rect 21177 13889 21189 13892
rect 21131 13883 21189 13889
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 21542 13880 21548 13932
rect 21600 13920 21606 13932
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 21600 13892 22385 13920
rect 21600 13880 21606 13892
rect 22373 13889 22385 13892
rect 22419 13920 22431 13923
rect 23155 13923 23213 13929
rect 23155 13920 23167 13923
rect 22419 13892 23167 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 23155 13889 23167 13892
rect 23201 13889 23213 13923
rect 23155 13883 23213 13889
rect 23274 13923 23332 13929
rect 23274 13889 23286 13923
rect 23320 13920 23332 13923
rect 23320 13889 23349 13920
rect 23274 13883 23349 13889
rect 19668 13824 20760 13852
rect 19668 13812 19674 13824
rect 14090 13784 14096 13796
rect 14003 13756 14096 13784
rect 14090 13744 14096 13756
rect 14148 13744 14154 13796
rect 14274 13744 14280 13796
rect 14332 13784 14338 13796
rect 17865 13787 17923 13793
rect 17865 13784 17877 13787
rect 14332 13756 17877 13784
rect 14332 13744 14338 13756
rect 17865 13753 17877 13756
rect 17911 13753 17923 13787
rect 17865 13747 17923 13753
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 18616 13784 18644 13812
rect 18012 13756 18644 13784
rect 23321 13784 23349 13883
rect 23382 13880 23388 13932
rect 23440 13920 23446 13932
rect 23569 13923 23627 13929
rect 23440 13892 23485 13920
rect 23440 13880 23446 13892
rect 23569 13889 23581 13923
rect 23615 13920 23627 13923
rect 23842 13920 23848 13932
rect 23615 13892 23848 13920
rect 23615 13889 23627 13892
rect 23569 13883 23627 13889
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 24118 13880 24124 13932
rect 24176 13920 24182 13932
rect 24397 13923 24455 13929
rect 24397 13920 24409 13923
rect 24176 13892 24409 13920
rect 24176 13880 24182 13892
rect 24397 13889 24409 13892
rect 24443 13920 24455 13923
rect 26973 13923 27031 13929
rect 26973 13920 26985 13923
rect 24443 13892 26985 13920
rect 24443 13889 24455 13892
rect 24397 13883 24455 13889
rect 26973 13889 26985 13892
rect 27019 13889 27031 13923
rect 26973 13883 27031 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 28626 13920 28632 13932
rect 27203 13892 28632 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 28626 13880 28632 13892
rect 28684 13880 28690 13932
rect 28721 13923 28779 13929
rect 28721 13889 28733 13923
rect 28767 13920 28779 13923
rect 30561 13923 30619 13929
rect 30561 13920 30573 13923
rect 28767 13892 30573 13920
rect 28767 13889 28779 13892
rect 28721 13883 28779 13889
rect 30561 13889 30573 13892
rect 30607 13889 30619 13923
rect 30561 13883 30619 13889
rect 28442 13852 28448 13864
rect 28403 13824 28448 13852
rect 28442 13812 28448 13824
rect 28500 13812 28506 13864
rect 30282 13852 30288 13864
rect 30243 13824 30288 13852
rect 30282 13812 30288 13824
rect 30340 13812 30346 13864
rect 30576 13852 30604 13883
rect 30742 13880 30748 13932
rect 30800 13920 30806 13932
rect 31205 13923 31263 13929
rect 31205 13920 31217 13923
rect 30800 13892 31217 13920
rect 30800 13880 30806 13892
rect 31205 13889 31217 13892
rect 31251 13889 31263 13923
rect 31386 13920 31392 13932
rect 31347 13892 31392 13920
rect 31205 13883 31263 13889
rect 31386 13880 31392 13892
rect 31444 13880 31450 13932
rect 31570 13920 31576 13932
rect 31531 13892 31576 13920
rect 31570 13880 31576 13892
rect 31628 13880 31634 13932
rect 33042 13920 33048 13932
rect 33003 13892 33048 13920
rect 33042 13880 33048 13892
rect 33100 13880 33106 13932
rect 33229 13923 33287 13929
rect 33229 13889 33241 13923
rect 33275 13920 33287 13923
rect 33318 13920 33324 13932
rect 33275 13892 33324 13920
rect 33275 13889 33287 13892
rect 33229 13883 33287 13889
rect 33318 13880 33324 13892
rect 33376 13880 33382 13932
rect 33413 13923 33471 13929
rect 33413 13889 33425 13923
rect 33459 13920 33471 13923
rect 33594 13920 33600 13932
rect 33459 13892 33600 13920
rect 33459 13889 33471 13892
rect 33413 13883 33471 13889
rect 33594 13880 33600 13892
rect 33652 13880 33658 13932
rect 34716 13929 34744 13960
rect 36277 13932 36305 13960
rect 36446 13948 36452 13960
rect 36504 13948 36510 14000
rect 34149 13923 34207 13929
rect 34149 13889 34161 13923
rect 34195 13889 34207 13923
rect 34149 13883 34207 13889
rect 34701 13923 34759 13929
rect 34701 13889 34713 13923
rect 34747 13889 34759 13923
rect 34701 13883 34759 13889
rect 30576 13824 32996 13852
rect 23382 13784 23388 13796
rect 23321 13756 23388 13784
rect 18012 13744 18018 13756
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 24302 13744 24308 13796
rect 24360 13784 24366 13796
rect 32858 13784 32864 13796
rect 24360 13756 32864 13784
rect 24360 13744 24366 13756
rect 32858 13744 32864 13756
rect 32916 13744 32922 13796
rect 32968 13784 32996 13824
rect 32968 13756 33180 13784
rect 2700 13688 3096 13716
rect 3513 13719 3571 13725
rect 3513 13685 3525 13719
rect 3559 13716 3571 13719
rect 3878 13716 3884 13728
rect 3559 13688 3884 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 8481 13719 8539 13725
rect 8481 13685 8493 13719
rect 8527 13716 8539 13719
rect 8754 13716 8760 13728
rect 8527 13688 8760 13716
rect 8527 13685 8539 13688
rect 8481 13679 8539 13685
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 10870 13676 10876 13728
rect 10928 13676 10934 13728
rect 12618 13716 12624 13728
rect 12579 13688 12624 13716
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 12802 13716 12808 13728
rect 12763 13688 12808 13716
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 21634 13716 21640 13728
rect 14608 13688 21640 13716
rect 14608 13676 14614 13688
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 23658 13676 23664 13728
rect 23716 13716 23722 13728
rect 24029 13719 24087 13725
rect 24029 13716 24041 13719
rect 23716 13688 24041 13716
rect 23716 13676 23722 13688
rect 24029 13685 24041 13688
rect 24075 13685 24087 13719
rect 24029 13679 24087 13685
rect 27154 13676 27160 13728
rect 27212 13716 27218 13728
rect 27341 13719 27399 13725
rect 27341 13716 27353 13719
rect 27212 13688 27353 13716
rect 27212 13676 27218 13688
rect 27341 13685 27353 13688
rect 27387 13685 27399 13719
rect 27890 13716 27896 13728
rect 27851 13688 27896 13716
rect 27341 13679 27399 13685
rect 27890 13676 27896 13688
rect 27948 13716 27954 13728
rect 28074 13716 28080 13728
rect 27948 13688 28080 13716
rect 27948 13676 27954 13688
rect 28074 13676 28080 13688
rect 28132 13676 28138 13728
rect 31018 13716 31024 13728
rect 30979 13688 31024 13716
rect 31018 13676 31024 13688
rect 31076 13676 31082 13728
rect 33152 13716 33180 13756
rect 34164 13716 34192 13883
rect 34790 13880 34796 13932
rect 34848 13920 34854 13932
rect 34885 13923 34943 13929
rect 34885 13920 34897 13923
rect 34848 13892 34897 13920
rect 34848 13880 34854 13892
rect 34885 13889 34897 13892
rect 34931 13889 34943 13923
rect 34885 13883 34943 13889
rect 34977 13923 35035 13929
rect 34977 13889 34989 13923
rect 35023 13889 35035 13923
rect 34977 13883 35035 13889
rect 34992 13852 35020 13883
rect 35066 13880 35072 13932
rect 35124 13920 35130 13932
rect 35124 13892 35169 13920
rect 35124 13880 35130 13892
rect 35526 13880 35532 13932
rect 35584 13920 35590 13932
rect 36170 13920 36176 13932
rect 35584 13892 36176 13920
rect 35584 13880 35590 13892
rect 36170 13880 36176 13892
rect 36228 13880 36234 13932
rect 36262 13926 36320 13932
rect 36262 13892 36274 13926
rect 36308 13892 36320 13926
rect 36262 13886 36320 13892
rect 35894 13852 35900 13864
rect 34992 13824 35112 13852
rect 35855 13824 35900 13852
rect 35084 13784 35112 13824
rect 35894 13812 35900 13824
rect 35952 13812 35958 13864
rect 36277 13784 36305 13886
rect 36354 13880 36360 13932
rect 36412 13920 36418 13932
rect 36556 13929 36584 14028
rect 39298 14016 39304 14028
rect 39356 14016 39362 14068
rect 39758 14016 39764 14068
rect 39816 14056 39822 14068
rect 40129 14059 40187 14065
rect 40129 14056 40141 14059
rect 39816 14028 40141 14056
rect 39816 14016 39822 14028
rect 40129 14025 40141 14028
rect 40175 14025 40187 14059
rect 40129 14019 40187 14025
rect 39942 13988 39948 14000
rect 39903 13960 39948 13988
rect 39942 13948 39948 13960
rect 40000 13948 40006 14000
rect 36541 13923 36599 13929
rect 36412 13892 36457 13920
rect 36412 13880 36418 13892
rect 36541 13889 36553 13923
rect 36587 13920 36599 13923
rect 39390 13920 39396 13932
rect 36587 13892 39396 13920
rect 36587 13889 36599 13892
rect 36541 13883 36599 13889
rect 39390 13880 39396 13892
rect 39448 13880 39454 13932
rect 39758 13920 39764 13932
rect 39719 13892 39764 13920
rect 39758 13880 39764 13892
rect 39816 13880 39822 13932
rect 39776 13852 39804 13880
rect 35084 13756 36305 13784
rect 36372 13824 39804 13852
rect 34238 13716 34244 13728
rect 33152 13688 34244 13716
rect 34238 13676 34244 13688
rect 34296 13676 34302 13728
rect 35158 13676 35164 13728
rect 35216 13716 35222 13728
rect 35526 13716 35532 13728
rect 35216 13688 35532 13716
rect 35216 13676 35222 13688
rect 35526 13676 35532 13688
rect 35584 13716 35590 13728
rect 36372 13716 36400 13824
rect 35584 13688 36400 13716
rect 35584 13676 35590 13688
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 1946 13512 1952 13524
rect 1907 13484 1952 13512
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 11422 13512 11428 13524
rect 10919 13484 11428 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 11422 13472 11428 13484
rect 11480 13512 11486 13524
rect 17313 13515 17371 13521
rect 17313 13512 17325 13515
rect 11480 13484 17325 13512
rect 11480 13472 11486 13484
rect 17313 13481 17325 13484
rect 17359 13481 17371 13515
rect 17313 13475 17371 13481
rect 2682 13444 2688 13456
rect 2424 13416 2688 13444
rect 2424 13385 2452 13416
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 12066 13444 12072 13456
rect 6503 13416 12072 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13345 2467 13379
rect 2409 13339 2467 13345
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 5077 13379 5135 13385
rect 5077 13376 5089 13379
rect 4120 13348 5089 13376
rect 4120 13336 4126 13348
rect 5077 13345 5089 13348
rect 5123 13345 5135 13379
rect 5077 13339 5135 13345
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 2590 13268 2596 13320
rect 2648 13308 2654 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2648 13280 2697 13308
rect 2648 13268 2654 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 5333 13311 5391 13317
rect 5333 13308 5345 13311
rect 4672 13280 5345 13308
rect 4672 13268 4678 13280
rect 5333 13277 5345 13280
rect 5379 13277 5391 13311
rect 5333 13271 5391 13277
rect 1765 13243 1823 13249
rect 1765 13209 1777 13243
rect 1811 13209 1823 13243
rect 1765 13203 1823 13209
rect 1780 13172 1808 13203
rect 6472 13172 6500 13407
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 13449 13447 13507 13453
rect 13449 13413 13461 13447
rect 13495 13444 13507 13447
rect 14274 13444 14280 13456
rect 13495 13416 14280 13444
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 14274 13404 14280 13416
rect 14332 13404 14338 13456
rect 17328 13444 17356 13475
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 21082 13512 21088 13524
rect 17460 13484 21088 13512
rect 17460 13472 17466 13484
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 21361 13515 21419 13521
rect 21361 13512 21373 13515
rect 21232 13484 21373 13512
rect 21232 13472 21238 13484
rect 21361 13481 21373 13484
rect 21407 13481 21419 13515
rect 21361 13475 21419 13481
rect 21634 13472 21640 13524
rect 21692 13512 21698 13524
rect 21692 13484 22048 13512
rect 21692 13472 21698 13484
rect 17328 13416 18736 13444
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8352 13348 8953 13376
rect 8352 13336 8358 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 11572 13348 11621 13376
rect 11572 13336 11578 13348
rect 11609 13345 11621 13348
rect 11655 13345 11667 13379
rect 11609 13339 11667 13345
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13136 13348 13553 13376
rect 13136 13336 13142 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 14056 13348 14105 13376
rect 14056 13336 14062 13348
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 14550 13376 14556 13388
rect 14511 13348 14556 13376
rect 14093 13339 14151 13345
rect 14550 13336 14556 13348
rect 14608 13336 14614 13388
rect 15378 13376 15384 13388
rect 15339 13348 15384 13376
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 18708 13385 18736 13416
rect 21450 13404 21456 13456
rect 21508 13444 21514 13456
rect 21821 13447 21879 13453
rect 21821 13444 21833 13447
rect 21508 13416 21833 13444
rect 21508 13404 21514 13416
rect 21821 13413 21833 13416
rect 21867 13413 21879 13447
rect 21821 13407 21879 13413
rect 18693 13379 18751 13385
rect 18693 13345 18705 13379
rect 18739 13345 18751 13379
rect 18693 13339 18751 13345
rect 18874 13336 18880 13388
rect 18932 13376 18938 13388
rect 20530 13376 20536 13388
rect 18932 13348 20536 13376
rect 18932 13336 18938 13348
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 21266 13376 21272 13388
rect 21179 13348 21272 13376
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7926 13308 7932 13320
rect 7147 13280 7932 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 9217 13311 9275 13317
rect 9217 13308 9229 13311
rect 8312 13280 9229 13308
rect 8312 13252 8340 13280
rect 9217 13277 9229 13280
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 10781 13311 10839 13317
rect 10781 13308 10793 13311
rect 10192 13280 10793 13308
rect 10192 13268 10198 13280
rect 10781 13277 10793 13280
rect 10827 13308 10839 13311
rect 10962 13308 10968 13320
rect 10827 13280 10968 13308
rect 10827 13277 10839 13280
rect 10781 13271 10839 13277
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11698 13268 11704 13320
rect 11756 13308 11762 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11756 13280 11897 13308
rect 11756 13268 11762 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 18414 13308 18420 13320
rect 18375 13280 18420 13308
rect 11885 13271 11943 13277
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 21192 13317 21220 13348
rect 21266 13336 21272 13348
rect 21324 13376 21330 13388
rect 21910 13376 21916 13388
rect 21324 13348 21916 13376
rect 21324 13336 21330 13348
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19392 13280 19625 13308
rect 19392 13268 19398 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21177 13311 21235 13317
rect 21177 13277 21189 13311
rect 21223 13277 21235 13311
rect 21177 13271 21235 13277
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13240 7343 13243
rect 8018 13240 8024 13252
rect 7331 13212 8024 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 8205 13243 8263 13249
rect 8205 13209 8217 13243
rect 8251 13209 8263 13243
rect 8205 13203 8263 13209
rect 6914 13172 6920 13184
rect 1780 13144 6500 13172
rect 6875 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 8220 13172 8248 13203
rect 8294 13200 8300 13252
rect 8352 13200 8358 13252
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 8444 13212 8489 13240
rect 8444 13200 8450 13212
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 13081 13243 13139 13249
rect 13081 13240 13093 13243
rect 11112 13212 13093 13240
rect 11112 13200 11118 13212
rect 13081 13209 13093 13212
rect 13127 13209 13139 13243
rect 13081 13203 13139 13209
rect 15648 13243 15706 13249
rect 15648 13209 15660 13243
rect 15694 13240 15706 13243
rect 17586 13240 17592 13252
rect 15694 13212 17592 13240
rect 15694 13209 15706 13212
rect 15648 13203 15706 13209
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 19429 13243 19487 13249
rect 19429 13240 19441 13243
rect 17972 13212 19441 13240
rect 9858 13172 9864 13184
rect 8220 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 16761 13175 16819 13181
rect 16761 13141 16773 13175
rect 16807 13172 16819 13175
rect 17972 13172 18000 13212
rect 19429 13209 19441 13212
rect 19475 13240 19487 13243
rect 20824 13240 20852 13271
rect 21726 13268 21732 13320
rect 21784 13308 21790 13320
rect 22020 13317 22048 13484
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 22649 13515 22707 13521
rect 22649 13512 22661 13515
rect 22612 13484 22661 13512
rect 22612 13472 22618 13484
rect 22649 13481 22661 13484
rect 22695 13481 22707 13515
rect 22649 13475 22707 13481
rect 21821 13311 21879 13317
rect 21821 13308 21833 13311
rect 21784 13280 21833 13308
rect 21784 13268 21790 13280
rect 21821 13277 21833 13280
rect 21867 13277 21879 13311
rect 21821 13271 21879 13277
rect 22005 13311 22063 13317
rect 22005 13277 22017 13311
rect 22051 13277 22063 13311
rect 22664 13308 22692 13475
rect 23014 13472 23020 13524
rect 23072 13512 23078 13524
rect 23201 13515 23259 13521
rect 23201 13512 23213 13515
rect 23072 13484 23213 13512
rect 23072 13472 23078 13484
rect 23201 13481 23213 13484
rect 23247 13481 23259 13515
rect 23201 13475 23259 13481
rect 28626 13472 28632 13524
rect 28684 13512 28690 13524
rect 28905 13515 28963 13521
rect 28905 13512 28917 13515
rect 28684 13484 28917 13512
rect 28684 13472 28690 13484
rect 28905 13481 28917 13484
rect 28951 13481 28963 13515
rect 32858 13512 32864 13524
rect 32819 13484 32864 13512
rect 28905 13475 28963 13481
rect 32858 13472 32864 13484
rect 32916 13472 32922 13524
rect 34149 13515 34207 13521
rect 34149 13481 34161 13515
rect 34195 13512 34207 13515
rect 34195 13484 34928 13512
rect 34195 13481 34207 13484
rect 34149 13475 34207 13481
rect 34900 13456 34928 13484
rect 35802 13472 35808 13524
rect 35860 13512 35866 13524
rect 37553 13515 37611 13521
rect 37553 13512 37565 13515
rect 35860 13484 37565 13512
rect 35860 13472 35866 13484
rect 37553 13481 37565 13484
rect 37599 13512 37611 13515
rect 37599 13484 41276 13512
rect 37599 13481 37611 13484
rect 37553 13475 37611 13481
rect 22738 13404 22744 13456
rect 22796 13444 22802 13456
rect 25498 13444 25504 13456
rect 22796 13416 25504 13444
rect 22796 13404 22802 13416
rect 25498 13404 25504 13416
rect 25556 13404 25562 13456
rect 29822 13404 29828 13456
rect 29880 13444 29886 13456
rect 30282 13444 30288 13456
rect 29880 13416 30288 13444
rect 29880 13404 29886 13416
rect 30282 13404 30288 13416
rect 30340 13444 30346 13456
rect 31846 13444 31852 13456
rect 30340 13416 31852 13444
rect 30340 13404 30346 13416
rect 23382 13336 23388 13388
rect 23440 13376 23446 13388
rect 26786 13376 26792 13388
rect 23440 13348 23612 13376
rect 26747 13348 26792 13376
rect 23440 13336 23446 13348
rect 23584 13317 23612 13348
rect 26786 13336 26792 13348
rect 26844 13376 26850 13388
rect 27525 13379 27583 13385
rect 27525 13376 27537 13379
rect 26844 13348 27537 13376
rect 26844 13336 26850 13348
rect 27525 13345 27537 13348
rect 27571 13345 27583 13379
rect 27525 13339 27583 13345
rect 29638 13336 29644 13388
rect 29696 13376 29702 13388
rect 31036 13385 31064 13416
rect 31846 13404 31852 13416
rect 31904 13444 31910 13456
rect 32306 13444 32312 13456
rect 31904 13416 32312 13444
rect 31904 13404 31910 13416
rect 32306 13404 32312 13416
rect 32364 13404 32370 13456
rect 32401 13447 32459 13453
rect 32401 13413 32413 13447
rect 32447 13444 32459 13447
rect 32582 13444 32588 13456
rect 32447 13416 32588 13444
rect 32447 13413 32459 13416
rect 32401 13407 32459 13413
rect 32582 13404 32588 13416
rect 32640 13444 32646 13456
rect 33410 13444 33416 13456
rect 32640 13416 33416 13444
rect 32640 13404 32646 13416
rect 33410 13404 33416 13416
rect 33468 13444 33474 13456
rect 34701 13447 34759 13453
rect 34701 13444 34713 13447
rect 33468 13416 34713 13444
rect 33468 13404 33474 13416
rect 34701 13413 34713 13416
rect 34747 13444 34759 13447
rect 34790 13444 34796 13456
rect 34747 13416 34796 13444
rect 34747 13413 34759 13416
rect 34701 13407 34759 13413
rect 34790 13404 34796 13416
rect 34848 13404 34854 13456
rect 34882 13404 34888 13456
rect 34940 13444 34946 13456
rect 36170 13444 36176 13456
rect 34940 13416 36176 13444
rect 34940 13404 34946 13416
rect 36170 13404 36176 13416
rect 36228 13404 36234 13456
rect 40126 13404 40132 13456
rect 40184 13444 40190 13456
rect 40184 13416 40264 13444
rect 40184 13404 40190 13416
rect 31021 13379 31079 13385
rect 29696 13348 30328 13376
rect 29696 13336 29702 13348
rect 23477 13311 23535 13317
rect 23477 13308 23489 13311
rect 22664 13280 23489 13308
rect 22005 13271 22063 13277
rect 23477 13277 23489 13280
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 23658 13268 23664 13320
rect 23716 13308 23722 13320
rect 23716 13280 23761 13308
rect 23716 13268 23722 13280
rect 23842 13268 23848 13320
rect 23900 13308 23906 13320
rect 25038 13308 25044 13320
rect 23900 13280 25044 13308
rect 23900 13268 23906 13280
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 29822 13268 29828 13320
rect 29880 13308 29886 13320
rect 30300 13317 30328 13348
rect 31021 13345 31033 13379
rect 31067 13345 31079 13379
rect 35621 13379 35679 13385
rect 31021 13339 31079 13345
rect 33336 13348 35480 13376
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 29880 13280 29929 13308
rect 29880 13268 29886 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 30285 13311 30343 13317
rect 30285 13277 30297 13311
rect 30331 13277 30343 13311
rect 30285 13271 30343 13277
rect 30466 13268 30472 13320
rect 30524 13308 30530 13320
rect 30742 13308 30748 13320
rect 30524 13280 30748 13308
rect 30524 13268 30530 13280
rect 30742 13268 30748 13280
rect 30800 13268 30806 13320
rect 33042 13308 33048 13320
rect 33003 13280 33048 13308
rect 33042 13268 33048 13280
rect 33100 13268 33106 13320
rect 33137 13311 33195 13317
rect 33137 13277 33149 13311
rect 33183 13308 33195 13311
rect 33336 13308 33364 13348
rect 35452 13317 35480 13348
rect 35621 13345 35633 13379
rect 35667 13376 35679 13379
rect 36354 13376 36360 13388
rect 35667 13348 36360 13376
rect 35667 13345 35679 13348
rect 35621 13339 35679 13345
rect 36354 13336 36360 13348
rect 36412 13336 36418 13388
rect 38933 13379 38991 13385
rect 38933 13345 38945 13379
rect 38979 13376 38991 13379
rect 39114 13376 39120 13388
rect 38979 13348 39120 13376
rect 38979 13345 38991 13348
rect 38933 13339 38991 13345
rect 39114 13336 39120 13348
rect 39172 13336 39178 13388
rect 33183 13280 33364 13308
rect 33413 13311 33471 13317
rect 33183 13277 33195 13280
rect 33137 13271 33195 13277
rect 33413 13277 33425 13311
rect 33459 13277 33471 13311
rect 33413 13271 33471 13277
rect 35437 13311 35495 13317
rect 35437 13277 35449 13311
rect 35483 13308 35495 13311
rect 35710 13308 35716 13320
rect 35483 13280 35716 13308
rect 35483 13277 35495 13280
rect 35437 13271 35495 13277
rect 20990 13240 20996 13252
rect 19475 13212 20852 13240
rect 20951 13212 20996 13240
rect 19475 13209 19487 13212
rect 19429 13203 19487 13209
rect 20990 13200 20996 13212
rect 21048 13200 21054 13252
rect 21085 13243 21143 13249
rect 21085 13209 21097 13243
rect 21131 13240 21143 13243
rect 23934 13240 23940 13252
rect 21131 13212 23940 13240
rect 21131 13209 21143 13212
rect 21085 13203 21143 13209
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 24118 13200 24124 13252
rect 24176 13240 24182 13252
rect 24581 13243 24639 13249
rect 24581 13240 24593 13243
rect 24176 13212 24593 13240
rect 24176 13200 24182 13212
rect 24581 13209 24593 13212
rect 24627 13240 24639 13243
rect 24670 13240 24676 13252
rect 24627 13212 24676 13240
rect 24627 13209 24639 13212
rect 24581 13203 24639 13209
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 24765 13243 24823 13249
rect 24765 13209 24777 13243
rect 24811 13240 24823 13243
rect 24811 13212 25452 13240
rect 24811 13209 24823 13212
rect 24765 13203 24823 13209
rect 16807 13144 18000 13172
rect 16807 13141 16819 13144
rect 16761 13135 16819 13141
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 18104 13144 19257 13172
rect 18104 13132 18110 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 24026 13132 24032 13184
rect 24084 13172 24090 13184
rect 24780 13172 24808 13203
rect 24946 13172 24952 13184
rect 24084 13144 24808 13172
rect 24907 13144 24952 13172
rect 24084 13132 24090 13144
rect 24946 13132 24952 13144
rect 25004 13132 25010 13184
rect 25424 13181 25452 13212
rect 25682 13200 25688 13252
rect 25740 13240 25746 13252
rect 26522 13243 26580 13249
rect 26522 13240 26534 13243
rect 25740 13212 26534 13240
rect 25740 13200 25746 13212
rect 26522 13209 26534 13212
rect 26568 13209 26580 13243
rect 26522 13203 26580 13209
rect 27614 13200 27620 13252
rect 27672 13240 27678 13252
rect 27770 13243 27828 13249
rect 27770 13240 27782 13243
rect 27672 13212 27782 13240
rect 27672 13200 27678 13212
rect 27770 13209 27782 13212
rect 27816 13209 27828 13243
rect 30006 13240 30012 13252
rect 29967 13212 30012 13240
rect 27770 13203 27828 13209
rect 30006 13200 30012 13212
rect 30064 13200 30070 13252
rect 30101 13243 30159 13249
rect 30101 13209 30113 13243
rect 30147 13240 30159 13243
rect 30374 13240 30380 13252
rect 30147 13212 30380 13240
rect 30147 13209 30159 13212
rect 30101 13203 30159 13209
rect 30374 13200 30380 13212
rect 30432 13200 30438 13252
rect 33229 13243 33287 13249
rect 33229 13209 33241 13243
rect 33275 13240 33287 13243
rect 33318 13240 33324 13252
rect 33275 13212 33324 13240
rect 33275 13209 33287 13212
rect 33229 13203 33287 13209
rect 33318 13200 33324 13212
rect 33376 13200 33382 13252
rect 25409 13175 25467 13181
rect 25409 13141 25421 13175
rect 25455 13141 25467 13175
rect 25409 13135 25467 13141
rect 29733 13175 29791 13181
rect 29733 13141 29745 13175
rect 29779 13172 29791 13175
rect 29822 13172 29828 13184
rect 29779 13144 29828 13172
rect 29779 13141 29791 13144
rect 29733 13135 29791 13141
rect 29822 13132 29828 13144
rect 29880 13132 29886 13184
rect 33042 13132 33048 13184
rect 33100 13172 33106 13184
rect 33428 13172 33456 13271
rect 35710 13268 35716 13280
rect 35768 13268 35774 13320
rect 39298 13268 39304 13320
rect 39356 13308 39362 13320
rect 40236 13317 40264 13416
rect 40328 13348 41092 13376
rect 40328 13317 40356 13348
rect 40129 13311 40187 13317
rect 40129 13308 40141 13311
rect 39356 13280 40141 13308
rect 39356 13268 39362 13280
rect 40129 13277 40141 13280
rect 40175 13277 40187 13311
rect 40129 13271 40187 13277
rect 40221 13311 40279 13317
rect 40221 13277 40233 13311
rect 40267 13277 40279 13311
rect 40221 13271 40279 13277
rect 40313 13311 40371 13317
rect 40313 13277 40325 13311
rect 40359 13277 40371 13311
rect 40313 13271 40371 13277
rect 40494 13268 40500 13320
rect 40552 13308 40558 13320
rect 40552 13280 40597 13308
rect 40552 13268 40558 13280
rect 34698 13200 34704 13252
rect 34756 13240 34762 13252
rect 35253 13243 35311 13249
rect 35253 13240 35265 13243
rect 34756 13212 35265 13240
rect 34756 13200 34762 13212
rect 35253 13209 35265 13212
rect 35299 13240 35311 13243
rect 35526 13240 35532 13252
rect 35299 13212 35532 13240
rect 35299 13209 35311 13212
rect 35253 13203 35311 13209
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 38688 13243 38746 13249
rect 38688 13209 38700 13243
rect 38734 13240 38746 13243
rect 39853 13243 39911 13249
rect 39853 13240 39865 13243
rect 38734 13212 39865 13240
rect 38734 13209 38746 13212
rect 38688 13203 38746 13209
rect 39853 13209 39865 13212
rect 39899 13209 39911 13243
rect 39853 13203 39911 13209
rect 39942 13200 39948 13252
rect 40000 13240 40006 13252
rect 40957 13243 41015 13249
rect 40957 13240 40969 13243
rect 40000 13212 40969 13240
rect 40000 13200 40006 13212
rect 40957 13209 40969 13212
rect 41003 13209 41015 13243
rect 41064 13240 41092 13348
rect 41141 13311 41199 13317
rect 41141 13277 41153 13311
rect 41187 13308 41199 13311
rect 41248 13308 41276 13484
rect 68094 13308 68100 13320
rect 41187 13280 41276 13308
rect 68055 13280 68100 13308
rect 41187 13277 41199 13280
rect 41141 13271 41199 13277
rect 68094 13268 68100 13280
rect 68152 13268 68158 13320
rect 41325 13243 41383 13249
rect 41325 13240 41337 13243
rect 41064 13212 41337 13240
rect 40957 13203 41015 13209
rect 41325 13209 41337 13212
rect 41371 13209 41383 13243
rect 41325 13203 41383 13209
rect 33100 13144 33456 13172
rect 33100 13132 33106 13144
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 4062 12928 4068 12980
rect 4120 12928 4126 12980
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 5721 12971 5779 12977
rect 5721 12968 5733 12971
rect 5408 12940 5733 12968
rect 5408 12928 5414 12940
rect 5721 12937 5733 12940
rect 5767 12937 5779 12971
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 5721 12931 5779 12937
rect 4080 12900 4108 12928
rect 3804 12872 4108 12900
rect 3804 12844 3832 12872
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2314 12832 2320 12844
rect 1995 12804 2320 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2314 12792 2320 12804
rect 2372 12832 2378 12844
rect 2685 12835 2743 12841
rect 2685 12832 2697 12835
rect 2372 12804 2697 12832
rect 2372 12792 2378 12804
rect 2685 12801 2697 12804
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12801 2927 12835
rect 3786 12832 3792 12844
rect 3699 12804 3792 12832
rect 2869 12795 2927 12801
rect 1394 12588 1400 12640
rect 1452 12628 1458 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 1452 12600 2145 12628
rect 1452 12588 1458 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 2884 12628 2912 12795
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4045 12835 4103 12841
rect 4045 12832 4057 12835
rect 3936 12804 4057 12832
rect 3936 12792 3942 12804
rect 4045 12801 4057 12804
rect 4091 12801 4103 12835
rect 5736 12832 5764 12931
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 9858 12968 9864 12980
rect 9819 12940 9864 12968
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10413 12971 10471 12977
rect 10413 12937 10425 12971
rect 10459 12968 10471 12971
rect 12158 12968 12164 12980
rect 10459 12940 12164 12968
rect 10459 12937 10471 12940
rect 10413 12931 10471 12937
rect 12158 12928 12164 12940
rect 12216 12968 12222 12980
rect 13265 12971 13323 12977
rect 12216 12940 12434 12968
rect 12216 12928 12222 12940
rect 8294 12900 8300 12912
rect 6840 12872 8300 12900
rect 6840 12841 6868 12872
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 9674 12900 9680 12912
rect 8680 12872 9680 12900
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 5736 12804 6745 12832
rect 4045 12795 4103 12801
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7101 12835 7159 12841
rect 6972 12804 7017 12832
rect 6972 12792 6978 12804
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 7190 12832 7196 12844
rect 7147 12804 7196 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 8110 12832 8116 12844
rect 7883 12804 8116 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8110 12792 8116 12804
rect 8168 12832 8174 12844
rect 8386 12832 8392 12844
rect 8168 12804 8392 12832
rect 8168 12792 8174 12804
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12832 8539 12835
rect 8680 12832 8708 12872
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 10965 12903 11023 12909
rect 10965 12869 10977 12903
rect 11011 12900 11023 12903
rect 11054 12900 11060 12912
rect 11011 12872 11060 12900
rect 11011 12869 11023 12872
rect 10965 12863 11023 12869
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 11977 12903 12035 12909
rect 11977 12900 11989 12903
rect 11756 12872 11989 12900
rect 11756 12860 11762 12872
rect 11977 12869 11989 12872
rect 12023 12869 12035 12903
rect 11977 12863 12035 12869
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12124 12872 12169 12900
rect 12124 12860 12130 12872
rect 8754 12841 8760 12844
rect 8527 12804 8708 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 8748 12795 8760 12841
rect 8812 12832 8818 12844
rect 11790 12832 11796 12844
rect 8812 12804 8848 12832
rect 11751 12804 11796 12832
rect 8754 12792 8760 12795
rect 8812 12792 8818 12804
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 11882 12724 11888 12776
rect 11940 12764 11946 12776
rect 12176 12764 12204 12795
rect 11940 12736 12204 12764
rect 12406 12764 12434 12940
rect 13265 12937 13277 12971
rect 13311 12968 13323 12971
rect 13354 12968 13360 12980
rect 13311 12940 13360 12968
rect 13311 12937 13323 12940
rect 13265 12931 13323 12937
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 15102 12968 15108 12980
rect 15063 12940 15108 12968
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 17126 12968 17132 12980
rect 17087 12940 17132 12968
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 17586 12968 17592 12980
rect 17547 12940 17592 12968
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 18966 12968 18972 12980
rect 18927 12940 18972 12968
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 21634 12968 21640 12980
rect 21232 12940 21640 12968
rect 21232 12928 21238 12940
rect 21634 12928 21640 12940
rect 21692 12968 21698 12980
rect 21821 12971 21879 12977
rect 21821 12968 21833 12971
rect 21692 12940 21833 12968
rect 21692 12928 21698 12940
rect 21821 12937 21833 12940
rect 21867 12937 21879 12971
rect 21821 12931 21879 12937
rect 24305 12971 24363 12977
rect 24305 12937 24317 12971
rect 24351 12968 24363 12971
rect 24486 12968 24492 12980
rect 24351 12940 24492 12968
rect 24351 12937 24363 12940
rect 24305 12931 24363 12937
rect 24486 12928 24492 12940
rect 24544 12928 24550 12980
rect 25682 12968 25688 12980
rect 25643 12940 25688 12968
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 25774 12928 25780 12980
rect 25832 12968 25838 12980
rect 27614 12968 27620 12980
rect 25832 12940 26234 12968
rect 27575 12940 27620 12968
rect 25832 12928 25838 12940
rect 15654 12860 15660 12912
rect 15712 12900 15718 12912
rect 17678 12900 17684 12912
rect 15712 12872 17684 12900
rect 15712 12860 15718 12872
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 18598 12860 18604 12912
rect 18656 12900 18662 12912
rect 20898 12900 20904 12912
rect 18656 12872 20904 12900
rect 18656 12860 18662 12872
rect 20898 12860 20904 12872
rect 20956 12900 20962 12912
rect 21269 12903 21327 12909
rect 21269 12900 21281 12903
rect 20956 12872 21281 12900
rect 20956 12860 20962 12872
rect 21269 12869 21281 12872
rect 21315 12900 21327 12903
rect 22002 12900 22008 12912
rect 21315 12872 22008 12900
rect 21315 12869 21327 12872
rect 21269 12863 21327 12869
rect 22002 12860 22008 12872
rect 22060 12860 22066 12912
rect 24026 12900 24032 12912
rect 23987 12872 24032 12900
rect 24026 12860 24032 12872
rect 24084 12860 24090 12912
rect 24946 12860 24952 12912
rect 25004 12900 25010 12912
rect 25004 12872 25176 12900
rect 25004 12860 25010 12872
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12801 13139 12835
rect 13262 12832 13268 12844
rect 13223 12804 13268 12832
rect 13081 12795 13139 12801
rect 13096 12764 13124 12795
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 14642 12832 14648 12844
rect 14599 12804 14648 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12832 15439 12835
rect 15470 12832 15476 12844
rect 15427 12804 15476 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 14458 12764 14464 12776
rect 12406 12736 13124 12764
rect 14419 12736 14464 12764
rect 11940 12724 11946 12736
rect 5169 12699 5227 12705
rect 5169 12665 5181 12699
rect 5215 12696 5227 12699
rect 12342 12696 12348 12708
rect 5215 12668 6776 12696
rect 12303 12668 12348 12696
rect 5215 12665 5227 12668
rect 5169 12659 5227 12665
rect 5184 12628 5212 12659
rect 2884 12600 5212 12628
rect 6457 12631 6515 12637
rect 2133 12591 2191 12597
rect 6457 12597 6469 12631
rect 6503 12628 6515 12631
rect 6638 12628 6644 12640
rect 6503 12600 6644 12628
rect 6503 12597 6515 12600
rect 6457 12591 6515 12597
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 6748 12628 6776 12668
rect 12342 12656 12348 12668
rect 12400 12656 12406 12708
rect 13096 12696 13124 12736
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 14550 12696 14556 12708
rect 13096 12668 14556 12696
rect 14550 12656 14556 12668
rect 14608 12656 14614 12708
rect 10594 12628 10600 12640
rect 6748 12600 10600 12628
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 12986 12628 12992 12640
rect 11296 12600 12992 12628
rect 11296 12588 11302 12600
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14274 12628 14280 12640
rect 14231 12600 14280 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 15212 12628 15240 12795
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 17862 12832 17868 12844
rect 17823 12804 17868 12832
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12801 18015 12835
rect 17957 12795 18015 12801
rect 17972 12764 18000 12795
rect 18046 12792 18052 12844
rect 18104 12832 18110 12844
rect 18104 12804 18149 12832
rect 18104 12792 18110 12804
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 18414 12832 18420 12844
rect 18288 12804 18420 12832
rect 18288 12792 18294 12804
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18966 12792 18972 12844
rect 19024 12832 19030 12844
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 19024 12804 19533 12832
rect 19024 12792 19030 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 20530 12792 20536 12844
rect 20588 12832 20594 12844
rect 22278 12832 22284 12844
rect 20588 12804 22284 12832
rect 20588 12792 20594 12804
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 23753 12835 23811 12841
rect 23753 12832 23765 12835
rect 23676 12804 23765 12832
rect 18322 12764 18328 12776
rect 17972 12736 18328 12764
rect 18322 12724 18328 12736
rect 18380 12724 18386 12776
rect 22186 12764 22192 12776
rect 19720 12736 22192 12764
rect 15286 12656 15292 12708
rect 15344 12696 15350 12708
rect 15933 12699 15991 12705
rect 15933 12696 15945 12699
rect 15344 12668 15945 12696
rect 15344 12656 15350 12668
rect 15933 12665 15945 12668
rect 15979 12696 15991 12699
rect 15979 12668 17632 12696
rect 15979 12665 15991 12668
rect 15933 12659 15991 12665
rect 15378 12628 15384 12640
rect 14424 12600 14469 12628
rect 15212 12600 15384 12628
rect 14424 12588 14430 12600
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 17604 12628 17632 12668
rect 19720 12628 19748 12736
rect 22186 12724 22192 12736
rect 22244 12764 22250 12776
rect 22738 12764 22744 12776
rect 22244 12736 22744 12764
rect 22244 12724 22250 12736
rect 22738 12724 22744 12736
rect 22796 12724 22802 12776
rect 22646 12628 22652 12640
rect 17604 12600 19748 12628
rect 22607 12600 22652 12628
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 23106 12588 23112 12640
rect 23164 12628 23170 12640
rect 23676 12628 23704 12804
rect 23753 12801 23765 12804
rect 23799 12801 23811 12835
rect 23753 12795 23811 12801
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 25038 12832 25044 12844
rect 24999 12804 25044 12832
rect 24121 12795 24179 12801
rect 23952 12764 23980 12795
rect 24026 12764 24032 12776
rect 23952 12736 24032 12764
rect 24026 12724 24032 12736
rect 24084 12724 24090 12776
rect 23934 12656 23940 12708
rect 23992 12696 23998 12708
rect 24136 12696 24164 12795
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25148 12832 25176 12872
rect 25204 12835 25262 12841
rect 25204 12832 25216 12835
rect 25148 12804 25216 12832
rect 25204 12801 25216 12804
rect 25250 12801 25262 12835
rect 25204 12795 25262 12801
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 24946 12724 24952 12776
rect 25004 12764 25010 12776
rect 25331 12764 25359 12795
rect 25426 12792 25432 12844
rect 25484 12841 25490 12844
rect 25484 12835 25513 12841
rect 25501 12801 25513 12835
rect 25484 12795 25513 12801
rect 25484 12792 25490 12795
rect 25004 12736 25359 12764
rect 26206 12764 26234 12940
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 31846 12928 31852 12980
rect 31904 12968 31910 12980
rect 37458 12968 37464 12980
rect 31904 12940 37464 12968
rect 31904 12928 31910 12940
rect 37458 12928 37464 12940
rect 37516 12928 37522 12980
rect 30374 12860 30380 12912
rect 30432 12900 30438 12912
rect 31389 12903 31447 12909
rect 31389 12900 31401 12903
rect 30432 12872 31401 12900
rect 30432 12860 30438 12872
rect 31389 12869 31401 12872
rect 31435 12900 31447 12903
rect 32493 12903 32551 12909
rect 32493 12900 32505 12903
rect 31435 12872 32505 12900
rect 31435 12869 31447 12872
rect 31389 12863 31447 12869
rect 32493 12869 32505 12872
rect 32539 12869 32551 12903
rect 32493 12863 32551 12869
rect 32600 12872 32996 12900
rect 26970 12832 26976 12844
rect 26931 12804 26976 12832
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27154 12841 27160 12844
rect 27152 12832 27160 12841
rect 27115 12804 27160 12832
rect 27152 12795 27160 12804
rect 27154 12792 27160 12795
rect 27212 12792 27218 12844
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 27387 12835 27445 12841
rect 27304 12804 27349 12832
rect 27304 12792 27310 12804
rect 27387 12801 27399 12835
rect 27433 12801 27445 12835
rect 27387 12795 27445 12801
rect 28445 12835 28503 12841
rect 28445 12801 28457 12835
rect 28491 12832 28503 12835
rect 28626 12832 28632 12844
rect 28491 12804 28632 12832
rect 28491 12801 28503 12804
rect 28445 12795 28503 12801
rect 26421 12767 26479 12773
rect 26421 12764 26433 12767
rect 26206 12736 26433 12764
rect 25004 12724 25010 12736
rect 26421 12733 26433 12736
rect 26467 12764 26479 12767
rect 27402 12764 27430 12795
rect 28626 12792 28632 12804
rect 28684 12832 28690 12844
rect 28997 12835 29055 12841
rect 28997 12832 29009 12835
rect 28684 12804 29009 12832
rect 28684 12792 28690 12804
rect 28997 12801 29009 12804
rect 29043 12801 29055 12835
rect 28997 12795 29055 12801
rect 30282 12792 30288 12844
rect 30340 12832 30346 12844
rect 31205 12835 31263 12841
rect 31205 12832 31217 12835
rect 30340 12804 31217 12832
rect 30340 12792 30346 12804
rect 31205 12801 31217 12804
rect 31251 12801 31263 12835
rect 31205 12795 31263 12801
rect 31297 12835 31355 12841
rect 31297 12801 31309 12835
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 31573 12835 31631 12841
rect 31573 12801 31585 12835
rect 31619 12832 31631 12835
rect 32306 12832 32312 12844
rect 31619 12804 31892 12832
rect 32267 12804 32312 12832
rect 31619 12801 31631 12804
rect 31573 12795 31631 12801
rect 26467 12736 27430 12764
rect 26467 12733 26479 12736
rect 26421 12727 26479 12733
rect 27522 12724 27528 12776
rect 27580 12764 27586 12776
rect 29638 12764 29644 12776
rect 27580 12736 29644 12764
rect 27580 12724 27586 12736
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 23992 12668 24164 12696
rect 23992 12656 23998 12668
rect 24670 12656 24676 12708
rect 24728 12696 24734 12708
rect 26142 12696 26148 12708
rect 24728 12668 26148 12696
rect 24728 12656 24734 12668
rect 26142 12656 26148 12668
rect 26200 12656 26206 12708
rect 31312 12696 31340 12795
rect 31754 12696 31760 12708
rect 31312 12668 31760 12696
rect 31754 12656 31760 12668
rect 31812 12656 31818 12708
rect 31864 12696 31892 12804
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 32401 12835 32459 12841
rect 32401 12801 32413 12835
rect 32447 12832 32459 12835
rect 32600 12832 32628 12872
rect 32447 12804 32628 12832
rect 32677 12835 32735 12841
rect 32447 12801 32459 12804
rect 32401 12795 32459 12801
rect 32677 12801 32689 12835
rect 32723 12801 32735 12835
rect 32677 12795 32735 12801
rect 31938 12724 31944 12776
rect 31996 12764 32002 12776
rect 32692 12764 32720 12795
rect 31996 12736 32720 12764
rect 31996 12724 32002 12736
rect 32766 12696 32772 12708
rect 31864 12668 32772 12696
rect 32766 12656 32772 12668
rect 32824 12656 32830 12708
rect 29086 12628 29092 12640
rect 23164 12600 23704 12628
rect 29047 12600 29092 12628
rect 23164 12588 23170 12600
rect 29086 12588 29092 12600
rect 29144 12588 29150 12640
rect 30374 12588 30380 12640
rect 30432 12628 30438 12640
rect 31021 12631 31079 12637
rect 31021 12628 31033 12631
rect 30432 12600 31033 12628
rect 30432 12588 30438 12600
rect 31021 12597 31033 12600
rect 31067 12597 31079 12631
rect 31021 12591 31079 12597
rect 31386 12588 31392 12640
rect 31444 12628 31450 12640
rect 32125 12631 32183 12637
rect 32125 12628 32137 12631
rect 31444 12600 32137 12628
rect 31444 12588 31450 12600
rect 32125 12597 32137 12600
rect 32171 12597 32183 12631
rect 32968 12628 32996 12872
rect 34238 12860 34244 12912
rect 34296 12900 34302 12912
rect 39025 12903 39083 12909
rect 39025 12900 39037 12903
rect 34296 12872 39037 12900
rect 34296 12860 34302 12872
rect 39025 12869 39037 12872
rect 39071 12900 39083 12903
rect 39071 12872 39620 12900
rect 39071 12869 39083 12872
rect 39025 12863 39083 12869
rect 33965 12835 34023 12841
rect 33965 12801 33977 12835
rect 34011 12832 34023 12835
rect 34330 12832 34336 12844
rect 34011 12804 34336 12832
rect 34011 12801 34023 12804
rect 33965 12795 34023 12801
rect 34330 12792 34336 12804
rect 34388 12792 34394 12844
rect 35434 12792 35440 12844
rect 35492 12832 35498 12844
rect 35814 12835 35872 12841
rect 35814 12832 35826 12835
rect 35492 12804 35826 12832
rect 35492 12792 35498 12804
rect 35814 12801 35826 12804
rect 35860 12801 35872 12835
rect 35814 12795 35872 12801
rect 36081 12835 36139 12841
rect 36081 12801 36093 12835
rect 36127 12832 36139 12835
rect 37090 12832 37096 12844
rect 36127 12804 37096 12832
rect 36127 12801 36139 12804
rect 36081 12795 36139 12801
rect 37090 12792 37096 12804
rect 37148 12792 37154 12844
rect 39592 12841 39620 12872
rect 39577 12835 39635 12841
rect 39577 12801 39589 12835
rect 39623 12801 39635 12835
rect 39577 12795 39635 12801
rect 39853 12835 39911 12841
rect 39853 12801 39865 12835
rect 39899 12832 39911 12835
rect 40494 12832 40500 12844
rect 39899 12804 40500 12832
rect 39899 12801 39911 12804
rect 39853 12795 39911 12801
rect 40494 12792 40500 12804
rect 40552 12792 40558 12844
rect 34238 12764 34244 12776
rect 34199 12736 34244 12764
rect 34238 12724 34244 12736
rect 34296 12724 34302 12776
rect 33042 12656 33048 12708
rect 33100 12696 33106 12708
rect 34701 12699 34759 12705
rect 34701 12696 34713 12699
rect 33100 12668 34713 12696
rect 33100 12656 33106 12668
rect 34701 12665 34713 12668
rect 34747 12665 34759 12699
rect 37366 12696 37372 12708
rect 34701 12659 34759 12665
rect 37292 12668 37372 12696
rect 37292 12628 37320 12668
rect 37366 12656 37372 12668
rect 37424 12656 37430 12708
rect 38838 12696 38844 12708
rect 38799 12668 38844 12696
rect 38838 12656 38844 12668
rect 38896 12656 38902 12708
rect 37458 12628 37464 12640
rect 32968 12600 37320 12628
rect 37419 12600 37464 12628
rect 32125 12591 32183 12597
rect 37458 12588 37464 12600
rect 37516 12588 37522 12640
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 1872 12396 5396 12424
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 1872 12229 1900 12396
rect 2774 12356 2780 12368
rect 2608 12328 2780 12356
rect 2608 12229 2636 12328
rect 2774 12316 2780 12328
rect 2832 12316 2838 12368
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 3970 12288 3976 12300
rect 3844 12260 3976 12288
rect 3844 12248 3850 12260
rect 3970 12248 3976 12260
rect 4028 12248 4034 12300
rect 1673 12223 1731 12229
rect 1673 12220 1685 12223
rect 1452 12192 1685 12220
rect 1452 12180 1458 12192
rect 1673 12189 1685 12192
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 2756 12223 2814 12229
rect 2961 12223 3019 12229
rect 2756 12220 2768 12223
rect 2593 12183 2651 12189
rect 2700 12192 2768 12220
rect 2406 12112 2412 12164
rect 2464 12152 2470 12164
rect 2700 12152 2728 12192
rect 2756 12189 2768 12192
rect 2802 12189 2814 12223
rect 2756 12183 2814 12189
rect 2869 12217 2927 12223
rect 2869 12183 2881 12217
rect 2915 12183 2927 12217
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3234 12220 3240 12232
rect 3007 12192 3240 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 2869 12177 2927 12183
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 2464 12124 2728 12152
rect 2464 12112 2470 12124
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 2222 12084 2228 12096
rect 2087 12056 2228 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 2884 12084 2912 12177
rect 3050 12112 3056 12164
rect 3108 12152 3114 12164
rect 4218 12155 4276 12161
rect 4218 12152 4230 12155
rect 3108 12124 4230 12152
rect 3108 12112 3114 12124
rect 4218 12121 4230 12124
rect 4264 12121 4276 12155
rect 4218 12115 4276 12121
rect 2648 12056 2912 12084
rect 3237 12087 3295 12093
rect 2648 12044 2654 12056
rect 3237 12053 3249 12087
rect 3283 12084 3295 12087
rect 4706 12084 4712 12096
rect 3283 12056 4712 12084
rect 3283 12053 3295 12056
rect 3237 12047 3295 12053
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 5368 12093 5396 12396
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 10689 12427 10747 12433
rect 8260 12396 10640 12424
rect 8260 12384 8266 12396
rect 7926 12356 7932 12368
rect 7839 12328 7932 12356
rect 7926 12316 7932 12328
rect 7984 12356 7990 12368
rect 9582 12356 9588 12368
rect 7984 12328 9588 12356
rect 7984 12316 7990 12328
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12325 10563 12359
rect 10612 12356 10640 12396
rect 10689 12393 10701 12427
rect 10735 12424 10747 12427
rect 11514 12424 11520 12436
rect 10735 12396 11520 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 12986 12424 12992 12436
rect 12947 12396 12992 12424
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 15289 12427 15347 12433
rect 13596 12396 14228 12424
rect 13596 12384 13602 12396
rect 14090 12356 14096 12368
rect 10612 12328 14096 12356
rect 10505 12319 10563 12325
rect 6546 12220 6552 12232
rect 6507 12192 6552 12220
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 6805 12223 6863 12229
rect 6805 12220 6817 12223
rect 6696 12192 6817 12220
rect 6696 12180 6702 12192
rect 6805 12189 6817 12192
rect 6851 12189 6863 12223
rect 6805 12183 6863 12189
rect 7834 12112 7840 12164
rect 7892 12152 7898 12164
rect 7892 12124 8340 12152
rect 7892 12112 7898 12124
rect 5353 12087 5411 12093
rect 5353 12053 5365 12087
rect 5399 12084 5411 12087
rect 7466 12084 7472 12096
rect 5399 12056 7472 12084
rect 5399 12053 5411 12056
rect 5353 12047 5411 12053
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 8312 12084 8340 12124
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10229 12155 10287 12161
rect 10229 12152 10241 12155
rect 9916 12124 10241 12152
rect 9916 12112 9922 12124
rect 10229 12121 10241 12124
rect 10275 12121 10287 12155
rect 10520 12152 10548 12319
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 14200 12356 14228 12396
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15654 12424 15660 12436
rect 15335 12396 15660 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 23661 12427 23719 12433
rect 15764 12396 20392 12424
rect 15764 12356 15792 12396
rect 17862 12356 17868 12368
rect 14200 12328 15792 12356
rect 17420 12328 17868 12356
rect 13078 12288 13084 12300
rect 13039 12260 13084 12288
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 14182 12248 14188 12300
rect 14240 12288 14246 12300
rect 14240 12260 15148 12288
rect 14240 12248 14246 12260
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 10962 12220 10968 12232
rect 10836 12192 10968 12220
rect 10836 12180 10842 12192
rect 10962 12180 10968 12192
rect 11020 12220 11026 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 11020 12192 11161 12220
rect 11020 12180 11026 12192
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12220 11483 12223
rect 11882 12220 11888 12232
rect 11471 12192 11888 12220
rect 11471 12189 11483 12192
rect 11425 12183 11483 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 13170 12220 13176 12232
rect 13131 12192 13176 12220
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 15120 12229 15148 12260
rect 17420 12232 17448 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 20254 12356 20260 12368
rect 19300 12328 20260 12356
rect 19300 12316 19306 12328
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 18230 12288 18236 12300
rect 18064 12260 18236 12288
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12220 17187 12223
rect 17402 12220 17408 12232
rect 17175 12192 17408 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 11606 12152 11612 12164
rect 10520 12124 11612 12152
rect 10229 12115 10287 12121
rect 11606 12112 11612 12124
rect 11664 12152 11670 12164
rect 14936 12152 14964 12183
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 18064 12229 18092 12260
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17552 12192 17969 12220
rect 17552 12180 17558 12192
rect 17957 12189 17969 12192
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18325 12223 18383 12229
rect 18196 12192 18241 12220
rect 18196 12180 18202 12192
rect 18325 12189 18337 12223
rect 18371 12220 18383 12223
rect 19242 12220 19248 12232
rect 18371 12192 19248 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 16022 12152 16028 12164
rect 11664 12124 14964 12152
rect 15672 12124 16028 12152
rect 11664 12112 11670 12124
rect 12434 12084 12440 12096
rect 8312 12056 12440 12084
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 12894 12084 12900 12096
rect 12851 12056 12900 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 14461 12087 14519 12093
rect 14461 12053 14473 12087
rect 14507 12084 14519 12087
rect 15470 12084 15476 12096
rect 14507 12056 15476 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 15470 12044 15476 12056
rect 15528 12084 15534 12096
rect 15672 12084 15700 12124
rect 16022 12112 16028 12124
rect 16080 12112 16086 12164
rect 16884 12155 16942 12161
rect 16884 12121 16896 12155
rect 16930 12152 16942 12155
rect 17681 12155 17739 12161
rect 17681 12152 17693 12155
rect 16930 12124 17693 12152
rect 16930 12121 16942 12124
rect 16884 12115 16942 12121
rect 17681 12121 17693 12124
rect 17727 12121 17739 12155
rect 18340 12152 18368 12183
rect 19242 12180 19248 12192
rect 19300 12220 19306 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 19300 12192 19809 12220
rect 19300 12180 19306 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19960 12217 20018 12223
rect 19960 12214 19972 12217
rect 19797 12183 19855 12189
rect 19904 12186 19972 12214
rect 17681 12115 17739 12121
rect 18064 12124 18368 12152
rect 18064 12096 18092 12124
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 19904 12152 19932 12186
rect 19960 12183 19972 12186
rect 20006 12183 20018 12217
rect 19960 12177 20018 12183
rect 20073 12180 20079 12232
rect 20131 12229 20137 12232
rect 20131 12223 20150 12229
rect 20138 12189 20150 12223
rect 20185 12223 20243 12229
rect 20185 12220 20197 12223
rect 20131 12183 20150 12189
rect 20180 12189 20197 12220
rect 20231 12189 20243 12223
rect 20364 12220 20392 12396
rect 23661 12393 23673 12427
rect 23707 12424 23719 12427
rect 24670 12424 24676 12436
rect 23707 12396 24676 12424
rect 23707 12393 23719 12396
rect 23661 12387 23719 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 26602 12384 26608 12436
rect 26660 12424 26666 12436
rect 26973 12427 27031 12433
rect 26973 12424 26985 12427
rect 26660 12396 26985 12424
rect 26660 12384 26666 12396
rect 26973 12393 26985 12396
rect 27019 12424 27031 12427
rect 27522 12424 27528 12436
rect 27019 12396 27528 12424
rect 27019 12393 27031 12396
rect 26973 12387 27031 12393
rect 27522 12384 27528 12396
rect 27580 12384 27586 12436
rect 28442 12384 28448 12436
rect 28500 12424 28506 12436
rect 28902 12424 28908 12436
rect 28500 12396 28908 12424
rect 28500 12384 28506 12396
rect 28902 12384 28908 12396
rect 28960 12384 28966 12436
rect 29822 12424 29828 12436
rect 29783 12396 29828 12424
rect 29822 12384 29828 12396
rect 29880 12384 29886 12436
rect 30282 12424 30288 12436
rect 30243 12396 30288 12424
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 30929 12427 30987 12433
rect 30929 12393 30941 12427
rect 30975 12424 30987 12427
rect 33594 12424 33600 12436
rect 30975 12396 33600 12424
rect 30975 12393 30987 12396
rect 30929 12387 30987 12393
rect 33594 12384 33600 12396
rect 33652 12384 33658 12436
rect 33796 12396 34744 12424
rect 24026 12316 24032 12368
rect 24084 12356 24090 12368
rect 28997 12359 29055 12365
rect 24084 12328 27614 12356
rect 24084 12316 24090 12328
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 22646 12288 22652 12300
rect 22066 12260 22652 12288
rect 22066 12220 22094 12260
rect 22646 12248 22652 12260
rect 22704 12288 22710 12300
rect 22833 12291 22891 12297
rect 22833 12288 22845 12291
rect 22704 12260 22845 12288
rect 22704 12248 22710 12260
rect 22833 12257 22845 12260
rect 22879 12257 22891 12291
rect 22833 12251 22891 12257
rect 25038 12248 25044 12300
rect 25096 12288 25102 12300
rect 25133 12291 25191 12297
rect 25133 12288 25145 12291
rect 25096 12260 25145 12288
rect 25096 12248 25102 12260
rect 25133 12257 25145 12260
rect 25179 12288 25191 12291
rect 26970 12288 26976 12300
rect 25179 12260 26976 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 26970 12248 26976 12260
rect 27028 12248 27034 12300
rect 27586 12288 27614 12328
rect 28997 12325 29009 12359
rect 29043 12356 29055 12359
rect 29043 12328 29960 12356
rect 29043 12325 29055 12328
rect 28997 12319 29055 12325
rect 28902 12288 28908 12300
rect 27586 12260 28672 12288
rect 28644 12232 28672 12260
rect 28736 12260 28908 12288
rect 20364 12192 22094 12220
rect 20180 12183 20243 12189
rect 20131 12180 20137 12183
rect 19024 12124 19932 12152
rect 19024 12112 19030 12124
rect 15528 12056 15700 12084
rect 15749 12087 15807 12093
rect 15528 12044 15534 12056
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 17862 12084 17868 12096
rect 15795 12056 17868 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 18046 12044 18052 12096
rect 18104 12044 18110 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 19116 12056 19349 12084
rect 19116 12044 19122 12056
rect 19337 12053 19349 12056
rect 19383 12084 19395 12087
rect 19426 12084 19432 12096
rect 19383 12056 19432 12084
rect 19383 12053 19395 12056
rect 19337 12047 19395 12053
rect 19426 12044 19432 12056
rect 19484 12084 19490 12096
rect 20180 12084 20208 12183
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 23014 12220 23020 12232
rect 22244 12192 23020 12220
rect 22244 12180 22250 12192
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 23845 12223 23903 12229
rect 23845 12220 23857 12223
rect 23768 12192 23857 12220
rect 20441 12155 20499 12161
rect 20441 12121 20453 12155
rect 20487 12152 20499 12155
rect 21146 12155 21204 12161
rect 21146 12152 21158 12155
rect 20487 12124 21158 12152
rect 20487 12121 20499 12124
rect 20441 12115 20499 12121
rect 21146 12121 21158 12124
rect 21192 12121 21204 12155
rect 21146 12115 21204 12121
rect 23768 12096 23796 12192
rect 23845 12189 23857 12192
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 24578 12180 24584 12232
rect 24636 12220 24642 12232
rect 24762 12220 24768 12232
rect 24636 12192 24768 12220
rect 24636 12180 24642 12192
rect 24762 12180 24768 12192
rect 24820 12220 24826 12232
rect 24857 12223 24915 12229
rect 24857 12220 24869 12223
rect 24820 12192 24869 12220
rect 24820 12180 24826 12192
rect 24857 12189 24869 12192
rect 24903 12189 24915 12223
rect 26142 12220 26148 12232
rect 26103 12192 26148 12220
rect 24857 12183 24915 12189
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 28445 12223 28503 12229
rect 28445 12220 28457 12223
rect 26252 12192 28457 12220
rect 24026 12112 24032 12164
rect 24084 12152 24090 12164
rect 26252 12152 26280 12192
rect 28445 12189 28457 12192
rect 28491 12189 28503 12223
rect 28626 12220 28632 12232
rect 28539 12192 28632 12220
rect 28445 12183 28503 12189
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 28736 12229 28764 12260
rect 28902 12248 28908 12260
rect 28960 12248 28966 12300
rect 29932 12297 29960 12328
rect 32398 12316 32404 12368
rect 32456 12356 32462 12368
rect 32950 12356 32956 12368
rect 32456 12328 32956 12356
rect 32456 12316 32462 12328
rect 32950 12316 32956 12328
rect 33008 12316 33014 12368
rect 33134 12316 33140 12368
rect 33192 12356 33198 12368
rect 33796 12356 33824 12396
rect 34514 12356 34520 12368
rect 33192 12328 33824 12356
rect 33980 12328 34520 12356
rect 33192 12316 33198 12328
rect 29917 12291 29975 12297
rect 29917 12257 29929 12291
rect 29963 12257 29975 12291
rect 29917 12251 29975 12257
rect 32309 12291 32367 12297
rect 32309 12257 32321 12291
rect 32355 12288 32367 12291
rect 32674 12288 32680 12300
rect 32355 12260 32680 12288
rect 32355 12257 32367 12260
rect 32309 12251 32367 12257
rect 32674 12248 32680 12260
rect 32732 12248 32738 12300
rect 33980 12288 34008 12328
rect 34514 12316 34520 12328
rect 34572 12316 34578 12368
rect 33888 12260 34008 12288
rect 28721 12223 28779 12229
rect 28721 12189 28733 12223
rect 28767 12189 28779 12223
rect 28721 12183 28779 12189
rect 28810 12180 28816 12232
rect 28868 12220 28874 12232
rect 28868 12192 28913 12220
rect 28868 12180 28874 12192
rect 29638 12180 29644 12232
rect 29696 12220 29702 12232
rect 29825 12223 29883 12229
rect 29825 12220 29837 12223
rect 29696 12192 29837 12220
rect 29696 12180 29702 12192
rect 29825 12189 29837 12192
rect 29871 12189 29883 12223
rect 29825 12183 29883 12189
rect 30101 12223 30159 12229
rect 30101 12189 30113 12223
rect 30147 12220 30159 12223
rect 31110 12220 31116 12232
rect 30147 12192 31116 12220
rect 30147 12189 30159 12192
rect 30101 12183 30159 12189
rect 31110 12180 31116 12192
rect 31168 12180 31174 12232
rect 33410 12180 33416 12232
rect 33468 12220 33474 12232
rect 33888 12229 33916 12260
rect 33735 12223 33793 12229
rect 33735 12220 33747 12223
rect 33468 12192 33747 12220
rect 33468 12180 33474 12192
rect 33735 12189 33747 12192
rect 33781 12189 33793 12223
rect 33735 12183 33793 12189
rect 33870 12223 33928 12229
rect 33870 12189 33882 12223
rect 33916 12189 33928 12223
rect 33870 12183 33928 12189
rect 33965 12223 34023 12229
rect 33965 12189 33977 12223
rect 34011 12220 34023 12223
rect 34149 12223 34207 12229
rect 34011 12192 34100 12220
rect 34011 12189 34023 12192
rect 33965 12183 34023 12189
rect 24084 12124 26280 12152
rect 26329 12155 26387 12161
rect 24084 12112 24090 12124
rect 26329 12121 26341 12155
rect 26375 12152 26387 12155
rect 28534 12152 28540 12164
rect 26375 12124 28540 12152
rect 26375 12121 26387 12124
rect 26329 12115 26387 12121
rect 28534 12112 28540 12124
rect 28592 12112 28598 12164
rect 32064 12155 32122 12161
rect 32064 12121 32076 12155
rect 32110 12152 32122 12155
rect 33505 12155 33563 12161
rect 33505 12152 33517 12155
rect 32110 12124 33517 12152
rect 32110 12121 32122 12124
rect 32064 12115 32122 12121
rect 33505 12121 33517 12124
rect 33551 12121 33563 12155
rect 34072 12152 34100 12192
rect 34149 12189 34161 12223
rect 34195 12220 34207 12223
rect 34238 12220 34244 12232
rect 34195 12192 34244 12220
rect 34195 12189 34207 12192
rect 34149 12183 34207 12189
rect 34238 12180 34244 12192
rect 34296 12180 34302 12232
rect 34716 12229 34744 12396
rect 35342 12384 35348 12436
rect 35400 12424 35406 12436
rect 37458 12424 37464 12436
rect 35400 12396 37464 12424
rect 35400 12384 35406 12396
rect 37458 12384 37464 12396
rect 37516 12384 37522 12436
rect 39025 12427 39083 12433
rect 39025 12393 39037 12427
rect 39071 12424 39083 12427
rect 39114 12424 39120 12436
rect 39071 12396 39120 12424
rect 39071 12393 39083 12396
rect 39025 12387 39083 12393
rect 39114 12384 39120 12396
rect 39172 12384 39178 12436
rect 35710 12356 35716 12368
rect 35671 12328 35716 12356
rect 35710 12316 35716 12328
rect 35768 12316 35774 12368
rect 34701 12223 34759 12229
rect 34701 12189 34713 12223
rect 34747 12189 34759 12223
rect 34701 12183 34759 12189
rect 34885 12223 34943 12229
rect 34885 12189 34897 12223
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 34330 12152 34336 12164
rect 34072 12124 34336 12152
rect 33505 12115 33563 12121
rect 34330 12112 34336 12124
rect 34388 12112 34394 12164
rect 34900 12152 34928 12183
rect 35894 12180 35900 12232
rect 35952 12220 35958 12232
rect 36826 12223 36884 12229
rect 36826 12220 36838 12223
rect 35952 12192 36838 12220
rect 35952 12180 35958 12192
rect 36826 12189 36838 12192
rect 36872 12189 36884 12223
rect 37090 12220 37096 12232
rect 37051 12192 37096 12220
rect 36826 12183 36884 12189
rect 37090 12180 37096 12192
rect 37148 12180 37154 12232
rect 37458 12180 37464 12232
rect 37516 12220 37522 12232
rect 37553 12223 37611 12229
rect 37553 12220 37565 12223
rect 37516 12192 37565 12220
rect 37516 12180 37522 12192
rect 37553 12189 37565 12192
rect 37599 12189 37611 12223
rect 37553 12183 37611 12189
rect 39022 12180 39028 12232
rect 39080 12220 39086 12232
rect 40037 12223 40095 12229
rect 40037 12220 40049 12223
rect 39080 12192 40049 12220
rect 39080 12180 39086 12192
rect 40037 12189 40049 12192
rect 40083 12189 40095 12223
rect 40037 12183 40095 12189
rect 40221 12217 40279 12223
rect 40221 12183 40233 12217
rect 40267 12183 40279 12217
rect 40221 12177 40279 12183
rect 40316 12217 40374 12223
rect 40316 12183 40328 12217
rect 40362 12183 40374 12217
rect 40316 12177 40374 12183
rect 40402 12180 40408 12232
rect 40460 12220 40466 12232
rect 41141 12223 41199 12229
rect 41141 12220 41153 12223
rect 40460 12192 41153 12220
rect 40460 12180 40466 12192
rect 41141 12189 41153 12192
rect 41187 12189 41199 12223
rect 41141 12183 41199 12189
rect 34532 12124 34928 12152
rect 22278 12084 22284 12096
rect 19484 12056 20208 12084
rect 22239 12056 22284 12084
rect 19484 12044 19490 12056
rect 22278 12044 22284 12056
rect 22336 12084 22342 12096
rect 23106 12084 23112 12096
rect 22336 12056 23112 12084
rect 22336 12044 22342 12056
rect 23106 12044 23112 12056
rect 23164 12044 23170 12096
rect 23201 12087 23259 12093
rect 23201 12053 23213 12087
rect 23247 12084 23259 12087
rect 23750 12084 23756 12096
rect 23247 12056 23756 12084
rect 23247 12053 23259 12056
rect 23201 12047 23259 12053
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 26510 12084 26516 12096
rect 26471 12056 26516 12084
rect 26510 12044 26516 12056
rect 26568 12044 26574 12096
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 31018 12084 31024 12096
rect 26660 12056 31024 12084
rect 26660 12044 26666 12056
rect 31018 12044 31024 12056
rect 31076 12044 31082 12096
rect 32950 12044 32956 12096
rect 33008 12084 33014 12096
rect 34532 12084 34560 12124
rect 40236 12096 40264 12177
rect 40328 12096 40356 12177
rect 40678 12152 40684 12164
rect 40639 12124 40684 12152
rect 40678 12112 40684 12124
rect 40736 12112 40742 12164
rect 33008 12056 34560 12084
rect 33008 12044 33014 12056
rect 34606 12044 34612 12096
rect 34664 12084 34670 12096
rect 34793 12087 34851 12093
rect 34793 12084 34805 12087
rect 34664 12056 34805 12084
rect 34664 12044 34670 12056
rect 34793 12053 34805 12056
rect 34839 12053 34851 12087
rect 34793 12047 34851 12053
rect 40218 12044 40224 12096
rect 40276 12044 40282 12096
rect 40310 12044 40316 12096
rect 40368 12044 40374 12096
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 2464 11852 3157 11880
rect 2464 11840 2470 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3145 11843 3203 11849
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 3292 11852 4077 11880
rect 3292 11840 3298 11852
rect 4065 11849 4077 11852
rect 4111 11880 4123 11883
rect 5350 11880 5356 11892
rect 4111 11852 5356 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 7248 11852 7389 11880
rect 7248 11840 7254 11852
rect 7377 11849 7389 11852
rect 7423 11849 7435 11883
rect 7377 11843 7435 11849
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 13081 11883 13139 11889
rect 7524 11852 12112 11880
rect 7524 11840 7530 11852
rect 2590 11812 2596 11824
rect 2332 11784 2596 11812
rect 1762 11704 1768 11756
rect 1820 11744 1826 11756
rect 2038 11744 2044 11756
rect 1820 11716 2044 11744
rect 1820 11704 1826 11716
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2332 11753 2360 11784
rect 2590 11772 2596 11784
rect 2648 11772 2654 11824
rect 3513 11815 3571 11821
rect 3513 11812 3525 11815
rect 3160 11784 3525 11812
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 2455 11747 2513 11753
rect 2455 11713 2467 11747
rect 2501 11744 2513 11747
rect 2501 11716 2636 11744
rect 2501 11713 2513 11716
rect 2455 11707 2513 11713
rect 2608 11676 2636 11716
rect 2682 11704 2688 11756
rect 2740 11744 2746 11756
rect 3160 11744 3188 11784
rect 3513 11781 3525 11784
rect 3559 11781 3571 11815
rect 3513 11775 3571 11781
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 9364 11784 9409 11812
rect 9364 11772 9370 11784
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 10229 11815 10287 11821
rect 10229 11812 10241 11815
rect 9640 11784 10088 11812
rect 9640 11772 9646 11784
rect 2740 11716 3188 11744
rect 3329 11747 3387 11753
rect 2740 11704 2746 11716
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 5810 11744 5816 11756
rect 3375 11716 5816 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 9030 11744 9036 11756
rect 8991 11716 9036 11744
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 9180 11716 9229 11744
rect 9180 11704 9186 11716
rect 9217 11713 9229 11716
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 9447 11747 9505 11753
rect 9447 11713 9459 11747
rect 9493 11744 9505 11747
rect 9674 11744 9680 11756
rect 9493 11716 9680 11744
rect 9493 11713 9505 11716
rect 9447 11707 9505 11713
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 10060 11753 10088 11784
rect 10152 11784 10241 11812
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 2866 11676 2872 11688
rect 2608 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 3142 11636 3148 11688
rect 3200 11676 3206 11688
rect 9306 11676 9312 11688
rect 3200 11648 9312 11676
rect 3200 11636 3206 11648
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 10152 11676 10180 11784
rect 10229 11781 10241 11784
rect 10275 11812 10287 11815
rect 11514 11812 11520 11824
rect 10275 11784 11520 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 11514 11772 11520 11784
rect 11572 11772 11578 11824
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 12084 11821 12112 11852
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 13630 11880 13636 11892
rect 13127 11852 13636 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 14608 11852 14657 11880
rect 14608 11840 14614 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 18138 11880 18144 11892
rect 18095 11852 18144 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18966 11840 18972 11892
rect 19024 11880 19030 11892
rect 19337 11883 19395 11889
rect 19337 11880 19349 11883
rect 19024 11852 19349 11880
rect 19024 11840 19030 11852
rect 19337 11849 19349 11852
rect 19383 11849 19395 11883
rect 19337 11843 19395 11849
rect 23382 11840 23388 11892
rect 23440 11880 23446 11892
rect 24578 11880 24584 11892
rect 23440 11852 24440 11880
rect 24539 11852 24584 11880
rect 23440 11840 23446 11852
rect 11977 11815 12035 11821
rect 11977 11812 11989 11815
rect 11756 11784 11989 11812
rect 11756 11772 11762 11784
rect 11977 11781 11989 11784
rect 12023 11781 12035 11815
rect 11977 11775 12035 11781
rect 12069 11815 12127 11821
rect 12069 11781 12081 11815
rect 12115 11781 12127 11815
rect 12069 11775 12127 11781
rect 13909 11815 13967 11821
rect 13909 11781 13921 11815
rect 13955 11812 13967 11815
rect 15746 11812 15752 11824
rect 13955 11784 15752 11812
rect 13955 11781 13967 11784
rect 13909 11775 13967 11781
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 17586 11772 17592 11824
rect 17644 11812 17650 11824
rect 17681 11815 17739 11821
rect 17681 11812 17693 11815
rect 17644 11784 17693 11812
rect 17644 11772 17650 11784
rect 17681 11781 17693 11784
rect 17727 11812 17739 11815
rect 19153 11815 19211 11821
rect 17727 11784 19012 11812
rect 17727 11781 17739 11784
rect 17681 11775 17739 11781
rect 18984 11756 19012 11784
rect 19153 11781 19165 11815
rect 19199 11812 19211 11815
rect 19702 11812 19708 11824
rect 19199 11784 19708 11812
rect 19199 11781 19211 11784
rect 19153 11775 19211 11781
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 22005 11815 22063 11821
rect 22005 11781 22017 11815
rect 22051 11812 22063 11815
rect 23566 11812 23572 11824
rect 22051 11784 23572 11812
rect 22051 11781 22063 11784
rect 22005 11775 22063 11781
rect 23566 11772 23572 11784
rect 23624 11812 23630 11824
rect 24412 11812 24440 11852
rect 24578 11840 24584 11852
rect 24636 11840 24642 11892
rect 25498 11880 25504 11892
rect 25459 11852 25504 11880
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 27246 11880 27252 11892
rect 26206 11852 27252 11880
rect 24946 11812 24952 11824
rect 23624 11784 23796 11812
rect 24412 11784 24952 11812
rect 23624 11772 23630 11784
rect 10318 11744 10324 11756
rect 10279 11716 10324 11744
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10962 11744 10968 11756
rect 10459 11716 10968 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 9416 11648 10180 11676
rect 2685 11611 2743 11617
rect 2685 11577 2697 11611
rect 2731 11608 2743 11611
rect 3050 11608 3056 11620
rect 2731 11580 3056 11608
rect 2731 11577 2743 11580
rect 2685 11571 2743 11577
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 9214 11608 9220 11620
rect 6932 11580 9220 11608
rect 6932 11552 6960 11580
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 6914 11540 6920 11552
rect 6875 11512 6920 11540
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 7984 11512 8401 11540
rect 7984 11500 7990 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 9416 11540 9444 11648
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10428 11608 10456 11707
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11793 11747 11851 11753
rect 11793 11744 11805 11747
rect 11388 11716 11805 11744
rect 11388 11704 11394 11716
rect 11793 11713 11805 11716
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11744 12955 11747
rect 13354 11744 13360 11756
rect 12943 11716 13360 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12176 11676 12204 11707
rect 13354 11704 13360 11716
rect 13412 11744 13418 11756
rect 13725 11747 13783 11753
rect 13725 11744 13737 11747
rect 13412 11716 13737 11744
rect 13412 11704 13418 11716
rect 13725 11713 13737 11716
rect 13771 11713 13783 11747
rect 13725 11707 13783 11713
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14550 11744 14556 11756
rect 14240 11716 14556 11744
rect 14240 11704 14246 11716
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 17862 11744 17868 11756
rect 17775 11716 17868 11744
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 18966 11744 18972 11756
rect 18927 11716 18972 11744
rect 18966 11704 18972 11716
rect 19024 11704 19030 11756
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19300 11716 19809 11744
rect 19300 11704 19306 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19978 11744 19984 11756
rect 19939 11716 19984 11744
rect 19797 11707 19855 11713
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20070 11704 20076 11756
rect 20128 11744 20134 11756
rect 20254 11753 20260 11756
rect 20211 11747 20260 11753
rect 20128 11716 20173 11744
rect 20128 11704 20134 11716
rect 20211 11713 20223 11747
rect 20257 11713 20260 11747
rect 20211 11707 20260 11713
rect 20254 11704 20260 11707
rect 20312 11744 20318 11756
rect 20622 11744 20628 11756
rect 20312 11716 20628 11744
rect 20312 11704 20318 11716
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 21082 11744 21088 11756
rect 21043 11716 21088 11744
rect 21082 11704 21088 11716
rect 21140 11704 21146 11756
rect 23768 11753 23796 11784
rect 24946 11772 24952 11784
rect 25004 11812 25010 11824
rect 26206 11812 26234 11852
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 27430 11840 27436 11892
rect 27488 11880 27494 11892
rect 30009 11883 30067 11889
rect 30009 11880 30021 11883
rect 27488 11852 30021 11880
rect 27488 11840 27494 11852
rect 30009 11849 30021 11852
rect 30055 11849 30067 11883
rect 30650 11880 30656 11892
rect 30611 11852 30656 11880
rect 30009 11843 30067 11849
rect 30650 11840 30656 11852
rect 30708 11840 30714 11892
rect 33134 11880 33140 11892
rect 31404 11852 33140 11880
rect 25004 11784 26234 11812
rect 25004 11772 25010 11784
rect 26510 11772 26516 11824
rect 26568 11812 26574 11824
rect 26568 11784 27179 11812
rect 26568 11772 26574 11784
rect 27151 11756 27179 11784
rect 23293 11747 23351 11753
rect 23293 11744 23305 11747
rect 22066 11716 23305 11744
rect 11940 11648 12204 11676
rect 11940 11636 11946 11648
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 12492 11648 17141 11676
rect 12492 11636 12498 11648
rect 17129 11645 17141 11648
rect 17175 11676 17187 11679
rect 17494 11676 17500 11688
rect 17175 11648 17500 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 17880 11676 17908 11704
rect 19518 11676 19524 11688
rect 17880 11648 19524 11676
rect 19518 11636 19524 11648
rect 19576 11636 19582 11688
rect 21910 11636 21916 11688
rect 21968 11676 21974 11688
rect 22066 11676 22094 11716
rect 23293 11713 23305 11716
rect 23339 11713 23351 11747
rect 23293 11707 23351 11713
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11713 23811 11747
rect 23753 11707 23811 11713
rect 23934 11704 23940 11756
rect 23992 11744 23998 11756
rect 23992 11716 24085 11744
rect 23992 11704 23998 11716
rect 24670 11704 24676 11756
rect 24728 11744 24734 11756
rect 24765 11747 24823 11753
rect 24765 11744 24777 11747
rect 24728 11716 24777 11744
rect 24728 11704 24734 11716
rect 24765 11713 24777 11716
rect 24811 11713 24823 11747
rect 25038 11744 25044 11756
rect 24999 11716 25044 11744
rect 24765 11707 24823 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25682 11744 25688 11756
rect 25643 11716 25688 11744
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 25958 11744 25964 11756
rect 25919 11716 25964 11744
rect 25958 11704 25964 11716
rect 26016 11704 26022 11756
rect 26970 11744 26976 11756
rect 26931 11716 26976 11744
rect 26970 11704 26976 11716
rect 27028 11704 27034 11756
rect 27136 11750 27194 11756
rect 27264 11753 27292 11840
rect 28534 11772 28540 11824
rect 28592 11812 28598 11824
rect 28721 11815 28779 11821
rect 28721 11812 28733 11815
rect 28592 11784 28733 11812
rect 28592 11772 28598 11784
rect 28721 11781 28733 11784
rect 28767 11781 28779 11815
rect 30834 11812 30840 11824
rect 28721 11775 28779 11781
rect 28920 11784 30840 11812
rect 27136 11716 27148 11750
rect 27182 11716 27194 11750
rect 27136 11710 27194 11716
rect 27249 11747 27307 11753
rect 27249 11713 27261 11747
rect 27295 11713 27307 11747
rect 27249 11707 27307 11713
rect 27387 11747 27445 11753
rect 27387 11713 27399 11747
rect 27433 11744 27445 11747
rect 27522 11744 27528 11756
rect 27433 11716 27528 11744
rect 27433 11713 27445 11716
rect 27387 11707 27445 11713
rect 27522 11704 27528 11716
rect 27580 11704 27586 11756
rect 28442 11744 28448 11756
rect 28403 11716 28448 11744
rect 28442 11704 28448 11716
rect 28500 11704 28506 11756
rect 28626 11744 28632 11756
rect 28587 11716 28632 11744
rect 28626 11704 28632 11716
rect 28684 11704 28690 11756
rect 28810 11744 28816 11756
rect 28771 11716 28816 11744
rect 28810 11704 28816 11716
rect 28868 11704 28874 11756
rect 23014 11676 23020 11688
rect 21968 11648 22094 11676
rect 22975 11648 23020 11676
rect 21968 11636 21974 11648
rect 23014 11636 23020 11648
rect 23072 11676 23078 11688
rect 23952 11676 23980 11704
rect 24854 11676 24860 11688
rect 23072 11648 23980 11676
rect 24815 11648 24860 11676
rect 23072 11636 23078 11648
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25774 11676 25780 11688
rect 25735 11648 25780 11676
rect 25774 11636 25780 11648
rect 25832 11636 25838 11688
rect 26602 11676 26608 11688
rect 25884 11648 26608 11676
rect 19794 11608 19800 11620
rect 9732 11580 10456 11608
rect 17880 11580 19800 11608
rect 9732 11568 9738 11580
rect 9582 11540 9588 11552
rect 9180 11512 9444 11540
rect 9543 11512 9588 11540
rect 9180 11500 9186 11512
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 10594 11540 10600 11552
rect 10555 11512 10600 11540
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 12345 11543 12403 11549
rect 12345 11509 12357 11543
rect 12391 11540 12403 11543
rect 17880 11540 17908 11580
rect 19794 11568 19800 11580
rect 19852 11568 19858 11620
rect 12391 11512 17908 11540
rect 12391 11509 12403 11512
rect 12345 11503 12403 11509
rect 18322 11500 18328 11552
rect 18380 11540 18386 11552
rect 20070 11540 20076 11552
rect 18380 11512 20076 11540
rect 18380 11500 18386 11512
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20438 11540 20444 11552
rect 20399 11512 20444 11540
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 20901 11543 20959 11549
rect 20901 11540 20913 11543
rect 20588 11512 20913 11540
rect 20588 11500 20594 11512
rect 20901 11509 20913 11512
rect 20947 11509 20959 11543
rect 23842 11540 23848 11552
rect 23803 11512 23848 11540
rect 20901 11503 20959 11509
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 25041 11543 25099 11549
rect 25041 11509 25053 11543
rect 25087 11540 25099 11543
rect 25884 11540 25912 11648
rect 26602 11636 26608 11648
rect 26660 11636 26666 11688
rect 28920 11676 28948 11784
rect 30834 11772 30840 11784
rect 30892 11772 30898 11824
rect 28994 11704 29000 11756
rect 29052 11744 29058 11756
rect 29549 11747 29607 11753
rect 29549 11744 29561 11747
rect 29052 11716 29561 11744
rect 29052 11704 29058 11716
rect 29549 11713 29561 11716
rect 29595 11713 29607 11747
rect 29549 11707 29607 11713
rect 29825 11747 29883 11753
rect 29825 11713 29837 11747
rect 29871 11744 29883 11747
rect 31294 11744 31300 11756
rect 29871 11716 31300 11744
rect 29871 11713 29883 11716
rect 29825 11707 29883 11713
rect 31294 11704 31300 11716
rect 31352 11704 31358 11756
rect 31404 11753 31432 11852
rect 33134 11840 33140 11852
rect 33192 11840 33198 11892
rect 33781 11883 33839 11889
rect 33781 11849 33793 11883
rect 33827 11880 33839 11883
rect 34330 11880 34336 11892
rect 33827 11852 34336 11880
rect 33827 11849 33839 11852
rect 33781 11843 33839 11849
rect 34330 11840 34336 11852
rect 34388 11840 34394 11892
rect 35345 11883 35403 11889
rect 35345 11849 35357 11883
rect 35391 11880 35403 11883
rect 35434 11880 35440 11892
rect 35391 11852 35440 11880
rect 35391 11849 35403 11852
rect 35345 11843 35403 11849
rect 35434 11840 35440 11852
rect 35492 11840 35498 11892
rect 39022 11880 39028 11892
rect 35829 11852 39028 11880
rect 32769 11815 32827 11821
rect 32769 11781 32781 11815
rect 32815 11812 32827 11815
rect 33042 11812 33048 11824
rect 32815 11784 33048 11812
rect 32815 11781 32827 11784
rect 32769 11775 32827 11781
rect 33042 11772 33048 11784
rect 33100 11772 33106 11824
rect 33594 11812 33600 11824
rect 33555 11784 33600 11812
rect 33594 11772 33600 11784
rect 33652 11772 33658 11824
rect 34514 11772 34520 11824
rect 34572 11812 34578 11824
rect 35710 11812 35716 11824
rect 34572 11784 35716 11812
rect 34572 11772 34578 11784
rect 31389 11747 31447 11753
rect 31389 11713 31401 11747
rect 31435 11713 31447 11747
rect 31389 11707 31447 11713
rect 32953 11747 33011 11753
rect 32953 11713 32965 11747
rect 32999 11744 33011 11747
rect 33410 11744 33416 11756
rect 32999 11716 33416 11744
rect 32999 11713 33011 11716
rect 32953 11707 33011 11713
rect 33410 11704 33416 11716
rect 33468 11704 33474 11756
rect 34238 11704 34244 11756
rect 34296 11744 34302 11756
rect 34992 11753 35020 11784
rect 35710 11772 35716 11784
rect 35768 11772 35774 11824
rect 34701 11747 34759 11753
rect 34701 11744 34713 11747
rect 34296 11716 34713 11744
rect 34296 11704 34302 11716
rect 34701 11713 34713 11716
rect 34747 11713 34759 11747
rect 34864 11747 34922 11753
rect 34864 11744 34876 11747
rect 34701 11707 34759 11713
rect 34808 11716 34876 11744
rect 27448 11648 28948 11676
rect 29641 11679 29699 11685
rect 25087 11512 25912 11540
rect 25961 11543 26019 11549
rect 25087 11509 25099 11512
rect 25041 11503 25099 11509
rect 25961 11509 25973 11543
rect 26007 11540 26019 11543
rect 27448 11540 27476 11648
rect 29641 11645 29653 11679
rect 29687 11645 29699 11679
rect 29641 11639 29699 11645
rect 28997 11611 29055 11617
rect 28997 11577 29009 11611
rect 29043 11608 29055 11611
rect 29656 11608 29684 11639
rect 30650 11636 30656 11688
rect 30708 11676 30714 11688
rect 31205 11679 31263 11685
rect 31205 11676 31217 11679
rect 30708 11648 31217 11676
rect 30708 11636 30714 11648
rect 31205 11645 31217 11648
rect 31251 11645 31263 11679
rect 31205 11639 31263 11645
rect 32585 11679 32643 11685
rect 32585 11645 32597 11679
rect 32631 11676 32643 11679
rect 34808 11676 34836 11716
rect 34864 11713 34876 11716
rect 34910 11713 34922 11747
rect 34864 11707 34922 11713
rect 34980 11747 35038 11753
rect 34980 11713 34992 11747
rect 35026 11713 35038 11747
rect 34980 11707 35038 11713
rect 35066 11704 35072 11756
rect 35124 11744 35130 11756
rect 35829 11753 35857 11852
rect 39022 11840 39028 11852
rect 39080 11840 39086 11892
rect 40218 11880 40224 11892
rect 40179 11852 40224 11880
rect 40218 11840 40224 11852
rect 40276 11840 40282 11892
rect 37090 11772 37096 11824
rect 37148 11812 37154 11824
rect 37148 11784 38792 11812
rect 37148 11772 37154 11784
rect 35805 11747 35863 11753
rect 35124 11716 35169 11744
rect 35124 11704 35130 11716
rect 35805 11713 35817 11747
rect 35851 11713 35863 11747
rect 35805 11707 35863 11713
rect 35968 11747 36026 11753
rect 35968 11713 35980 11747
rect 36014 11713 36026 11747
rect 36084 11747 36142 11753
rect 36084 11744 36096 11747
rect 35968 11707 36026 11713
rect 36083 11713 36096 11744
rect 36130 11713 36142 11747
rect 36083 11707 36142 11713
rect 36219 11747 36277 11753
rect 36219 11713 36231 11747
rect 36265 11744 36277 11747
rect 36265 11742 36305 11744
rect 36354 11742 36360 11756
rect 36265 11714 36360 11742
rect 36265 11713 36277 11714
rect 36219 11707 36277 11713
rect 32631 11648 34836 11676
rect 32631 11645 32643 11648
rect 32585 11639 32643 11645
rect 35434 11636 35440 11688
rect 35492 11676 35498 11688
rect 35983 11676 36011 11707
rect 35492 11648 36011 11676
rect 36083 11676 36111 11707
rect 36354 11704 36360 11714
rect 36412 11744 36418 11756
rect 37274 11744 37280 11756
rect 36412 11716 37280 11744
rect 36412 11704 36418 11716
rect 37274 11704 37280 11716
rect 37332 11704 37338 11756
rect 38764 11753 38792 11784
rect 39758 11772 39764 11824
rect 39816 11812 39822 11824
rect 39853 11815 39911 11821
rect 39853 11812 39865 11815
rect 39816 11784 39865 11812
rect 39816 11772 39822 11784
rect 39853 11781 39865 11784
rect 39899 11781 39911 11815
rect 40678 11812 40684 11824
rect 39853 11775 39911 11781
rect 39960 11784 40684 11812
rect 38493 11747 38551 11753
rect 38493 11713 38505 11747
rect 38539 11744 38551 11747
rect 38749 11747 38807 11753
rect 38539 11716 38700 11744
rect 38539 11713 38551 11716
rect 38493 11707 38551 11713
rect 36446 11676 36452 11688
rect 36083 11648 36452 11676
rect 35492 11636 35498 11648
rect 36446 11636 36452 11648
rect 36504 11636 36510 11688
rect 38672 11676 38700 11716
rect 38749 11713 38761 11747
rect 38795 11744 38807 11747
rect 39114 11744 39120 11756
rect 38795 11716 39120 11744
rect 38795 11713 38807 11716
rect 38749 11707 38807 11713
rect 39114 11704 39120 11716
rect 39172 11704 39178 11756
rect 39960 11676 39988 11784
rect 40678 11772 40684 11784
rect 40736 11772 40742 11824
rect 40037 11747 40095 11753
rect 40037 11713 40049 11747
rect 40083 11713 40095 11747
rect 40037 11707 40095 11713
rect 38672 11648 39988 11676
rect 31386 11608 31392 11620
rect 29043 11580 29684 11608
rect 29840 11580 31392 11608
rect 29043 11577 29055 11580
rect 28997 11571 29055 11577
rect 27614 11540 27620 11552
rect 26007 11512 27476 11540
rect 27575 11512 27620 11540
rect 26007 11509 26019 11512
rect 25961 11503 26019 11509
rect 27614 11500 27620 11512
rect 27672 11500 27678 11552
rect 29840 11549 29868 11580
rect 31386 11568 31392 11580
rect 31444 11568 31450 11620
rect 34422 11568 34428 11620
rect 34480 11608 34486 11620
rect 37369 11611 37427 11617
rect 37369 11608 37381 11611
rect 34480 11580 37381 11608
rect 34480 11568 34486 11580
rect 37369 11577 37381 11580
rect 37415 11577 37427 11611
rect 37369 11571 37427 11577
rect 29825 11543 29883 11549
rect 29825 11509 29837 11543
rect 29871 11509 29883 11543
rect 29825 11503 29883 11509
rect 31573 11543 31631 11549
rect 31573 11509 31585 11543
rect 31619 11540 31631 11543
rect 34146 11540 34152 11552
rect 31619 11512 34152 11540
rect 31619 11509 31631 11512
rect 31573 11503 31631 11509
rect 34146 11500 34152 11512
rect 34204 11500 34210 11552
rect 36449 11543 36507 11549
rect 36449 11509 36461 11543
rect 36495 11540 36507 11543
rect 36814 11540 36820 11552
rect 36495 11512 36820 11540
rect 36495 11509 36507 11512
rect 36449 11503 36507 11509
rect 36814 11500 36820 11512
rect 36872 11500 36878 11552
rect 37384 11540 37412 11571
rect 40052 11540 40080 11707
rect 67634 11608 67640 11620
rect 67595 11580 67640 11608
rect 67634 11568 67640 11580
rect 67692 11568 67698 11620
rect 37384 11512 40080 11540
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 6546 11336 6552 11348
rect 4028 11308 6552 11336
rect 4028 11296 4034 11308
rect 6546 11296 6552 11308
rect 6604 11336 6610 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6604 11308 6745 11336
rect 6604 11296 6610 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 7282 11336 7288 11348
rect 7064 11308 7288 11336
rect 7064 11296 7070 11308
rect 7282 11296 7288 11308
rect 7340 11336 7346 11348
rect 9674 11336 9680 11348
rect 7340 11308 9680 11336
rect 7340 11296 7346 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 11020 11308 11529 11336
rect 11020 11296 11026 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 11517 11299 11575 11305
rect 12713 11339 12771 11345
rect 12713 11305 12725 11339
rect 12759 11336 12771 11339
rect 13170 11336 13176 11348
rect 12759 11308 13176 11336
rect 12759 11305 12771 11308
rect 12713 11299 12771 11305
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13538 11336 13544 11348
rect 13311 11308 13544 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 16390 11336 16396 11348
rect 16351 11308 16396 11336
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20073 11339 20131 11345
rect 20073 11336 20085 11339
rect 20036 11308 20085 11336
rect 20036 11296 20042 11308
rect 20073 11305 20085 11308
rect 20119 11305 20131 11339
rect 20073 11299 20131 11305
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 20714 11336 20720 11348
rect 20404 11308 20720 11336
rect 20404 11296 20410 11308
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 22465 11339 22523 11345
rect 22465 11336 22477 11339
rect 21008 11308 22477 11336
rect 5810 11228 5816 11280
rect 5868 11268 5874 11280
rect 10318 11268 10324 11280
rect 5868 11240 10324 11268
rect 5868 11228 5874 11240
rect 10318 11228 10324 11240
rect 10376 11228 10382 11280
rect 15654 11228 15660 11280
rect 15712 11268 15718 11280
rect 16209 11271 16267 11277
rect 16209 11268 16221 11271
rect 15712 11240 16221 11268
rect 15712 11228 15718 11240
rect 16209 11237 16221 11240
rect 16255 11237 16267 11271
rect 19426 11268 19432 11280
rect 16209 11231 16267 11237
rect 17144 11240 19432 11268
rect 2866 11200 2872 11212
rect 2779 11172 2872 11200
rect 2866 11160 2872 11172
rect 2924 11200 2930 11212
rect 7006 11200 7012 11212
rect 2924 11172 7012 11200
rect 2924 11160 2930 11172
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 7190 11160 7196 11212
rect 7248 11200 7254 11212
rect 9766 11200 9772 11212
rect 7248 11172 8340 11200
rect 7248 11160 7254 11172
rect 5074 11092 5080 11144
rect 5132 11132 5138 11144
rect 7926 11132 7932 11144
rect 5132 11104 7932 11132
rect 5132 11092 5138 11104
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 5445 11067 5503 11073
rect 5445 11033 5457 11067
rect 5491 11064 5503 11067
rect 6914 11064 6920 11076
rect 5491 11036 6920 11064
rect 5491 11033 5503 11036
rect 5445 11027 5503 11033
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 8036 11064 8064 11095
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8312 11141 8340 11172
rect 9324 11172 9772 11200
rect 9324 11141 9352 11172
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 13262 11200 13268 11212
rect 11716 11172 13268 11200
rect 8297 11135 8355 11141
rect 8168 11104 8213 11132
rect 8168 11092 8174 11104
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9490 11132 9496 11144
rect 9451 11104 9496 11132
rect 9309 11095 9367 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 8386 11064 8392 11076
rect 8036 11036 8392 11064
rect 8386 11024 8392 11036
rect 8444 11064 8450 11076
rect 8754 11064 8760 11076
rect 8444 11036 8760 11064
rect 8444 11024 8450 11036
rect 8754 11024 8760 11036
rect 8812 11064 8818 11076
rect 9600 11064 9628 11095
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 9732 11104 10425 11132
rect 9732 11092 9738 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 10413 11095 10471 11101
rect 11054 11092 11060 11104
rect 11112 11132 11118 11144
rect 11716 11141 11744 11172
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 16482 11200 16488 11212
rect 16443 11172 16488 11200
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 11112 11104 11529 11132
rect 11112 11092 11118 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 8812 11036 9628 11064
rect 8812 11024 8818 11036
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 11716 11064 11744 11095
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 14332 11104 14381 11132
rect 14332 11092 14338 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 16574 11132 16580 11144
rect 16535 11104 16580 11132
rect 14369 11095 14427 11101
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 17144 11132 17172 11240
rect 19426 11228 19432 11240
rect 19484 11228 19490 11280
rect 21008 11268 21036 11308
rect 22465 11305 22477 11308
rect 22511 11336 22523 11339
rect 24026 11336 24032 11348
rect 22511 11308 24032 11336
rect 22511 11305 22523 11308
rect 22465 11299 22523 11305
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24210 11296 24216 11348
rect 24268 11336 24274 11348
rect 24397 11339 24455 11345
rect 24397 11336 24409 11339
rect 24268 11308 24409 11336
rect 24268 11296 24274 11308
rect 24397 11305 24409 11308
rect 24443 11305 24455 11339
rect 24397 11299 24455 11305
rect 25682 11296 25688 11348
rect 25740 11336 25746 11348
rect 28353 11339 28411 11345
rect 25740 11308 28304 11336
rect 25740 11296 25746 11308
rect 19904 11240 21036 11268
rect 17221 11203 17279 11209
rect 17221 11169 17233 11203
rect 17267 11200 17279 11203
rect 17267 11172 18276 11200
rect 17267 11169 17279 11172
rect 17221 11163 17279 11169
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 17144 11104 17417 11132
rect 17405 11101 17417 11104
rect 17451 11101 17463 11135
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 17405 11095 17463 11101
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18248 11141 18276 11172
rect 19334 11160 19340 11212
rect 19392 11160 19398 11212
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18322 11092 18328 11144
rect 18380 11132 18386 11144
rect 18506 11141 18512 11144
rect 18463 11135 18512 11141
rect 18380 11104 18425 11132
rect 18380 11092 18386 11104
rect 18463 11101 18475 11135
rect 18509 11101 18512 11135
rect 18463 11095 18512 11101
rect 18506 11092 18512 11095
rect 18564 11092 18570 11144
rect 18966 11092 18972 11144
rect 19024 11132 19030 11144
rect 19352 11132 19380 11160
rect 19904 11141 19932 11240
rect 23474 11228 23480 11280
rect 23532 11228 23538 11280
rect 23842 11228 23848 11280
rect 23900 11228 23906 11280
rect 19889 11135 19947 11141
rect 19024 11104 19748 11132
rect 19024 11092 19030 11104
rect 13354 11064 13360 11076
rect 9916 11036 11744 11064
rect 13315 11036 13360 11064
rect 9916 11024 9922 11036
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 14636 11067 14694 11073
rect 14636 11033 14648 11067
rect 14682 11064 14694 11067
rect 14826 11064 14832 11076
rect 14682 11036 14832 11064
rect 14682 11033 14694 11036
rect 14636 11027 14694 11033
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 18693 11067 18751 11073
rect 18693 11033 18705 11067
rect 18739 11064 18751 11067
rect 19334 11064 19340 11076
rect 18739 11036 19340 11064
rect 18739 11033 18751 11036
rect 18693 11027 18751 11033
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 19720 11073 19748 11104
rect 19889 11101 19901 11135
rect 19935 11101 19947 11135
rect 20530 11132 20536 11144
rect 19889 11095 19947 11101
rect 19996 11104 20536 11132
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 19996 11064 20024 11104
rect 20530 11092 20536 11104
rect 20588 11092 20594 11144
rect 20622 11092 20628 11144
rect 20680 11132 20686 11144
rect 23492 11141 23520 11228
rect 23860 11200 23888 11228
rect 23584 11172 23888 11200
rect 23584 11141 23612 11172
rect 23934 11160 23940 11212
rect 23992 11200 23998 11212
rect 26973 11203 27031 11209
rect 26973 11200 26985 11203
rect 23992 11172 26985 11200
rect 23992 11160 23998 11172
rect 26973 11169 26985 11172
rect 27019 11169 27031 11203
rect 28276 11200 28304 11308
rect 28353 11305 28365 11339
rect 28399 11336 28411 11339
rect 28534 11336 28540 11348
rect 28399 11308 28540 11336
rect 28399 11305 28411 11308
rect 28353 11299 28411 11305
rect 28534 11296 28540 11308
rect 28592 11296 28598 11348
rect 28994 11336 29000 11348
rect 28955 11308 29000 11336
rect 28994 11296 29000 11308
rect 29052 11296 29058 11348
rect 29914 11336 29920 11348
rect 29875 11308 29920 11336
rect 29914 11296 29920 11308
rect 29972 11296 29978 11348
rect 31110 11336 31116 11348
rect 31071 11308 31116 11336
rect 31110 11296 31116 11308
rect 31168 11296 31174 11348
rect 31294 11296 31300 11348
rect 31352 11336 31358 11348
rect 32125 11339 32183 11345
rect 32125 11336 32137 11339
rect 31352 11308 32137 11336
rect 31352 11296 31358 11308
rect 32125 11305 32137 11308
rect 32171 11305 32183 11339
rect 32125 11299 32183 11305
rect 35253 11339 35311 11345
rect 35253 11305 35265 11339
rect 35299 11336 35311 11339
rect 35434 11336 35440 11348
rect 35299 11308 35440 11336
rect 35299 11305 35311 11308
rect 35253 11299 35311 11305
rect 35434 11296 35440 11308
rect 35492 11296 35498 11348
rect 38930 11336 38936 11348
rect 36188 11308 38936 11336
rect 29638 11268 29644 11280
rect 29599 11240 29644 11268
rect 29638 11228 29644 11240
rect 29696 11228 29702 11280
rect 31018 11268 31024 11280
rect 29748 11240 31024 11268
rect 29748 11200 29776 11240
rect 31018 11228 31024 11240
rect 31076 11228 31082 11280
rect 35713 11271 35771 11277
rect 35713 11237 35725 11271
rect 35759 11237 35771 11271
rect 36188 11268 36216 11308
rect 38930 11296 38936 11308
rect 38988 11296 38994 11348
rect 37550 11268 37556 11280
rect 35713 11231 35771 11237
rect 36096 11240 36216 11268
rect 37511 11240 37556 11268
rect 32122 11200 32128 11212
rect 28276 11172 29776 11200
rect 29840 11172 32128 11200
rect 26973 11163 27031 11169
rect 21085 11135 21143 11141
rect 20680 11104 20725 11132
rect 20680 11092 20686 11104
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 23477 11135 23535 11141
rect 21131 11104 23152 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 19751 11036 20024 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20438 11024 20444 11076
rect 20496 11064 20502 11076
rect 21330 11067 21388 11073
rect 21330 11064 21342 11067
rect 20496 11036 21342 11064
rect 20496 11024 20502 11036
rect 21330 11033 21342 11036
rect 21376 11033 21388 11067
rect 21330 11027 21388 11033
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 7653 10999 7711 11005
rect 7653 10996 7665 10999
rect 7616 10968 7665 10996
rect 7616 10956 7622 10968
rect 7653 10965 7665 10968
rect 7699 10965 7711 10999
rect 7653 10959 7711 10965
rect 9953 10999 10011 11005
rect 9953 10965 9965 10999
rect 9999 10996 10011 10999
rect 10042 10996 10048 11008
rect 9999 10968 10048 10996
rect 9999 10965 10011 10968
rect 9953 10959 10011 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 15749 10999 15807 11005
rect 15749 10965 15761 10999
rect 15795 10996 15807 10999
rect 15930 10996 15936 11008
rect 15795 10968 15936 10996
rect 15795 10965 15807 10968
rect 15749 10959 15807 10965
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 22370 10996 22376 11008
rect 18380 10968 22376 10996
rect 18380 10956 18386 10968
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 23124 10996 23152 11104
rect 23477 11101 23489 11135
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 23569 11135 23627 11141
rect 23569 11101 23581 11135
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 23658 11092 23664 11144
rect 23716 11132 23722 11144
rect 23845 11135 23903 11141
rect 23716 11104 23761 11132
rect 23716 11092 23722 11104
rect 23845 11101 23857 11135
rect 23891 11132 23903 11135
rect 24210 11132 24216 11144
rect 23891 11104 24216 11132
rect 23891 11101 23903 11104
rect 23845 11095 23903 11101
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 24762 11092 24768 11144
rect 24820 11132 24826 11144
rect 24949 11135 25007 11141
rect 24949 11132 24961 11135
rect 24820 11104 24961 11132
rect 24820 11092 24826 11104
rect 24949 11101 24961 11104
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11132 25283 11135
rect 25314 11132 25320 11144
rect 25271 11104 25320 11132
rect 25271 11101 25283 11104
rect 25225 11095 25283 11101
rect 25314 11092 25320 11104
rect 25372 11092 25378 11144
rect 27240 11135 27298 11141
rect 27240 11101 27252 11135
rect 27286 11132 27298 11135
rect 27614 11132 27620 11144
rect 27286 11104 27620 11132
rect 27286 11101 27298 11104
rect 27240 11095 27298 11101
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 29840 11141 29868 11172
rect 32122 11160 32128 11172
rect 32180 11160 32186 11212
rect 35728 11200 35756 11231
rect 32416 11172 35756 11200
rect 29825 11135 29883 11141
rect 29825 11101 29837 11135
rect 29871 11101 29883 11135
rect 29825 11095 29883 11101
rect 29914 11092 29920 11144
rect 29972 11132 29978 11144
rect 29972 11104 30017 11132
rect 29972 11092 29978 11104
rect 31202 11092 31208 11144
rect 31260 11132 31266 11144
rect 31297 11135 31355 11141
rect 31297 11132 31309 11135
rect 31260 11104 31309 11132
rect 31260 11092 31266 11104
rect 31297 11101 31309 11104
rect 31343 11101 31355 11135
rect 31297 11095 31355 11101
rect 31386 11092 31392 11144
rect 31444 11132 31450 11144
rect 31662 11132 31668 11144
rect 31444 11104 31489 11132
rect 31623 11104 31668 11132
rect 31444 11092 31450 11104
rect 31662 11092 31668 11104
rect 31720 11092 31726 11144
rect 32416 11141 32444 11172
rect 32309 11135 32367 11141
rect 32309 11101 32321 11135
rect 32355 11101 32367 11135
rect 32309 11095 32367 11101
rect 32401 11135 32459 11141
rect 32401 11101 32413 11135
rect 32447 11101 32459 11135
rect 32674 11132 32680 11144
rect 32635 11104 32680 11132
rect 32401 11095 32459 11101
rect 23201 11067 23259 11073
rect 23201 11033 23213 11067
rect 23247 11064 23259 11067
rect 24026 11064 24032 11076
rect 23247 11036 24032 11064
rect 23247 11033 23259 11036
rect 23201 11027 23259 11033
rect 24026 11024 24032 11036
rect 24084 11024 24090 11076
rect 24118 11024 24124 11076
rect 24176 11064 24182 11076
rect 30101 11067 30159 11073
rect 30101 11064 30113 11067
rect 24176 11036 30113 11064
rect 24176 11024 24182 11036
rect 30101 11033 30113 11036
rect 30147 11064 30159 11067
rect 30561 11067 30619 11073
rect 30561 11064 30573 11067
rect 30147 11036 30573 11064
rect 30147 11033 30159 11036
rect 30101 11027 30159 11033
rect 30561 11033 30573 11036
rect 30607 11033 30619 11067
rect 30561 11027 30619 11033
rect 31481 11067 31539 11073
rect 31481 11033 31493 11067
rect 31527 11033 31539 11067
rect 31481 11027 31539 11033
rect 23934 10996 23940 11008
rect 23124 10968 23940 10996
rect 23934 10956 23940 10968
rect 23992 10956 23998 11008
rect 31386 10956 31392 11008
rect 31444 10996 31450 11008
rect 31496 10996 31524 11027
rect 31570 11024 31576 11076
rect 31628 11064 31634 11076
rect 32324 11064 32352 11095
rect 32674 11092 32680 11104
rect 32732 11092 32738 11144
rect 33410 11092 33416 11144
rect 33468 11132 33474 11144
rect 33873 11135 33931 11141
rect 33873 11132 33885 11135
rect 33468 11104 33885 11132
rect 33468 11092 33474 11104
rect 33873 11101 33885 11104
rect 33919 11101 33931 11135
rect 33873 11095 33931 11101
rect 34149 11135 34207 11141
rect 34149 11101 34161 11135
rect 34195 11132 34207 11135
rect 34422 11132 34428 11144
rect 34195 11104 34428 11132
rect 34195 11101 34207 11104
rect 34149 11095 34207 11101
rect 32490 11064 32496 11076
rect 31628 11036 32352 11064
rect 32451 11036 32496 11064
rect 31628 11024 31634 11036
rect 32490 11024 32496 11036
rect 32548 11024 32554 11076
rect 33888 11064 33916 11095
rect 34422 11092 34428 11104
rect 34480 11092 34486 11144
rect 34698 11092 34704 11144
rect 34756 11132 34762 11144
rect 35084 11141 35112 11172
rect 34885 11135 34943 11141
rect 34885 11132 34897 11135
rect 34756 11104 34897 11132
rect 34756 11092 34762 11104
rect 34885 11101 34897 11104
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11101 35127 11135
rect 35069 11095 35127 11101
rect 36096 11064 36124 11240
rect 37550 11228 37556 11240
rect 37608 11228 37614 11280
rect 38933 11203 38991 11209
rect 38933 11200 38945 11203
rect 38856 11172 38945 11200
rect 38856 11144 38884 11172
rect 38933 11169 38945 11172
rect 38979 11200 38991 11203
rect 39114 11200 39120 11212
rect 38979 11172 39120 11200
rect 38979 11169 38991 11172
rect 38933 11163 38991 11169
rect 39114 11160 39120 11172
rect 39172 11160 39178 11212
rect 40402 11200 40408 11212
rect 40144 11172 40408 11200
rect 40144 11144 40172 11172
rect 40402 11160 40408 11172
rect 40460 11160 40466 11212
rect 37090 11132 37096 11144
rect 36740 11104 37096 11132
rect 36740 11076 36768 11104
rect 37090 11092 37096 11104
rect 37148 11092 37154 11144
rect 38838 11092 38844 11144
rect 38896 11092 38902 11144
rect 40126 11132 40132 11144
rect 40087 11104 40132 11132
rect 40126 11092 40132 11104
rect 40184 11092 40190 11144
rect 40221 11135 40279 11141
rect 40221 11101 40233 11135
rect 40267 11101 40279 11135
rect 40221 11095 40279 11101
rect 33888 11036 36124 11064
rect 36722 11024 36728 11076
rect 36780 11024 36786 11076
rect 36814 11024 36820 11076
rect 36872 11073 36878 11076
rect 36872 11064 36884 11073
rect 38688 11067 38746 11073
rect 36872 11036 36917 11064
rect 36872 11027 36884 11036
rect 38688 11033 38700 11067
rect 38734 11064 38746 11067
rect 39853 11067 39911 11073
rect 39853 11064 39865 11067
rect 38734 11036 39865 11064
rect 38734 11033 38746 11036
rect 38688 11027 38746 11033
rect 39853 11033 39865 11036
rect 39899 11033 39911 11067
rect 39853 11027 39911 11033
rect 36872 11024 36878 11027
rect 40236 11008 40264 11095
rect 40310 11092 40316 11144
rect 40368 11132 40374 11144
rect 40368 11104 40413 11132
rect 40368 11092 40374 11104
rect 40494 11092 40500 11144
rect 40552 11132 40558 11144
rect 40552 11104 40597 11132
rect 40552 11092 40558 11104
rect 31444 10968 31524 10996
rect 31444 10956 31450 10968
rect 35710 10956 35716 11008
rect 35768 10996 35774 11008
rect 40218 10996 40224 11008
rect 35768 10968 40224 10996
rect 35768 10956 35774 10968
rect 40218 10956 40224 10968
rect 40276 10956 40282 11008
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 2593 10795 2651 10801
rect 2593 10792 2605 10795
rect 1912 10764 2605 10792
rect 1912 10752 1918 10764
rect 2593 10761 2605 10764
rect 2639 10792 2651 10795
rect 3142 10792 3148 10804
rect 2639 10764 3148 10792
rect 2639 10761 2651 10764
rect 2593 10755 2651 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 5810 10792 5816 10804
rect 5771 10764 5816 10792
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 8110 10792 8116 10804
rect 6503 10764 8116 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9309 10795 9367 10801
rect 9309 10761 9321 10795
rect 9355 10792 9367 10795
rect 9490 10792 9496 10804
rect 9355 10764 9496 10792
rect 9355 10761 9367 10764
rect 9309 10755 9367 10761
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 13541 10795 13599 10801
rect 13541 10792 13553 10795
rect 12584 10764 13553 10792
rect 12584 10752 12590 10764
rect 13541 10761 13553 10764
rect 13587 10792 13599 10795
rect 18322 10792 18328 10804
rect 13587 10764 18328 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 20162 10792 20168 10804
rect 19576 10764 20168 10792
rect 19576 10752 19582 10764
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 23293 10795 23351 10801
rect 20680 10764 23244 10792
rect 20680 10752 20686 10764
rect 1394 10724 1400 10736
rect 1355 10696 1400 10724
rect 1394 10684 1400 10696
rect 1452 10684 1458 10736
rect 1581 10727 1639 10733
rect 1581 10693 1593 10727
rect 1627 10724 1639 10727
rect 5258 10724 5264 10736
rect 1627 10696 5264 10724
rect 1627 10693 1639 10696
rect 1581 10687 1639 10693
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 8938 10724 8944 10736
rect 6604 10696 8944 10724
rect 6604 10684 6610 10696
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3706 10659 3764 10665
rect 3706 10656 3718 10659
rect 3200 10628 3718 10656
rect 3200 10616 3206 10628
rect 3706 10625 3718 10628
rect 3752 10625 3764 10659
rect 3970 10656 3976 10668
rect 3931 10628 3976 10656
rect 3706 10619 3764 10625
rect 3970 10616 3976 10628
rect 4028 10656 4034 10668
rect 4706 10665 4712 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4028 10628 4445 10656
rect 4028 10616 4034 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4700 10656 4712 10665
rect 4667 10628 4712 10656
rect 4433 10619 4491 10625
rect 4700 10619 4712 10628
rect 4706 10616 4712 10619
rect 4764 10616 4770 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 7006 10656 7012 10668
rect 6871 10628 7012 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 6656 10452 6684 10619
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7300 10665 7328 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 11698 10724 11704 10736
rect 11659 10696 11704 10724
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 13630 10684 13636 10736
rect 13688 10724 13694 10736
rect 23106 10724 23112 10736
rect 13688 10696 18828 10724
rect 13688 10684 13694 10696
rect 7558 10665 7564 10668
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7552 10656 7564 10665
rect 7519 10628 7564 10656
rect 7285 10619 7343 10625
rect 7552 10619 7564 10628
rect 7558 10616 7564 10619
rect 7616 10616 7622 10668
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 9493 10619 9551 10625
rect 9508 10588 9536 10619
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11112 10628 11529 10656
rect 11112 10616 11118 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11790 10656 11796 10668
rect 11751 10628 11796 10656
rect 11517 10619 11575 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 11940 10628 11985 10656
rect 11940 10616 11946 10628
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 13354 10656 13360 10668
rect 12492 10628 13360 10656
rect 12492 10616 12498 10628
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 14090 10656 14096 10668
rect 14051 10628 14096 10656
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 14182 10616 14188 10668
rect 14240 10656 14246 10668
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 14240 10628 14289 10656
rect 14240 10616 14246 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 14645 10659 14703 10665
rect 14424 10628 14469 10656
rect 14424 10616 14430 10628
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 15930 10656 15936 10668
rect 14691 10628 15936 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 17310 10656 17316 10668
rect 17271 10628 17316 10656
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18230 10656 18236 10668
rect 18187 10628 18236 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18230 10616 18236 10628
rect 18288 10656 18294 10668
rect 18506 10656 18512 10668
rect 18288 10628 18512 10656
rect 18288 10616 18294 10628
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 11330 10588 11336 10600
rect 9508 10560 11336 10588
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10588 14519 10591
rect 15470 10588 15476 10600
rect 14507 10560 15476 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 15470 10548 15476 10560
rect 15528 10548 15534 10600
rect 17218 10588 17224 10600
rect 17179 10560 17224 10588
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 18800 10588 18828 10696
rect 18892 10696 23112 10724
rect 18892 10665 18920 10696
rect 23106 10684 23112 10696
rect 23164 10684 23170 10736
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10656 19027 10659
rect 19518 10656 19524 10668
rect 19015 10628 19524 10656
rect 19015 10625 19027 10628
rect 18969 10619 19027 10625
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 19150 10588 19156 10600
rect 18800 10560 19156 10588
rect 19150 10548 19156 10560
rect 19208 10588 19214 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19208 10560 19441 10588
rect 19208 10548 19214 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 12066 10520 12072 10532
rect 12027 10492 12072 10520
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 12250 10480 12256 10532
rect 12308 10520 12314 10532
rect 19444 10520 19472 10551
rect 19518 10520 19524 10532
rect 12308 10492 17172 10520
rect 19444 10492 19524 10520
rect 12308 10480 12314 10492
rect 8665 10455 8723 10461
rect 8665 10452 8677 10455
rect 6656 10424 8677 10452
rect 8665 10421 8677 10424
rect 8711 10452 8723 10455
rect 9030 10452 9036 10464
rect 8711 10424 9036 10452
rect 8711 10421 8723 10424
rect 8665 10415 8723 10421
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 14826 10452 14832 10464
rect 14787 10424 14832 10452
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 16945 10455 17003 10461
rect 16945 10421 16957 10455
rect 16991 10452 17003 10455
rect 17034 10452 17040 10464
rect 16991 10424 17040 10452
rect 16991 10421 17003 10424
rect 16945 10415 17003 10421
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 17144 10461 17172 10492
rect 19518 10480 19524 10492
rect 19576 10480 19582 10532
rect 19628 10520 19656 10619
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20533 10659 20591 10665
rect 20533 10656 20545 10659
rect 20128 10628 20545 10656
rect 20128 10616 20134 10628
rect 20533 10625 20545 10628
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 20990 10616 20996 10668
rect 21048 10656 21054 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21048 10628 21833 10656
rect 21048 10616 21054 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10656 22063 10659
rect 22370 10656 22376 10668
rect 22051 10628 22376 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 22370 10616 22376 10628
rect 22428 10656 22434 10668
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 22428 10628 22477 10656
rect 22428 10616 22434 10628
rect 22465 10625 22477 10628
rect 22511 10625 22523 10659
rect 22465 10619 22523 10625
rect 20257 10591 20315 10597
rect 20257 10557 20269 10591
rect 20303 10588 20315 10591
rect 23216 10588 23244 10764
rect 23293 10761 23305 10795
rect 23339 10792 23351 10795
rect 23474 10792 23480 10804
rect 23339 10764 23480 10792
rect 23339 10761 23351 10764
rect 23293 10755 23351 10761
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 24670 10752 24676 10804
rect 24728 10792 24734 10804
rect 27522 10792 27528 10804
rect 24728 10764 27528 10792
rect 24728 10752 24734 10764
rect 27522 10752 27528 10764
rect 27580 10752 27586 10804
rect 30006 10792 30012 10804
rect 29967 10764 30012 10792
rect 30006 10752 30012 10764
rect 30064 10752 30070 10804
rect 30561 10795 30619 10801
rect 30561 10761 30573 10795
rect 30607 10792 30619 10795
rect 30650 10792 30656 10804
rect 30607 10764 30656 10792
rect 30607 10761 30619 10764
rect 30561 10755 30619 10761
rect 30650 10752 30656 10764
rect 30708 10752 30714 10804
rect 31021 10795 31079 10801
rect 31021 10761 31033 10795
rect 31067 10761 31079 10795
rect 32122 10792 32128 10804
rect 32083 10764 32128 10792
rect 31021 10755 31079 10761
rect 26694 10684 26700 10736
rect 26752 10724 26758 10736
rect 26752 10696 27476 10724
rect 26752 10684 26758 10696
rect 23750 10656 23756 10668
rect 23711 10628 23756 10656
rect 23750 10616 23756 10628
rect 23808 10616 23814 10668
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 24670 10656 24676 10668
rect 23900 10628 24676 10656
rect 23900 10616 23906 10628
rect 24670 10616 24676 10628
rect 24728 10616 24734 10668
rect 24946 10656 24952 10668
rect 24907 10628 24952 10656
rect 24946 10616 24952 10628
rect 25004 10616 25010 10668
rect 27448 10665 27476 10696
rect 27433 10659 27491 10665
rect 27433 10625 27445 10659
rect 27479 10625 27491 10659
rect 29546 10656 29552 10668
rect 29507 10628 29552 10656
rect 27433 10619 27491 10625
rect 29546 10616 29552 10628
rect 29604 10616 29610 10668
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10656 29883 10659
rect 31036 10656 31064 10755
rect 32122 10752 32128 10764
rect 32180 10752 32186 10804
rect 38654 10792 38660 10804
rect 32600 10764 38660 10792
rect 31386 10724 31392 10736
rect 31347 10696 31392 10724
rect 31386 10684 31392 10696
rect 31444 10724 31450 10736
rect 32490 10724 32496 10736
rect 31444 10696 32496 10724
rect 31444 10684 31450 10696
rect 32490 10684 32496 10696
rect 32548 10684 32554 10736
rect 31202 10656 31208 10668
rect 29871 10628 31064 10656
rect 31115 10628 31208 10656
rect 29871 10625 29883 10628
rect 29825 10619 29883 10625
rect 31202 10616 31208 10628
rect 31260 10616 31266 10668
rect 31294 10616 31300 10668
rect 31352 10656 31358 10668
rect 31573 10659 31631 10665
rect 31352 10628 31397 10656
rect 31352 10616 31358 10628
rect 31573 10625 31585 10659
rect 31619 10656 31631 10659
rect 32214 10656 32220 10668
rect 31619 10628 32220 10656
rect 31619 10625 31631 10628
rect 31573 10619 31631 10625
rect 32214 10616 32220 10628
rect 32272 10616 32278 10668
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32401 10659 32459 10665
rect 32401 10625 32413 10659
rect 32447 10656 32459 10659
rect 32600 10656 32628 10764
rect 38654 10752 38660 10764
rect 38712 10752 38718 10804
rect 39577 10795 39635 10801
rect 39577 10761 39589 10795
rect 39623 10792 39635 10795
rect 40310 10792 40316 10804
rect 39623 10764 40316 10792
rect 39623 10761 39635 10764
rect 39577 10755 39635 10761
rect 40310 10752 40316 10764
rect 40368 10752 40374 10804
rect 34330 10724 34336 10736
rect 32692 10696 34336 10724
rect 32692 10665 32720 10696
rect 34330 10684 34336 10696
rect 34388 10684 34394 10736
rect 34606 10684 34612 10736
rect 34664 10724 34670 10736
rect 35529 10727 35587 10733
rect 35529 10724 35541 10727
rect 34664 10696 35541 10724
rect 34664 10684 34670 10696
rect 35529 10693 35541 10696
rect 35575 10693 35587 10727
rect 35529 10687 35587 10693
rect 36265 10727 36323 10733
rect 36265 10693 36277 10727
rect 36311 10724 36323 10727
rect 36354 10724 36360 10736
rect 36311 10696 36360 10724
rect 36311 10693 36323 10696
rect 36265 10687 36323 10693
rect 36354 10684 36360 10696
rect 36412 10684 36418 10736
rect 37550 10684 37556 10736
rect 37608 10724 37614 10736
rect 39393 10727 39451 10733
rect 39393 10724 39405 10727
rect 37608 10696 39405 10724
rect 37608 10684 37614 10696
rect 39393 10693 39405 10696
rect 39439 10693 39451 10727
rect 40126 10724 40132 10736
rect 40087 10696 40132 10724
rect 39393 10687 39451 10693
rect 40126 10684 40132 10696
rect 40184 10684 40190 10736
rect 32447 10628 32628 10656
rect 32677 10659 32735 10665
rect 32447 10625 32459 10628
rect 32401 10619 32459 10625
rect 32677 10625 32689 10659
rect 32723 10625 32735 10659
rect 33318 10656 33324 10668
rect 33279 10628 33324 10656
rect 32677 10619 32735 10625
rect 28442 10588 28448 10600
rect 20303 10560 20944 10588
rect 23216 10560 28448 10588
rect 20303 10557 20315 10560
rect 20257 10551 20315 10557
rect 20916 10532 20944 10560
rect 28442 10548 28448 10560
rect 28500 10548 28506 10600
rect 28994 10548 29000 10600
rect 29052 10588 29058 10600
rect 29641 10591 29699 10597
rect 29641 10588 29653 10591
rect 29052 10560 29653 10588
rect 29052 10548 29058 10560
rect 29641 10557 29653 10560
rect 29687 10557 29699 10591
rect 31220 10588 31248 10616
rect 32324 10588 32352 10619
rect 33318 10616 33324 10628
rect 33376 10616 33382 10668
rect 34146 10656 34152 10668
rect 34107 10628 34152 10656
rect 34146 10616 34152 10628
rect 34204 10616 34210 10668
rect 34425 10659 34483 10665
rect 34425 10625 34437 10659
rect 34471 10656 34483 10659
rect 34698 10656 34704 10668
rect 34471 10628 34704 10656
rect 34471 10625 34483 10628
rect 34425 10619 34483 10625
rect 34698 10616 34704 10628
rect 34756 10616 34762 10668
rect 38930 10616 38936 10668
rect 38988 10656 38994 10668
rect 39209 10659 39267 10665
rect 39209 10656 39221 10659
rect 38988 10628 39221 10656
rect 38988 10616 38994 10628
rect 39209 10625 39221 10628
rect 39255 10656 39267 10659
rect 39942 10656 39948 10668
rect 39255 10628 39948 10656
rect 39255 10625 39267 10628
rect 39209 10619 39267 10625
rect 39942 10616 39948 10628
rect 40000 10616 40006 10668
rect 33137 10591 33195 10597
rect 33137 10588 33149 10591
rect 31220 10560 32352 10588
rect 32416 10560 33149 10588
rect 29641 10551 29699 10557
rect 31588 10532 31616 10560
rect 20806 10520 20812 10532
rect 19628 10492 20812 10520
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 20898 10480 20904 10532
rect 20956 10520 20962 10532
rect 21913 10523 21971 10529
rect 21913 10520 21925 10523
rect 20956 10492 21925 10520
rect 20956 10480 20962 10492
rect 21913 10489 21925 10492
rect 21959 10489 21971 10523
rect 21913 10483 21971 10489
rect 27614 10480 27620 10532
rect 27672 10520 27678 10532
rect 27672 10492 27717 10520
rect 27672 10480 27678 10492
rect 31570 10480 31576 10532
rect 31628 10480 31634 10532
rect 17129 10455 17187 10461
rect 17129 10421 17141 10455
rect 17175 10421 17187 10455
rect 17129 10415 17187 10421
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18601 10455 18659 10461
rect 18601 10452 18613 10455
rect 18196 10424 18613 10452
rect 18196 10412 18202 10424
rect 18601 10421 18613 10424
rect 18647 10421 18659 10455
rect 18782 10452 18788 10464
rect 18743 10424 18788 10452
rect 18601 10415 18659 10421
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 19797 10455 19855 10461
rect 19797 10421 19809 10455
rect 19843 10452 19855 10455
rect 21082 10452 21088 10464
rect 19843 10424 21088 10452
rect 19843 10421 19855 10424
rect 19797 10415 19855 10421
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 23937 10455 23995 10461
rect 23937 10421 23949 10455
rect 23983 10452 23995 10455
rect 24210 10452 24216 10464
rect 23983 10424 24216 10452
rect 23983 10421 23995 10424
rect 23937 10415 23995 10421
rect 24210 10412 24216 10424
rect 24268 10412 24274 10464
rect 26421 10455 26479 10461
rect 26421 10421 26433 10455
rect 26467 10452 26479 10455
rect 26694 10452 26700 10464
rect 26467 10424 26700 10452
rect 26467 10421 26479 10424
rect 26421 10415 26479 10421
rect 26694 10412 26700 10424
rect 26752 10412 26758 10464
rect 29825 10455 29883 10461
rect 29825 10421 29837 10455
rect 29871 10452 29883 10455
rect 30374 10452 30380 10464
rect 29871 10424 30380 10452
rect 29871 10421 29883 10424
rect 29825 10415 29883 10421
rect 30374 10412 30380 10424
rect 30432 10412 30438 10464
rect 30650 10412 30656 10464
rect 30708 10452 30714 10464
rect 32416 10452 32444 10560
rect 33137 10557 33149 10560
rect 33183 10557 33195 10591
rect 33137 10551 33195 10557
rect 35713 10591 35771 10597
rect 35713 10557 35725 10591
rect 35759 10588 35771 10591
rect 36446 10588 36452 10600
rect 35759 10560 36452 10588
rect 35759 10557 35771 10560
rect 35713 10551 35771 10557
rect 36446 10548 36452 10560
rect 36504 10548 36510 10600
rect 30708 10424 32444 10452
rect 33505 10455 33563 10461
rect 30708 10412 30714 10424
rect 33505 10421 33517 10455
rect 33551 10452 33563 10455
rect 34422 10452 34428 10464
rect 33551 10424 34428 10452
rect 33551 10421 33563 10424
rect 33505 10415 33563 10421
rect 34422 10412 34428 10424
rect 34480 10412 34486 10464
rect 36354 10412 36360 10464
rect 36412 10452 36418 10464
rect 39758 10452 39764 10464
rect 36412 10424 39764 10452
rect 36412 10412 36418 10424
rect 39758 10412 39764 10424
rect 39816 10412 39822 10464
rect 67634 10452 67640 10464
rect 67595 10424 67640 10452
rect 67634 10412 67640 10424
rect 67692 10412 67698 10464
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 3053 10251 3111 10257
rect 3053 10217 3065 10251
rect 3099 10248 3111 10251
rect 3142 10248 3148 10260
rect 3099 10220 3148 10248
rect 3099 10217 3111 10220
rect 3053 10211 3111 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7248 10220 7481 10248
rect 7248 10208 7254 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 7469 10211 7527 10217
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 19426 10208 19432 10260
rect 19484 10248 19490 10260
rect 20622 10248 20628 10260
rect 19484 10220 20628 10248
rect 19484 10208 19490 10220
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 22005 10251 22063 10257
rect 22005 10248 22017 10251
rect 21876 10220 22017 10248
rect 21876 10208 21882 10220
rect 22005 10217 22017 10220
rect 22051 10217 22063 10251
rect 22005 10211 22063 10217
rect 27525 10251 27583 10257
rect 27525 10217 27537 10251
rect 27571 10217 27583 10251
rect 28994 10248 29000 10260
rect 28955 10220 29000 10248
rect 27525 10211 27583 10217
rect 14090 10140 14096 10192
rect 14148 10180 14154 10192
rect 27540 10180 27568 10211
rect 28994 10208 29000 10220
rect 29052 10208 29058 10260
rect 29914 10208 29920 10260
rect 29972 10248 29978 10260
rect 30101 10251 30159 10257
rect 30101 10248 30113 10251
rect 29972 10220 30113 10248
rect 29972 10208 29978 10220
rect 30101 10217 30113 10220
rect 30147 10217 30159 10251
rect 35710 10248 35716 10260
rect 35671 10220 35716 10248
rect 30101 10211 30159 10217
rect 35710 10208 35716 10220
rect 35768 10208 35774 10260
rect 30558 10180 30564 10192
rect 14148 10152 15792 10180
rect 27540 10152 30564 10180
rect 14148 10140 14154 10152
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 1995 10084 2636 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 1394 10004 1400 10056
rect 1452 10044 1458 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 1452 10016 1593 10044
rect 1452 10004 1458 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10044 1823 10047
rect 1854 10044 1860 10056
rect 1811 10016 1860 10044
rect 1811 10013 1823 10016
rect 1765 10007 1823 10013
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 2038 10004 2044 10056
rect 2096 10044 2102 10056
rect 2608 10053 2636 10084
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 8018 10112 8024 10124
rect 7064 10084 8024 10112
rect 7064 10072 7070 10084
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8938 10072 8944 10124
rect 8996 10112 9002 10124
rect 9953 10115 10011 10121
rect 9953 10112 9965 10115
rect 8996 10084 9965 10112
rect 8996 10072 9002 10084
rect 9953 10081 9965 10084
rect 9999 10081 10011 10115
rect 15565 10115 15623 10121
rect 15565 10112 15577 10115
rect 9953 10075 10011 10081
rect 13464 10084 15577 10112
rect 2409 10047 2467 10053
rect 2409 10044 2421 10047
rect 2096 10016 2421 10044
rect 2096 10004 2102 10016
rect 2409 10013 2421 10016
rect 2455 10013 2467 10047
rect 2409 10007 2467 10013
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10013 2743 10047
rect 2685 10007 2743 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 2823 10016 3801 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3789 10013 3801 10016
rect 3835 10044 3847 10047
rect 5074 10044 5080 10056
rect 3835 10016 5080 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 2700 9976 2728 10007
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10209 10047 10267 10053
rect 10209 10044 10221 10047
rect 10100 10016 10221 10044
rect 10100 10004 10106 10016
rect 10209 10013 10221 10016
rect 10255 10013 10267 10047
rect 13464 10044 13492 10084
rect 15565 10081 15577 10084
rect 15611 10081 15623 10115
rect 15565 10075 15623 10081
rect 10209 10007 10267 10013
rect 12406 10016 13492 10044
rect 13541 10047 13599 10053
rect 2608 9948 2728 9976
rect 2608 9920 2636 9948
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 12406 9976 12434 10016
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 14274 10044 14280 10056
rect 13587 10016 14280 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 15470 10044 15476 10056
rect 15431 10016 15476 10044
rect 15289 10007 15347 10013
rect 8352 9948 12434 9976
rect 13296 9979 13354 9985
rect 8352 9936 8358 9948
rect 13296 9945 13308 9979
rect 13342 9976 13354 9979
rect 13446 9976 13452 9988
rect 13342 9948 13452 9976
rect 13342 9945 13354 9948
rect 13296 9939 13354 9945
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 15304 9976 15332 10007
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 15654 10044 15660 10056
rect 15615 10016 15660 10044
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 15764 10044 15792 10152
rect 30558 10140 30564 10152
rect 30616 10140 30622 10192
rect 31294 10140 31300 10192
rect 31352 10180 31358 10192
rect 38286 10180 38292 10192
rect 31352 10152 38292 10180
rect 31352 10140 31358 10152
rect 38286 10140 38292 10152
rect 38344 10140 38350 10192
rect 40218 10140 40224 10192
rect 40276 10140 40282 10192
rect 16390 10072 16396 10124
rect 16448 10112 16454 10124
rect 17313 10115 17371 10121
rect 17313 10112 17325 10115
rect 16448 10084 17325 10112
rect 16448 10072 16454 10084
rect 17313 10081 17325 10084
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 17460 10084 19257 10112
rect 17460 10072 17466 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 19245 10075 19303 10081
rect 23845 10115 23903 10121
rect 23845 10081 23857 10115
rect 23891 10112 23903 10115
rect 23934 10112 23940 10124
rect 23891 10084 23940 10112
rect 23891 10081 23903 10084
rect 23845 10075 23903 10081
rect 23934 10072 23940 10084
rect 23992 10072 23998 10124
rect 24670 10112 24676 10124
rect 24631 10084 24676 10112
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 27338 10112 27344 10124
rect 27299 10084 27344 10112
rect 27338 10072 27344 10084
rect 27396 10072 27402 10124
rect 28902 10112 28908 10124
rect 27448 10084 28908 10112
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 15764 10016 15853 10044
rect 15841 10013 15853 10016
rect 15887 10044 15899 10047
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 15887 10016 16957 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 16945 10013 16957 10016
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 17092 10016 17141 10044
rect 17092 10004 17098 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10013 17279 10047
rect 17494 10044 17500 10056
rect 17455 10016 17500 10044
rect 17221 10007 17279 10013
rect 16114 9976 16120 9988
rect 15304 9948 16120 9976
rect 16114 9936 16120 9948
rect 16172 9936 16178 9988
rect 17236 9976 17264 10007
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19501 10047 19559 10053
rect 19501 10044 19513 10047
rect 19392 10016 19513 10044
rect 19392 10004 19398 10016
rect 19501 10013 19513 10016
rect 19547 10013 19559 10047
rect 21450 10044 21456 10056
rect 21411 10016 21456 10044
rect 19501 10007 19559 10013
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 21821 10047 21879 10053
rect 21821 10013 21833 10047
rect 21867 10044 21879 10047
rect 21910 10044 21916 10056
rect 21867 10016 21916 10044
rect 21867 10013 21879 10016
rect 21821 10007 21879 10013
rect 21910 10004 21916 10016
rect 21968 10004 21974 10056
rect 23578 10047 23636 10053
rect 23578 10013 23590 10047
rect 23624 10044 23636 10047
rect 24026 10044 24032 10056
rect 23624 10016 24032 10044
rect 23624 10013 23636 10016
rect 23578 10007 23636 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10044 25007 10047
rect 25222 10044 25228 10056
rect 24995 10016 25228 10044
rect 24995 10013 25007 10016
rect 24949 10007 25007 10013
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 25682 10004 25688 10056
rect 25740 10044 25746 10056
rect 25961 10047 26019 10053
rect 25961 10044 25973 10047
rect 25740 10016 25973 10044
rect 25740 10004 25746 10016
rect 25961 10013 25973 10016
rect 26007 10013 26019 10047
rect 26234 10044 26240 10056
rect 26195 10016 26240 10044
rect 25961 10007 26019 10013
rect 26234 10004 26240 10016
rect 26292 10044 26298 10056
rect 27448 10044 27476 10084
rect 26292 10016 27476 10044
rect 27525 10047 27583 10053
rect 26292 10004 26298 10016
rect 27525 10013 27537 10047
rect 27571 10044 27583 10047
rect 28350 10044 28356 10056
rect 27571 10016 28356 10044
rect 27571 10013 27583 10016
rect 27525 10007 27583 10013
rect 28350 10004 28356 10016
rect 28408 10004 28414 10056
rect 28828 10053 28856 10084
rect 28902 10072 28908 10084
rect 28960 10112 28966 10124
rect 28960 10084 29960 10112
rect 28960 10072 28966 10084
rect 28445 10047 28503 10053
rect 28445 10013 28457 10047
rect 28491 10013 28503 10047
rect 28445 10007 28503 10013
rect 28813 10047 28871 10053
rect 28813 10013 28825 10047
rect 28859 10044 28871 10047
rect 28859 10016 28893 10044
rect 28859 10013 28871 10016
rect 28813 10007 28871 10013
rect 17954 9976 17960 9988
rect 17236 9948 17960 9976
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 21358 9936 21364 9988
rect 21416 9976 21422 9988
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 21416 9948 21649 9976
rect 21416 9936 21422 9948
rect 21637 9945 21649 9948
rect 21683 9945 21695 9979
rect 21637 9939 21695 9945
rect 21729 9979 21787 9985
rect 21729 9945 21741 9979
rect 21775 9976 21787 9979
rect 27246 9976 27252 9988
rect 21775 9948 22094 9976
rect 27207 9948 27252 9976
rect 21775 9945 21787 9948
rect 21729 9939 21787 9945
rect 2590 9868 2596 9920
rect 2648 9868 2654 9920
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 9640 9880 12173 9908
rect 9640 9868 9646 9880
rect 12161 9877 12173 9880
rect 12207 9908 12219 9911
rect 13170 9908 13176 9920
rect 12207 9880 13176 9908
rect 12207 9877 12219 9880
rect 12161 9871 12219 9877
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 15105 9911 15163 9917
rect 15105 9908 15117 9911
rect 15068 9880 15117 9908
rect 15068 9868 15074 9880
rect 15105 9877 15117 9880
rect 15151 9877 15163 9911
rect 15105 9871 15163 9877
rect 17681 9911 17739 9917
rect 17681 9877 17693 9911
rect 17727 9908 17739 9911
rect 18322 9908 18328 9920
rect 17727 9880 18328 9908
rect 17727 9877 17739 9880
rect 17681 9871 17739 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 22066 9908 22094 9948
rect 27246 9936 27252 9948
rect 27304 9936 27310 9988
rect 22465 9911 22523 9917
rect 22465 9908 22477 9911
rect 22066 9880 22477 9908
rect 22465 9877 22477 9880
rect 22511 9908 22523 9911
rect 22554 9908 22560 9920
rect 22511 9880 22560 9908
rect 22511 9877 22523 9880
rect 22465 9871 22523 9877
rect 22554 9868 22560 9880
rect 22612 9868 22618 9920
rect 23106 9868 23112 9920
rect 23164 9908 23170 9920
rect 27709 9911 27767 9917
rect 27709 9908 27721 9911
rect 23164 9880 27721 9908
rect 23164 9868 23170 9880
rect 27709 9877 27721 9880
rect 27755 9877 27767 9911
rect 28460 9908 28488 10007
rect 29454 10004 29460 10056
rect 29512 10044 29518 10056
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 29512 10016 29561 10044
rect 29512 10004 29518 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29822 10044 29828 10056
rect 29783 10016 29828 10044
rect 29549 10007 29607 10013
rect 29822 10004 29828 10016
rect 29880 10004 29886 10056
rect 29932 10053 29960 10084
rect 33134 10072 33140 10124
rect 33192 10112 33198 10124
rect 33229 10115 33287 10121
rect 33229 10112 33241 10115
rect 33192 10084 33241 10112
rect 33192 10072 33198 10084
rect 33229 10081 33241 10084
rect 33275 10081 33287 10115
rect 33229 10075 33287 10081
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 31570 10004 31576 10056
rect 31628 10044 31634 10056
rect 31849 10047 31907 10053
rect 31849 10044 31861 10047
rect 31628 10016 31861 10044
rect 31628 10004 31634 10016
rect 31849 10013 31861 10016
rect 31895 10013 31907 10047
rect 31849 10007 31907 10013
rect 32125 10047 32183 10053
rect 32125 10013 32137 10047
rect 32171 10044 32183 10047
rect 32306 10044 32312 10056
rect 32171 10016 32312 10044
rect 32171 10013 32183 10016
rect 32125 10007 32183 10013
rect 32306 10004 32312 10016
rect 32364 10044 32370 10056
rect 32953 10047 33011 10053
rect 32953 10044 32965 10047
rect 32364 10016 32965 10044
rect 32364 10004 32370 10016
rect 32953 10013 32965 10016
rect 32999 10013 33011 10047
rect 32953 10007 33011 10013
rect 37550 10004 37556 10056
rect 37608 10044 37614 10056
rect 39117 10047 39175 10053
rect 39117 10044 39129 10047
rect 37608 10016 39129 10044
rect 37608 10004 37614 10016
rect 39117 10013 39129 10016
rect 39163 10013 39175 10047
rect 39117 10007 39175 10013
rect 39758 10004 39764 10056
rect 39816 10044 39822 10056
rect 40236 10053 40264 10140
rect 40129 10047 40187 10053
rect 40129 10044 40141 10047
rect 39816 10016 40141 10044
rect 39816 10004 39822 10016
rect 40129 10013 40141 10016
rect 40175 10013 40187 10047
rect 40129 10007 40187 10013
rect 40221 10047 40279 10053
rect 40221 10013 40233 10047
rect 40267 10013 40279 10047
rect 40221 10007 40279 10013
rect 40313 10047 40371 10053
rect 40313 10013 40325 10047
rect 40359 10013 40371 10047
rect 40494 10044 40500 10056
rect 40455 10016 40500 10044
rect 40313 10007 40371 10013
rect 28626 9976 28632 9988
rect 28587 9948 28632 9976
rect 28626 9936 28632 9948
rect 28684 9936 28690 9988
rect 28721 9979 28779 9985
rect 28721 9945 28733 9979
rect 28767 9976 28779 9979
rect 29362 9976 29368 9988
rect 28767 9948 29368 9976
rect 28767 9945 28779 9948
rect 28721 9939 28779 9945
rect 29362 9936 29368 9948
rect 29420 9936 29426 9988
rect 29730 9976 29736 9988
rect 29691 9948 29736 9976
rect 29730 9936 29736 9948
rect 29788 9936 29794 9988
rect 34422 9936 34428 9988
rect 34480 9976 34486 9988
rect 34701 9979 34759 9985
rect 34701 9976 34713 9979
rect 34480 9948 34713 9976
rect 34480 9936 34486 9948
rect 34701 9945 34713 9948
rect 34747 9945 34759 9979
rect 34882 9976 34888 9988
rect 34843 9948 34888 9976
rect 34701 9939 34759 9945
rect 34882 9936 34888 9948
rect 34940 9936 34946 9988
rect 35618 9976 35624 9988
rect 35579 9948 35624 9976
rect 35618 9936 35624 9948
rect 35676 9936 35682 9988
rect 38930 9976 38936 9988
rect 38891 9948 38936 9976
rect 38930 9936 38936 9948
rect 38988 9936 38994 9988
rect 39301 9979 39359 9985
rect 39301 9945 39313 9979
rect 39347 9976 39359 9979
rect 40328 9976 40356 10007
rect 40494 10004 40500 10016
rect 40552 10004 40558 10056
rect 39347 9948 40356 9976
rect 39347 9945 39359 9948
rect 39301 9939 39359 9945
rect 28994 9908 29000 9920
rect 28460 9880 29000 9908
rect 27709 9871 27767 9877
rect 28994 9868 29000 9880
rect 29052 9868 29058 9920
rect 34790 9868 34796 9920
rect 34848 9908 34854 9920
rect 35069 9911 35127 9917
rect 35069 9908 35081 9911
rect 34848 9880 35081 9908
rect 34848 9868 34854 9880
rect 35069 9877 35081 9880
rect 35115 9877 35127 9911
rect 39850 9908 39856 9920
rect 39811 9880 39856 9908
rect 35069 9871 35127 9877
rect 39850 9868 39856 9880
rect 39908 9868 39914 9920
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2682 9704 2688 9716
rect 1452 9676 2688 9704
rect 1452 9664 1458 9676
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 5258 9704 5264 9716
rect 5171 9676 5264 9704
rect 5258 9664 5264 9676
rect 5316 9704 5322 9716
rect 11790 9704 11796 9716
rect 5316 9676 11796 9704
rect 5316 9664 5322 9676
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 13446 9704 13452 9716
rect 13407 9676 13452 9704
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 19337 9707 19395 9713
rect 19337 9673 19349 9707
rect 19383 9704 19395 9707
rect 19426 9704 19432 9716
rect 19383 9676 19432 9704
rect 19383 9673 19395 9676
rect 19337 9667 19395 9673
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 21910 9704 21916 9716
rect 21871 9676 21916 9704
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 30285 9707 30343 9713
rect 30285 9673 30297 9707
rect 30331 9704 30343 9707
rect 32398 9704 32404 9716
rect 30331 9676 32404 9704
rect 30331 9673 30343 9676
rect 30285 9667 30343 9673
rect 1762 9596 1768 9648
rect 1820 9636 1826 9648
rect 2777 9639 2835 9645
rect 1820 9608 2268 9636
rect 1820 9596 1826 9608
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 2096 9540 2145 9568
rect 2096 9528 2102 9540
rect 2133 9537 2145 9540
rect 2179 9537 2191 9571
rect 2240 9568 2268 9608
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 4126 9639 4184 9645
rect 4126 9636 4138 9639
rect 2823 9608 4138 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 4126 9605 4138 9608
rect 4172 9605 4184 9639
rect 4126 9599 4184 9605
rect 7650 9596 7656 9648
rect 7708 9636 7714 9648
rect 8021 9639 8079 9645
rect 8021 9636 8033 9639
rect 7708 9608 8033 9636
rect 7708 9596 7714 9608
rect 8021 9605 8033 9608
rect 8067 9605 8079 9639
rect 8021 9599 8079 9605
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 10321 9639 10379 9645
rect 10321 9636 10333 9639
rect 8812 9608 9260 9636
rect 8812 9596 8818 9608
rect 2296 9571 2354 9577
rect 2296 9568 2308 9571
rect 2240 9540 2308 9568
rect 2133 9531 2191 9537
rect 2296 9537 2308 9540
rect 2342 9537 2354 9571
rect 2296 9531 2354 9537
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 3878 9568 3884 9580
rect 2547 9540 2774 9568
rect 3839 9540 3884 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2424 9500 2452 9531
rect 2590 9500 2596 9512
rect 2424 9472 2596 9500
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 2746 9500 2774 9540
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 9122 9568 9128 9580
rect 3988 9540 9128 9568
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 2746 9472 3341 9500
rect 3329 9469 3341 9472
rect 3375 9500 3387 9503
rect 3988 9500 4016 9540
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9232 9577 9260 9608
rect 9324 9608 10333 9636
rect 9324 9577 9352 9608
rect 10321 9605 10333 9608
rect 10367 9605 10379 9639
rect 10870 9636 10876 9648
rect 10831 9608 10876 9636
rect 10321 9599 10379 9605
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 11698 9636 11704 9648
rect 11659 9608 11704 9636
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 20993 9639 21051 9645
rect 20993 9605 21005 9639
rect 21039 9636 21051 9639
rect 21450 9636 21456 9648
rect 21039 9608 21456 9636
rect 21039 9605 21051 9608
rect 20993 9599 21051 9605
rect 21450 9596 21456 9608
rect 21508 9596 21514 9648
rect 22554 9596 22560 9648
rect 22612 9636 22618 9648
rect 23477 9639 23535 9645
rect 23477 9636 23489 9639
rect 22612 9608 23489 9636
rect 22612 9596 22618 9608
rect 23477 9605 23489 9608
rect 23523 9605 23535 9639
rect 23658 9636 23664 9648
rect 23619 9608 23664 9636
rect 23477 9599 23535 9605
rect 23658 9596 23664 9608
rect 23716 9596 23722 9648
rect 28626 9636 28632 9648
rect 25792 9608 28632 9636
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 9766 9568 9772 9580
rect 9539 9540 9772 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9950 9568 9956 9580
rect 9911 9540 9956 9568
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 11054 9568 11060 9580
rect 10183 9540 11060 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 3375 9472 4016 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 11532 9500 11560 9531
rect 6880 9472 11560 9500
rect 6880 9460 6886 9472
rect 4890 9392 4896 9444
rect 4948 9432 4954 9444
rect 11808 9432 11836 9531
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 11940 9540 11985 9568
rect 11940 9528 11946 9540
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12584 9540 12725 9568
rect 12584 9528 12590 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12894 9568 12900 9580
rect 12855 9540 12900 9568
rect 12713 9531 12771 9537
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 15010 9577 15016 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 13228 9540 13277 9568
rect 13228 9528 13234 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 15004 9568 15016 9577
rect 14971 9540 15016 9568
rect 13265 9531 13323 9537
rect 15004 9531 15016 9540
rect 15010 9528 15016 9531
rect 15068 9528 15074 9580
rect 18322 9528 18328 9580
rect 18380 9577 18386 9580
rect 18380 9568 18392 9577
rect 18380 9540 18425 9568
rect 18380 9531 18392 9540
rect 18380 9528 18386 9531
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 21140 9540 21189 9568
rect 21140 9528 21146 9540
rect 21177 9537 21189 9540
rect 21223 9568 21235 9571
rect 21634 9568 21640 9580
rect 21223 9540 21640 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 21726 9528 21732 9580
rect 21784 9568 21790 9580
rect 21821 9571 21879 9577
rect 21821 9568 21833 9571
rect 21784 9540 21833 9568
rect 21784 9528 21790 9540
rect 21821 9537 21833 9540
rect 21867 9537 21879 9571
rect 22002 9568 22008 9580
rect 21963 9540 22008 9568
rect 21821 9531 21879 9537
rect 22002 9528 22008 9540
rect 22060 9568 22066 9580
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 22060 9540 22477 9568
rect 22060 9528 22066 9540
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9568 23351 9571
rect 23750 9568 23756 9580
rect 23339 9540 23756 9568
rect 23339 9537 23351 9540
rect 23293 9531 23351 9537
rect 23750 9528 23756 9540
rect 23808 9528 23814 9580
rect 25792 9577 25820 9608
rect 28626 9596 28632 9608
rect 28684 9636 28690 9648
rect 29730 9636 29736 9648
rect 28684 9608 29736 9636
rect 28684 9596 28690 9608
rect 29730 9596 29736 9608
rect 29788 9596 29794 9648
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 27617 9571 27675 9577
rect 27617 9537 27629 9571
rect 27663 9537 27675 9571
rect 27798 9568 27804 9580
rect 27759 9540 27804 9568
rect 27617 9531 27675 9537
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12406 9472 13001 9500
rect 12406 9432 12434 9472
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9500 13139 9503
rect 13538 9500 13544 9512
rect 13127 9472 13544 9500
rect 13127 9469 13139 9472
rect 13081 9463 13139 9469
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 14737 9503 14795 9509
rect 14737 9500 14749 9503
rect 14332 9472 14749 9500
rect 14332 9460 14338 9472
rect 14737 9469 14749 9472
rect 14783 9469 14795 9503
rect 18598 9500 18604 9512
rect 18559 9472 18604 9500
rect 14737 9463 14795 9469
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 25498 9500 25504 9512
rect 25459 9472 25504 9500
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 27632 9500 27660 9531
rect 27798 9528 27804 9540
rect 27856 9528 27862 9580
rect 27893 9571 27951 9577
rect 27893 9537 27905 9571
rect 27939 9537 27951 9571
rect 27893 9531 27951 9537
rect 27706 9500 27712 9512
rect 27632 9472 27712 9500
rect 27706 9460 27712 9472
rect 27764 9460 27770 9512
rect 27908 9500 27936 9531
rect 27982 9528 27988 9580
rect 28040 9568 28046 9580
rect 32140 9577 32168 9676
rect 32398 9664 32404 9676
rect 32456 9664 32462 9716
rect 32674 9664 32680 9716
rect 32732 9704 32738 9716
rect 37550 9704 37556 9716
rect 32732 9676 37556 9704
rect 32732 9664 32738 9676
rect 37550 9664 37556 9676
rect 37608 9664 37614 9716
rect 39758 9704 39764 9716
rect 39719 9676 39764 9704
rect 39758 9664 39764 9676
rect 39816 9664 39822 9716
rect 34790 9636 34796 9648
rect 34440 9608 34796 9636
rect 28721 9571 28779 9577
rect 28721 9568 28733 9571
rect 28040 9540 28733 9568
rect 28040 9528 28046 9540
rect 28721 9537 28733 9540
rect 28767 9537 28779 9571
rect 28721 9531 28779 9537
rect 32125 9571 32183 9577
rect 32125 9537 32137 9571
rect 32171 9537 32183 9571
rect 32125 9531 32183 9537
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9568 32367 9571
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 32355 9540 33057 9568
rect 32355 9537 32367 9540
rect 32309 9531 32367 9537
rect 33045 9537 33057 9540
rect 33091 9568 33103 9571
rect 33318 9568 33324 9580
rect 33091 9540 33324 9568
rect 33091 9537 33103 9540
rect 33045 9531 33103 9537
rect 28074 9500 28080 9512
rect 27908 9472 28080 9500
rect 28074 9460 28080 9472
rect 28132 9460 28138 9512
rect 27246 9432 27252 9444
rect 4948 9404 11836 9432
rect 11900 9404 12434 9432
rect 15672 9404 17356 9432
rect 4948 9392 4954 9404
rect 8846 9364 8852 9376
rect 8807 9336 8852 9364
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9950 9364 9956 9376
rect 9732 9336 9956 9364
rect 9732 9324 9738 9336
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 11900 9364 11928 9404
rect 10100 9336 11928 9364
rect 12069 9367 12127 9373
rect 10100 9324 10106 9336
rect 12069 9333 12081 9367
rect 12115 9364 12127 9367
rect 15672 9364 15700 9404
rect 16114 9364 16120 9376
rect 12115 9336 15700 9364
rect 16075 9336 16120 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17218 9364 17224 9376
rect 16908 9336 17224 9364
rect 16908 9324 16914 9336
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17328 9364 17356 9404
rect 18616 9404 27252 9432
rect 18616 9364 18644 9404
rect 27246 9392 27252 9404
rect 27304 9392 27310 9444
rect 17328 9336 18644 9364
rect 19886 9324 19892 9376
rect 19944 9364 19950 9376
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19944 9336 19993 9364
rect 19944 9324 19950 9336
rect 19981 9333 19993 9336
rect 20027 9333 20039 9367
rect 19981 9327 20039 9333
rect 20346 9324 20352 9376
rect 20404 9364 20410 9376
rect 20809 9367 20867 9373
rect 20809 9364 20821 9367
rect 20404 9336 20821 9364
rect 20404 9324 20410 9336
rect 20809 9333 20821 9336
rect 20855 9333 20867 9367
rect 28258 9364 28264 9376
rect 28219 9336 28264 9364
rect 20809 9327 20867 9333
rect 28258 9324 28264 9336
rect 28316 9324 28322 9376
rect 28736 9364 28764 9531
rect 33318 9528 33324 9540
rect 33376 9528 33382 9580
rect 34054 9528 34060 9580
rect 34112 9568 34118 9580
rect 34440 9577 34468 9608
rect 34790 9596 34796 9608
rect 34848 9596 34854 9648
rect 34885 9639 34943 9645
rect 34885 9605 34897 9639
rect 34931 9636 34943 9639
rect 36458 9639 36516 9645
rect 36458 9636 36470 9639
rect 34931 9608 36470 9636
rect 34931 9605 34943 9608
rect 34885 9599 34943 9605
rect 36458 9605 36470 9608
rect 36504 9605 36516 9639
rect 36458 9599 36516 9605
rect 38688 9639 38746 9645
rect 38688 9605 38700 9639
rect 38734 9636 38746 9639
rect 39850 9636 39856 9648
rect 38734 9608 39856 9636
rect 38734 9605 38746 9608
rect 38688 9599 38746 9605
rect 39850 9596 39856 9608
rect 39908 9596 39914 9648
rect 34241 9571 34299 9577
rect 34241 9568 34253 9571
rect 34112 9540 34253 9568
rect 34112 9528 34118 9540
rect 34241 9537 34253 9540
rect 34287 9537 34299 9571
rect 34241 9531 34299 9537
rect 34425 9571 34483 9577
rect 34425 9537 34437 9571
rect 34471 9537 34483 9571
rect 34425 9531 34483 9537
rect 34517 9571 34575 9577
rect 34517 9537 34529 9571
rect 34563 9537 34575 9571
rect 34517 9531 34575 9537
rect 34609 9571 34667 9577
rect 34609 9537 34621 9571
rect 34655 9568 34667 9571
rect 34698 9568 34704 9580
rect 34655 9540 34704 9568
rect 34655 9537 34667 9540
rect 34609 9531 34667 9537
rect 31294 9500 31300 9512
rect 31255 9472 31300 9500
rect 31294 9460 31300 9472
rect 31352 9460 31358 9512
rect 31573 9503 31631 9509
rect 31573 9469 31585 9503
rect 31619 9500 31631 9503
rect 32582 9500 32588 9512
rect 31619 9472 32588 9500
rect 31619 9469 31631 9472
rect 31573 9463 31631 9469
rect 32582 9460 32588 9472
rect 32640 9500 32646 9512
rect 32769 9503 32827 9509
rect 32769 9500 32781 9503
rect 32640 9472 32781 9500
rect 32640 9460 32646 9472
rect 32769 9469 32781 9472
rect 32815 9469 32827 9503
rect 32769 9463 32827 9469
rect 34532 9500 34560 9531
rect 34698 9528 34704 9540
rect 34756 9528 34762 9580
rect 38838 9528 38844 9580
rect 38896 9568 38902 9580
rect 38933 9571 38991 9577
rect 38933 9568 38945 9571
rect 38896 9540 38945 9568
rect 38896 9528 38902 9540
rect 38933 9537 38945 9540
rect 38979 9537 38991 9571
rect 38933 9531 38991 9537
rect 35618 9500 35624 9512
rect 34532 9472 35624 9500
rect 32217 9435 32275 9441
rect 32217 9401 32229 9435
rect 32263 9432 32275 9435
rect 34532 9432 34560 9472
rect 35618 9460 35624 9472
rect 35676 9460 35682 9512
rect 36722 9500 36728 9512
rect 36683 9472 36728 9500
rect 36722 9460 36728 9472
rect 36780 9460 36786 9512
rect 32263 9404 34560 9432
rect 34716 9404 35857 9432
rect 32263 9401 32275 9404
rect 32217 9395 32275 9401
rect 34716 9364 34744 9404
rect 28736 9336 34744 9364
rect 34790 9324 34796 9376
rect 34848 9364 34854 9376
rect 35345 9367 35403 9373
rect 35345 9364 35357 9367
rect 34848 9336 35357 9364
rect 34848 9324 34854 9336
rect 35345 9333 35357 9336
rect 35391 9333 35403 9367
rect 35829 9364 35857 9404
rect 36354 9364 36360 9376
rect 35829 9336 36360 9364
rect 35345 9327 35403 9333
rect 36354 9324 36360 9336
rect 36412 9324 36418 9376
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 11054 9160 11060 9172
rect 10367 9132 11060 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 15286 9160 15292 9172
rect 13780 9132 15292 9160
rect 13780 9120 13786 9132
rect 15286 9120 15292 9132
rect 15344 9160 15350 9172
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 15344 9132 16313 9160
rect 15344 9120 15350 9132
rect 16301 9129 16313 9132
rect 16347 9129 16359 9163
rect 16301 9123 16359 9129
rect 24397 9163 24455 9169
rect 24397 9129 24409 9163
rect 24443 9160 24455 9163
rect 24854 9160 24860 9172
rect 24443 9132 24860 9160
rect 24443 9129 24455 9132
rect 24397 9123 24455 9129
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 26145 9163 26203 9169
rect 26145 9129 26157 9163
rect 26191 9160 26203 9163
rect 27338 9160 27344 9172
rect 26191 9132 27344 9160
rect 26191 9129 26203 9132
rect 26145 9123 26203 9129
rect 27338 9120 27344 9132
rect 27396 9120 27402 9172
rect 27798 9120 27804 9172
rect 27856 9160 27862 9172
rect 27893 9163 27951 9169
rect 27893 9160 27905 9163
rect 27856 9132 27905 9160
rect 27856 9120 27862 9132
rect 27893 9129 27905 9132
rect 27939 9129 27951 9163
rect 27893 9123 27951 9129
rect 28350 9120 28356 9172
rect 28408 9160 28414 9172
rect 31389 9163 31447 9169
rect 31389 9160 31401 9163
rect 28408 9132 31401 9160
rect 28408 9120 28414 9132
rect 31389 9129 31401 9132
rect 31435 9129 31447 9163
rect 31389 9123 31447 9129
rect 33686 9120 33692 9172
rect 33744 9160 33750 9172
rect 34698 9160 34704 9172
rect 33744 9132 34704 9160
rect 33744 9120 33750 9132
rect 34698 9120 34704 9132
rect 34756 9120 34762 9172
rect 14366 9052 14372 9104
rect 14424 9092 14430 9104
rect 16853 9095 16911 9101
rect 16853 9092 16865 9095
rect 14424 9064 16865 9092
rect 14424 9052 14430 9064
rect 16853 9061 16865 9064
rect 16899 9061 16911 9095
rect 16853 9055 16911 9061
rect 21358 9052 21364 9104
rect 21416 9092 21422 9104
rect 25498 9092 25504 9104
rect 21416 9064 25504 9092
rect 21416 9052 21422 9064
rect 2038 8984 2044 9036
rect 2096 9024 2102 9036
rect 2317 9027 2375 9033
rect 2317 9024 2329 9027
rect 2096 8996 2329 9024
rect 2096 8984 2102 8996
rect 2317 8993 2329 8996
rect 2363 8993 2375 9027
rect 2317 8987 2375 8993
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 9024 2651 9027
rect 2958 9024 2964 9036
rect 2639 8996 2964 9024
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 2958 8984 2964 8996
rect 3016 9024 3022 9036
rect 3234 9024 3240 9036
rect 3016 8996 3240 9024
rect 3016 8984 3022 8996
rect 3234 8984 3240 8996
rect 3292 8984 3298 9036
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 4028 8996 5457 9024
rect 4028 8984 4034 8996
rect 5445 8993 5457 8996
rect 5491 9024 5503 9027
rect 8754 9024 8760 9036
rect 5491 8996 5580 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 5552 8968 5580 8996
rect 7668 8996 8760 9024
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 2740 8928 3801 8956
rect 2740 8916 2746 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 3936 8928 5028 8956
rect 3936 8916 3942 8928
rect 3973 8891 4031 8897
rect 3973 8857 3985 8891
rect 4019 8888 4031 8891
rect 4890 8888 4896 8900
rect 4019 8860 4896 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 5000 8888 5028 8928
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 7668 8965 7696 8996
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 8938 9024 8944 9036
rect 8899 8996 8944 9024
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 15381 9027 15439 9033
rect 15381 9024 15393 9027
rect 15252 8996 15393 9024
rect 15252 8984 15258 8996
rect 15381 8993 15393 8996
rect 15427 8993 15439 9027
rect 15381 8987 15439 8993
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 16390 9024 16396 9036
rect 15528 8996 16396 9024
rect 15528 8984 15534 8996
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 20898 9024 20904 9036
rect 19444 8996 19656 9024
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 5644 8928 7573 8956
rect 5644 8888 5672 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 5000 8860 5672 8888
rect 5712 8891 5770 8897
rect 5712 8857 5724 8891
rect 5758 8888 5770 8891
rect 7285 8891 7343 8897
rect 7285 8888 7297 8891
rect 5758 8860 7297 8888
rect 5758 8857 5770 8860
rect 5712 8851 5770 8857
rect 7285 8857 7297 8860
rect 7331 8857 7343 8891
rect 7576 8888 7604 8919
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 7929 8959 7987 8965
rect 7800 8928 7845 8956
rect 7800 8916 7806 8928
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 7944 8888 7972 8919
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 9197 8959 9255 8965
rect 9197 8956 9209 8959
rect 8904 8928 9209 8956
rect 8904 8916 8910 8928
rect 9197 8925 9209 8928
rect 9243 8925 9255 8959
rect 9197 8919 9255 8925
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 15105 8959 15163 8965
rect 15105 8956 15117 8959
rect 14516 8928 15117 8956
rect 14516 8916 14522 8928
rect 15105 8925 15117 8928
rect 15151 8925 15163 8959
rect 15105 8919 15163 8925
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15657 8959 15715 8965
rect 15657 8925 15669 8959
rect 15703 8956 15715 8959
rect 17310 8956 17316 8968
rect 15703 8928 17316 8956
rect 15703 8925 15715 8928
rect 15657 8919 15715 8925
rect 9766 8888 9772 8900
rect 7576 8860 7696 8888
rect 7944 8860 9772 8888
rect 7285 8851 7343 8857
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 3234 8820 3240 8832
rect 3191 8792 3240 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 3384 8792 4169 8820
rect 3384 8780 3390 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 7668 8820 7696 8860
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 11238 8848 11244 8900
rect 11296 8888 11302 8900
rect 12161 8891 12219 8897
rect 12161 8888 12173 8891
rect 11296 8860 12173 8888
rect 11296 8848 11302 8860
rect 12161 8857 12173 8860
rect 12207 8857 12219 8891
rect 15304 8888 15332 8919
rect 17310 8916 17316 8928
rect 17368 8916 17374 8968
rect 19444 8965 19472 8996
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 18616 8928 19441 8956
rect 16298 8888 16304 8900
rect 12161 8851 12219 8857
rect 12406 8860 14688 8888
rect 15304 8860 16304 8888
rect 8202 8820 8208 8832
rect 7668 8792 8208 8820
rect 4157 8783 4215 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 10870 8820 10876 8832
rect 9180 8792 10876 8820
rect 9180 8780 9186 8792
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11701 8823 11759 8829
rect 11701 8789 11713 8823
rect 11747 8820 11759 8823
rect 11882 8820 11888 8832
rect 11747 8792 11888 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 11882 8780 11888 8792
rect 11940 8820 11946 8832
rect 12406 8820 12434 8860
rect 14660 8832 14688 8860
rect 16298 8848 16304 8860
rect 16356 8848 16362 8900
rect 11940 8792 12434 8820
rect 12805 8823 12863 8829
rect 11940 8780 11946 8792
rect 12805 8789 12817 8823
rect 12851 8820 12863 8823
rect 12986 8820 12992 8832
rect 12851 8792 12992 8820
rect 12851 8789 12863 8792
rect 12805 8783 12863 8789
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13446 8820 13452 8832
rect 13407 8792 13452 8820
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 14642 8820 14648 8832
rect 14603 8792 14648 8820
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15378 8820 15384 8832
rect 15068 8792 15384 8820
rect 15068 8780 15074 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15838 8820 15844 8832
rect 15799 8792 15844 8820
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 18616 8829 18644 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19521 8959 19579 8965
rect 19521 8925 19533 8959
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 18966 8848 18972 8900
rect 19024 8888 19030 8900
rect 19536 8888 19564 8919
rect 19024 8860 19564 8888
rect 19024 8848 19030 8860
rect 18601 8823 18659 8829
rect 18601 8820 18613 8823
rect 16080 8792 18613 8820
rect 16080 8780 16086 8792
rect 18601 8789 18613 8792
rect 18647 8789 18659 8823
rect 19628 8820 19656 8996
rect 20456 8996 20904 9024
rect 20162 8956 20168 8968
rect 20123 8928 20168 8956
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 20346 8956 20352 8968
rect 20307 8928 20352 8956
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 20456 8965 20484 8996
rect 20898 8984 20904 8996
rect 20956 8984 20962 9036
rect 22830 9024 22836 9036
rect 21008 8996 22836 9024
rect 20441 8959 20499 8965
rect 20441 8925 20453 8959
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 20530 8916 20536 8968
rect 20588 8956 20594 8968
rect 21008 8956 21036 8996
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 20588 8928 21036 8956
rect 20588 8916 20594 8928
rect 21910 8916 21916 8968
rect 21968 8956 21974 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 21968 8928 24593 8956
rect 21968 8916 21974 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 19705 8891 19763 8897
rect 19705 8857 19717 8891
rect 19751 8888 19763 8891
rect 24486 8888 24492 8900
rect 19751 8860 24492 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 24486 8848 24492 8860
rect 24544 8848 24550 8900
rect 20346 8820 20352 8832
rect 19628 8792 20352 8820
rect 18601 8783 18659 8789
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 20806 8820 20812 8832
rect 20767 8792 20812 8820
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 24596 8820 24624 8919
rect 24670 8916 24676 8968
rect 24728 8956 24734 8968
rect 24946 8956 24952 8968
rect 24728 8928 24773 8956
rect 24907 8928 24952 8956
rect 24728 8916 24734 8928
rect 24946 8916 24952 8928
rect 25004 8916 25010 8968
rect 24765 8891 24823 8897
rect 24765 8857 24777 8891
rect 24811 8888 24823 8891
rect 25319 8888 25347 9064
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 26602 9092 26608 9104
rect 25608 9064 26608 9092
rect 25608 8965 25636 9064
rect 26602 9052 26608 9064
rect 26660 9052 26666 9104
rect 27522 9052 27528 9104
rect 27580 9092 27586 9104
rect 29546 9092 29552 9104
rect 27580 9064 29552 9092
rect 27580 9052 27586 9064
rect 29546 9052 29552 9064
rect 29604 9052 29610 9104
rect 33505 9095 33563 9101
rect 33505 9061 33517 9095
rect 33551 9092 33563 9095
rect 33551 9064 35020 9092
rect 33551 9061 33563 9064
rect 33505 9055 33563 9061
rect 27614 8984 27620 9036
rect 27672 9024 27678 9036
rect 27798 9024 27804 9036
rect 27672 8996 27804 9024
rect 27672 8984 27678 8996
rect 27798 8984 27804 8996
rect 27856 8984 27862 9036
rect 28258 8984 28264 9036
rect 28316 9024 28322 9036
rect 28316 8996 29684 9024
rect 28316 8984 28322 8996
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8925 25651 8959
rect 25593 8919 25651 8925
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8925 25835 8959
rect 25777 8919 25835 8925
rect 25961 8959 26019 8965
rect 25961 8925 25973 8959
rect 26007 8956 26019 8959
rect 26234 8956 26240 8968
rect 26007 8928 26240 8956
rect 26007 8925 26019 8928
rect 25961 8919 26019 8925
rect 25792 8888 25820 8919
rect 26234 8916 26240 8928
rect 26292 8916 26298 8968
rect 29546 8956 29552 8968
rect 29507 8928 29552 8956
rect 29546 8916 29552 8928
rect 29604 8916 29610 8968
rect 29656 8956 29684 8996
rect 31294 8984 31300 9036
rect 31352 9024 31358 9036
rect 34790 9024 34796 9036
rect 31352 8996 31800 9024
rect 31352 8984 31358 8996
rect 29805 8959 29863 8965
rect 29805 8956 29817 8959
rect 29656 8928 29817 8956
rect 29805 8925 29817 8928
rect 29851 8925 29863 8959
rect 31570 8956 31576 8968
rect 31531 8928 31576 8956
rect 29805 8919 29863 8925
rect 31570 8916 31576 8928
rect 31628 8916 31634 8968
rect 31772 8965 31800 8996
rect 33060 8996 34796 9024
rect 31757 8959 31815 8965
rect 31757 8925 31769 8959
rect 31803 8925 31815 8959
rect 31938 8956 31944 8968
rect 31899 8928 31944 8956
rect 31757 8919 31815 8925
rect 31938 8916 31944 8928
rect 31996 8916 32002 8968
rect 32306 8916 32312 8968
rect 32364 8956 32370 8968
rect 33060 8965 33088 8996
rect 34790 8984 34796 8996
rect 34848 8984 34854 9036
rect 32677 8959 32735 8965
rect 32677 8956 32689 8959
rect 32364 8928 32689 8956
rect 32364 8916 32370 8928
rect 32677 8925 32689 8928
rect 32723 8925 32735 8959
rect 32677 8919 32735 8925
rect 33045 8959 33103 8965
rect 33045 8925 33057 8959
rect 33091 8925 33103 8959
rect 33045 8919 33103 8925
rect 33686 8916 33692 8968
rect 33744 8956 33750 8968
rect 33781 8959 33839 8965
rect 33781 8956 33793 8959
rect 33744 8928 33793 8956
rect 33744 8916 33750 8928
rect 33781 8925 33793 8928
rect 33827 8925 33839 8959
rect 33781 8919 33839 8925
rect 33873 8959 33931 8965
rect 33873 8925 33885 8959
rect 33919 8925 33931 8959
rect 33873 8919 33931 8925
rect 24811 8860 25820 8888
rect 25869 8891 25927 8897
rect 24811 8857 24823 8860
rect 24765 8851 24823 8857
rect 25869 8857 25881 8891
rect 25915 8857 25927 8891
rect 25869 8851 25927 8857
rect 25682 8820 25688 8832
rect 24596 8792 25688 8820
rect 25682 8780 25688 8792
rect 25740 8780 25746 8832
rect 25884 8820 25912 8851
rect 27246 8848 27252 8900
rect 27304 8888 27310 8900
rect 27525 8891 27583 8897
rect 27525 8888 27537 8891
rect 27304 8860 27537 8888
rect 27304 8848 27310 8860
rect 27525 8857 27537 8860
rect 27571 8857 27583 8891
rect 27525 8851 27583 8857
rect 27709 8891 27767 8897
rect 27709 8857 27721 8891
rect 27755 8857 27767 8891
rect 27709 8851 27767 8857
rect 27614 8820 27620 8832
rect 25884 8792 27620 8820
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 27724 8820 27752 8851
rect 31478 8848 31484 8900
rect 31536 8888 31542 8900
rect 31665 8891 31723 8897
rect 31665 8888 31677 8891
rect 31536 8860 31677 8888
rect 31536 8848 31542 8860
rect 31665 8857 31677 8860
rect 31711 8857 31723 8891
rect 32766 8888 32772 8900
rect 32727 8860 32772 8888
rect 31665 8851 31723 8857
rect 32766 8848 32772 8860
rect 32824 8848 32830 8900
rect 32861 8891 32919 8897
rect 32861 8857 32873 8891
rect 32907 8857 32919 8891
rect 32861 8851 32919 8857
rect 29822 8820 29828 8832
rect 27724 8792 29828 8820
rect 29822 8780 29828 8792
rect 29880 8820 29886 8832
rect 30929 8823 30987 8829
rect 30929 8820 30941 8823
rect 29880 8792 30941 8820
rect 29880 8780 29886 8792
rect 30929 8789 30941 8792
rect 30975 8789 30987 8823
rect 32490 8820 32496 8832
rect 32451 8792 32496 8820
rect 30929 8783 30987 8789
rect 32490 8780 32496 8792
rect 32548 8780 32554 8832
rect 32582 8780 32588 8832
rect 32640 8820 32646 8832
rect 32876 8820 32904 8851
rect 32640 8792 32904 8820
rect 33888 8820 33916 8919
rect 33962 8916 33968 8968
rect 34020 8956 34026 8968
rect 34149 8959 34207 8965
rect 34020 8928 34065 8956
rect 34020 8916 34026 8928
rect 34149 8925 34161 8959
rect 34195 8956 34207 8959
rect 34238 8956 34244 8968
rect 34195 8928 34244 8956
rect 34195 8925 34207 8928
rect 34149 8919 34207 8925
rect 34238 8916 34244 8928
rect 34296 8916 34302 8968
rect 34992 8888 35020 9064
rect 36633 9027 36691 9033
rect 36633 8993 36645 9027
rect 36679 9024 36691 9027
rect 36722 9024 36728 9036
rect 36679 8996 36728 9024
rect 36679 8993 36691 8996
rect 36633 8987 36691 8993
rect 36722 8984 36728 8996
rect 36780 8984 36786 9036
rect 68094 8956 68100 8968
rect 68055 8928 68100 8956
rect 68094 8916 68100 8928
rect 68152 8916 68158 8968
rect 36366 8891 36424 8897
rect 36366 8888 36378 8891
rect 34992 8860 36378 8888
rect 36366 8857 36378 8860
rect 36412 8857 36424 8891
rect 36366 8851 36424 8857
rect 34606 8820 34612 8832
rect 33888 8792 34612 8820
rect 32640 8780 32646 8792
rect 34606 8780 34612 8792
rect 34664 8780 34670 8832
rect 35250 8820 35256 8832
rect 35211 8792 35256 8820
rect 35250 8780 35256 8792
rect 35308 8780 35314 8832
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 4801 8619 4859 8625
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 4890 8616 4896 8628
rect 4847 8588 4896 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 7561 8619 7619 8625
rect 7561 8585 7573 8619
rect 7607 8616 7619 8619
rect 7742 8616 7748 8628
rect 7607 8588 7748 8616
rect 7607 8585 7619 8588
rect 7561 8579 7619 8585
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8113 8619 8171 8625
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8202 8616 8208 8628
rect 8159 8588 8208 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 9968 8588 11284 8616
rect 3326 8548 3332 8560
rect 2516 8520 3332 8548
rect 2038 8440 2044 8492
rect 2096 8480 2102 8492
rect 2516 8489 2544 8520
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 3970 8548 3976 8560
rect 3436 8520 3976 8548
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 2096 8452 2329 8480
rect 2096 8440 2102 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 3142 8480 3148 8492
rect 2731 8452 3148 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2608 8356 2636 8443
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3436 8489 3464 8520
rect 3970 8508 3976 8520
rect 4028 8508 4034 8560
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 7377 8551 7435 8557
rect 7377 8548 7389 8551
rect 6880 8520 7389 8548
rect 6880 8508 6886 8520
rect 7377 8517 7389 8520
rect 7423 8517 7435 8551
rect 7377 8511 7435 8517
rect 7926 8508 7932 8560
rect 7984 8548 7990 8560
rect 9582 8548 9588 8560
rect 7984 8520 9588 8548
rect 7984 8508 7990 8520
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8449 3479 8483
rect 3677 8483 3735 8489
rect 3677 8480 3689 8483
rect 3421 8443 3479 8449
rect 3528 8452 3689 8480
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 3528 8412 3556 8452
rect 3677 8449 3689 8452
rect 3723 8449 3735 8483
rect 3677 8443 3735 8449
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 7064 8452 7205 8480
rect 7064 8440 7070 8452
rect 7193 8449 7205 8452
rect 7239 8480 7251 8483
rect 9674 8480 9680 8492
rect 7239 8452 9680 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 9968 8412 9996 8588
rect 10134 8508 10140 8560
rect 10192 8548 10198 8560
rect 10192 8520 11008 8548
rect 10192 8508 10198 8520
rect 10980 8489 11008 8520
rect 10709 8483 10767 8489
rect 10709 8449 10721 8483
rect 10755 8480 10767 8483
rect 10965 8483 11023 8489
rect 10755 8452 10916 8480
rect 10755 8449 10767 8452
rect 10709 8443 10767 8449
rect 3007 8384 3556 8412
rect 9600 8384 9996 8412
rect 10888 8412 10916 8452
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 11256 8480 11284 8588
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 14090 8616 14096 8628
rect 12584 8588 14096 8616
rect 12584 8576 12590 8588
rect 14090 8576 14096 8588
rect 14148 8616 14154 8628
rect 14148 8588 14596 8616
rect 14148 8576 14154 8588
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11256 8452 11713 8480
rect 10965 8443 11023 8449
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11701 8443 11759 8449
rect 11808 8452 12081 8480
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 10888 8384 11529 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 2590 8304 2596 8356
rect 2648 8304 2654 8356
rect 5813 8347 5871 8353
rect 5813 8313 5825 8347
rect 5859 8344 5871 8347
rect 5902 8344 5908 8356
rect 5859 8316 5908 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 6178 8304 6184 8356
rect 6236 8344 6242 8356
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 6236 8316 6653 8344
rect 6236 8304 6242 8316
rect 6641 8313 6653 8316
rect 6687 8313 6699 8347
rect 9030 8344 9036 8356
rect 8991 8316 9036 8344
rect 6641 8307 6699 8313
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 9214 8304 9220 8356
rect 9272 8344 9278 8356
rect 9600 8353 9628 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 9585 8347 9643 8353
rect 9585 8344 9597 8347
rect 9272 8316 9597 8344
rect 9272 8304 9278 8316
rect 9585 8313 9597 8316
rect 9631 8313 9643 8347
rect 9585 8307 9643 8313
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11808 8344 11836 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12250 8480 12256 8492
rect 12211 8452 12256 8480
rect 12069 8443 12127 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 13998 8480 14004 8492
rect 14056 8489 14062 8492
rect 13968 8452 14004 8480
rect 13998 8440 14004 8452
rect 14056 8443 14068 8489
rect 14568 8480 14596 8588
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 20254 8616 20260 8628
rect 14976 8588 20260 8616
rect 14976 8576 14982 8588
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 21450 8576 21456 8628
rect 21508 8616 21514 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 21508 8588 21833 8616
rect 21508 8576 21514 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 25685 8619 25743 8625
rect 25685 8585 25697 8619
rect 25731 8616 25743 8619
rect 25774 8616 25780 8628
rect 25731 8588 25780 8616
rect 25731 8585 25743 8588
rect 25685 8579 25743 8585
rect 25774 8576 25780 8588
rect 25832 8576 25838 8628
rect 29362 8616 29368 8628
rect 27448 8588 29368 8616
rect 15838 8508 15844 8560
rect 15896 8548 15902 8560
rect 18794 8551 18852 8557
rect 18794 8548 18806 8551
rect 15896 8520 18806 8548
rect 15896 8508 15902 8520
rect 18794 8517 18806 8520
rect 18840 8517 18852 8551
rect 18794 8511 18852 8517
rect 20806 8508 20812 8560
rect 20864 8548 20870 8560
rect 22934 8551 22992 8557
rect 22934 8548 22946 8551
rect 20864 8520 22946 8548
rect 20864 8508 20870 8520
rect 22934 8517 22946 8520
rect 22980 8517 22992 8551
rect 22934 8511 22992 8517
rect 23842 8508 23848 8560
rect 23900 8548 23906 8560
rect 24397 8551 24455 8557
rect 24397 8548 24409 8551
rect 23900 8520 24409 8548
rect 23900 8508 23906 8520
rect 24397 8517 24409 8520
rect 24443 8548 24455 8551
rect 24670 8548 24676 8560
rect 24443 8520 24676 8548
rect 24443 8517 24455 8520
rect 24397 8511 24455 8517
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 25961 8551 26019 8557
rect 25961 8517 25973 8551
rect 26007 8548 26019 8551
rect 26418 8548 26424 8560
rect 26007 8520 26424 8548
rect 26007 8517 26019 8520
rect 25961 8511 26019 8517
rect 26418 8508 26424 8520
rect 26476 8508 26482 8560
rect 27448 8557 27476 8588
rect 29362 8576 29368 8588
rect 29420 8576 29426 8628
rect 29638 8576 29644 8628
rect 29696 8616 29702 8628
rect 32125 8619 32183 8625
rect 32125 8616 32137 8619
rect 29696 8588 32137 8616
rect 29696 8576 29702 8588
rect 32125 8585 32137 8588
rect 32171 8585 32183 8619
rect 33962 8616 33968 8628
rect 33923 8588 33968 8616
rect 32125 8579 32183 8585
rect 33962 8576 33968 8588
rect 34020 8576 34026 8628
rect 34330 8576 34336 8628
rect 34388 8616 34394 8628
rect 37369 8619 37427 8625
rect 37369 8616 37381 8619
rect 34388 8588 37381 8616
rect 34388 8576 34394 8588
rect 27433 8551 27491 8557
rect 27433 8517 27445 8551
rect 27479 8517 27491 8551
rect 27433 8511 27491 8517
rect 27617 8551 27675 8557
rect 27617 8517 27629 8551
rect 27663 8548 27675 8551
rect 28721 8551 28779 8557
rect 27663 8520 28304 8548
rect 27663 8517 27675 8520
rect 27617 8511 27675 8517
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14568 8452 15117 8480
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 19150 8480 19156 8492
rect 15105 8443 15163 8449
rect 16868 8452 19156 8480
rect 14056 8440 14062 8443
rect 11885 8415 11943 8421
rect 11885 8381 11897 8415
rect 11931 8381 11943 8415
rect 11885 8375 11943 8381
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8412 12035 8415
rect 12618 8412 12624 8424
rect 12023 8384 12624 8412
rect 12023 8381 12035 8384
rect 11977 8375 12035 8381
rect 11020 8316 11836 8344
rect 11020 8304 11026 8316
rect 10594 8236 10600 8288
rect 10652 8276 10658 8288
rect 11054 8276 11060 8288
rect 10652 8248 11060 8276
rect 10652 8236 10658 8248
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11900 8276 11928 8375
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 14274 8412 14280 8424
rect 14235 8384 14280 8412
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14700 8384 14841 8412
rect 14700 8372 14706 8384
rect 14829 8381 14841 8384
rect 14875 8412 14887 8415
rect 16868 8412 16896 8452
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 20441 8483 20499 8489
rect 20441 8449 20453 8483
rect 20487 8480 20499 8483
rect 21358 8480 21364 8492
rect 20487 8452 21364 8480
rect 20487 8449 20499 8452
rect 20441 8443 20499 8449
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8480 23259 8483
rect 23934 8480 23940 8492
rect 23247 8452 23940 8480
rect 23247 8449 23259 8452
rect 23201 8443 23259 8449
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 24210 8480 24216 8492
rect 24171 8452 24216 8480
rect 24210 8440 24216 8452
rect 24268 8480 24274 8492
rect 24762 8480 24768 8492
rect 24268 8452 24768 8480
rect 24268 8440 24274 8452
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 25682 8440 25688 8492
rect 25740 8480 25746 8492
rect 25869 8483 25927 8489
rect 25869 8480 25881 8483
rect 25740 8452 25881 8480
rect 25740 8440 25746 8452
rect 25869 8449 25881 8452
rect 25915 8449 25927 8483
rect 25869 8443 25927 8449
rect 26053 8483 26111 8489
rect 26053 8449 26065 8483
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 26237 8483 26295 8489
rect 26237 8449 26249 8483
rect 26283 8480 26295 8483
rect 26510 8480 26516 8492
rect 26283 8452 26516 8480
rect 26283 8449 26295 8452
rect 26237 8443 26295 8449
rect 14875 8384 16896 8412
rect 19061 8415 19119 8421
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 19061 8381 19073 8415
rect 19107 8381 19119 8415
rect 20162 8412 20168 8424
rect 20123 8384 20168 8412
rect 19061 8375 19119 8381
rect 16850 8344 16856 8356
rect 14292 8316 16856 8344
rect 11204 8248 11928 8276
rect 12897 8279 12955 8285
rect 11204 8236 11210 8248
rect 12897 8245 12909 8279
rect 12943 8276 12955 8279
rect 13078 8276 13084 8288
rect 12943 8248 13084 8276
rect 12943 8245 12955 8248
rect 12897 8239 12955 8245
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 14292 8276 14320 8316
rect 16850 8304 16856 8316
rect 16908 8304 16914 8356
rect 16942 8304 16948 8356
rect 17000 8344 17006 8356
rect 17037 8347 17095 8353
rect 17037 8344 17049 8347
rect 17000 8316 17049 8344
rect 17000 8304 17006 8316
rect 17037 8313 17049 8316
rect 17083 8313 17095 8347
rect 17037 8307 17095 8313
rect 17310 8304 17316 8356
rect 17368 8344 17374 8356
rect 17681 8347 17739 8353
rect 17681 8344 17693 8347
rect 17368 8316 17693 8344
rect 17368 8304 17374 8316
rect 17681 8313 17693 8316
rect 17727 8313 17739 8347
rect 17681 8307 17739 8313
rect 13688 8248 14320 8276
rect 13688 8236 13694 8248
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 19076 8276 19104 8375
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 24581 8415 24639 8421
rect 24581 8381 24593 8415
rect 24627 8412 24639 8415
rect 25130 8412 25136 8424
rect 24627 8384 25136 8412
rect 24627 8381 24639 8384
rect 24581 8375 24639 8381
rect 25130 8372 25136 8384
rect 25188 8372 25194 8424
rect 25498 8372 25504 8424
rect 25556 8412 25562 8424
rect 26068 8412 26096 8443
rect 26510 8440 26516 8452
rect 26568 8440 26574 8492
rect 27246 8480 27252 8492
rect 27207 8452 27252 8480
rect 27246 8440 27252 8452
rect 27304 8440 27310 8492
rect 27706 8440 27712 8492
rect 27764 8480 27770 8492
rect 28276 8489 28304 8520
rect 28721 8517 28733 8551
rect 28767 8548 28779 8551
rect 30478 8551 30536 8557
rect 30478 8548 30490 8551
rect 28767 8520 30490 8548
rect 28767 8517 28779 8520
rect 28721 8511 28779 8517
rect 30478 8517 30490 8520
rect 30524 8517 30536 8551
rect 30478 8511 30536 8517
rect 31570 8508 31576 8560
rect 31628 8548 31634 8560
rect 31628 8520 32720 8548
rect 31628 8508 31634 8520
rect 28077 8483 28135 8489
rect 28077 8480 28089 8483
rect 27764 8452 28089 8480
rect 27764 8440 27770 8452
rect 28077 8449 28089 8452
rect 28123 8449 28135 8483
rect 28077 8443 28135 8449
rect 28261 8483 28319 8489
rect 28261 8449 28273 8483
rect 28307 8449 28319 8483
rect 28261 8443 28319 8449
rect 28353 8483 28411 8489
rect 28353 8449 28365 8483
rect 28399 8449 28411 8483
rect 28353 8443 28411 8449
rect 28445 8483 28503 8489
rect 28445 8449 28457 8483
rect 28491 8480 28503 8483
rect 29086 8480 29092 8492
rect 28491 8452 29092 8480
rect 28491 8449 28503 8452
rect 28445 8443 28503 8449
rect 25556 8384 26096 8412
rect 25556 8372 25562 8384
rect 28166 8372 28172 8424
rect 28224 8412 28230 8424
rect 28368 8412 28396 8443
rect 29086 8440 29092 8452
rect 29144 8440 29150 8492
rect 31754 8480 31760 8492
rect 29196 8452 31760 8480
rect 28224 8384 28396 8412
rect 28224 8372 28230 8384
rect 24486 8304 24492 8356
rect 24544 8344 24550 8356
rect 29196 8344 29224 8452
rect 31754 8440 31760 8452
rect 31812 8480 31818 8492
rect 32306 8480 32312 8492
rect 31812 8452 32312 8480
rect 31812 8440 31818 8452
rect 32306 8440 32312 8452
rect 32364 8440 32370 8492
rect 32401 8483 32459 8489
rect 32401 8449 32413 8483
rect 32447 8449 32459 8483
rect 32401 8443 32459 8449
rect 30745 8415 30803 8421
rect 30745 8381 30757 8415
rect 30791 8412 30803 8415
rect 30926 8412 30932 8424
rect 30791 8384 30932 8412
rect 30791 8381 30803 8384
rect 30745 8375 30803 8381
rect 30926 8372 30932 8384
rect 30984 8372 30990 8424
rect 24544 8316 29224 8344
rect 32416 8344 32444 8443
rect 32490 8440 32496 8492
rect 32548 8480 32554 8492
rect 32692 8489 32720 8520
rect 32766 8508 32772 8560
rect 32824 8548 32830 8560
rect 33781 8551 33839 8557
rect 33781 8548 33793 8551
rect 32824 8520 33793 8548
rect 32824 8508 32830 8520
rect 33781 8517 33793 8520
rect 33827 8548 33839 8551
rect 35250 8548 35256 8560
rect 33827 8520 35256 8548
rect 33827 8517 33839 8520
rect 33781 8511 33839 8517
rect 35250 8508 35256 8520
rect 35308 8508 35314 8560
rect 35728 8557 35756 8588
rect 37369 8585 37381 8588
rect 37415 8585 37427 8619
rect 37369 8579 37427 8585
rect 35713 8551 35771 8557
rect 35713 8517 35725 8551
rect 35759 8517 35771 8551
rect 36354 8548 36360 8560
rect 36315 8520 36360 8548
rect 35713 8511 35771 8517
rect 36354 8508 36360 8520
rect 36412 8508 36418 8560
rect 32677 8483 32735 8489
rect 32548 8452 32593 8480
rect 32548 8440 32554 8452
rect 32677 8449 32689 8483
rect 32723 8449 32735 8483
rect 32677 8443 32735 8449
rect 33597 8483 33655 8489
rect 33597 8449 33609 8483
rect 33643 8480 33655 8483
rect 34146 8480 34152 8492
rect 33643 8452 34152 8480
rect 33643 8449 33655 8452
rect 33597 8443 33655 8449
rect 34146 8440 34152 8452
rect 34204 8440 34210 8492
rect 35526 8480 35532 8492
rect 35487 8452 35532 8480
rect 35526 8440 35532 8452
rect 35584 8440 35590 8492
rect 37274 8440 37280 8492
rect 37332 8480 37338 8492
rect 38482 8483 38540 8489
rect 38482 8480 38494 8483
rect 37332 8452 38494 8480
rect 37332 8440 37338 8452
rect 38482 8449 38494 8452
rect 38528 8449 38540 8483
rect 38482 8443 38540 8449
rect 38749 8483 38807 8489
rect 38749 8449 38761 8483
rect 38795 8480 38807 8483
rect 38838 8480 38844 8492
rect 38795 8452 38844 8480
rect 38795 8449 38807 8452
rect 38749 8443 38807 8449
rect 38838 8440 38844 8452
rect 38896 8440 38902 8492
rect 33962 8344 33968 8356
rect 32416 8316 33968 8344
rect 24544 8304 24550 8316
rect 33962 8304 33968 8316
rect 34020 8304 34026 8356
rect 18748 8248 19104 8276
rect 18748 8236 18754 8248
rect 25038 8236 25044 8288
rect 25096 8276 25102 8288
rect 25133 8279 25191 8285
rect 25133 8276 25145 8279
rect 25096 8248 25145 8276
rect 25096 8236 25102 8248
rect 25133 8245 25145 8248
rect 25179 8245 25191 8279
rect 25133 8239 25191 8245
rect 35897 8279 35955 8285
rect 35897 8245 35909 8279
rect 35943 8276 35955 8279
rect 36262 8276 36268 8288
rect 35943 8248 36268 8276
rect 35943 8245 35955 8248
rect 35897 8239 35955 8245
rect 36262 8236 36268 8248
rect 36320 8236 36326 8288
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 3142 8072 3148 8084
rect 3055 8044 3148 8072
rect 3142 8032 3148 8044
rect 3200 8072 3206 8084
rect 3878 8072 3884 8084
rect 3200 8044 3884 8072
rect 3200 8032 3206 8044
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 13265 8075 13323 8081
rect 9232 8044 13216 8072
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 9232 7945 9260 8044
rect 11882 8004 11888 8016
rect 10336 7976 11888 8004
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 5592 7908 5733 7936
rect 5592 7896 5598 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 7975 7908 9229 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5123 7840 6316 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 2501 7803 2559 7809
rect 2501 7800 2513 7803
rect 2188 7772 2513 7800
rect 2188 7760 2194 7772
rect 2501 7769 2513 7772
rect 2547 7769 2559 7803
rect 5966 7803 6024 7809
rect 5966 7800 5978 7803
rect 2501 7763 2559 7769
rect 5276 7772 5978 7800
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 2406 7732 2412 7744
rect 2087 7704 2412 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 3878 7732 3884 7744
rect 3839 7704 3884 7732
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4617 7735 4675 7741
rect 4617 7701 4629 7735
rect 4663 7732 4675 7735
rect 5074 7732 5080 7744
rect 4663 7704 5080 7732
rect 4663 7701 4675 7704
rect 4617 7695 4675 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5276 7741 5304 7772
rect 5966 7769 5978 7772
rect 6012 7769 6024 7803
rect 6288 7800 6316 7840
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7432 7840 7757 7868
rect 7432 7828 7438 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 10226 7868 10232 7880
rect 8987 7840 10232 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 7561 7803 7619 7809
rect 7561 7800 7573 7803
rect 6288 7772 7573 7800
rect 5966 7763 6024 7769
rect 7561 7769 7573 7772
rect 7607 7769 7619 7803
rect 7561 7763 7619 7769
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7701 5319 7735
rect 5261 7695 5319 7701
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 7834 7732 7840 7744
rect 7147 7704 7840 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 10336 7732 10364 7976
rect 11882 7964 11888 7976
rect 11940 7964 11946 8016
rect 13188 8004 13216 8044
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 13998 8072 14004 8084
rect 13311 8044 14004 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 16816 8044 18092 8072
rect 16816 8032 16822 8044
rect 14458 8004 14464 8016
rect 13188 7976 14464 8004
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 14829 8007 14887 8013
rect 14829 7973 14841 8007
rect 14875 8004 14887 8007
rect 16298 8004 16304 8016
rect 14875 7976 16304 8004
rect 14875 7973 14887 7976
rect 14829 7967 14887 7973
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 17770 7964 17776 8016
rect 17828 8004 17834 8016
rect 17828 7976 17908 8004
rect 17828 7964 17834 7976
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 12805 7939 12863 7945
rect 12805 7936 12817 7939
rect 11112 7908 12817 7936
rect 11112 7896 11118 7908
rect 12805 7905 12817 7908
rect 12851 7905 12863 7939
rect 14476 7936 14504 7964
rect 17880 7945 17908 7976
rect 17865 7939 17923 7945
rect 14476 7908 15608 7936
rect 12805 7899 12863 7905
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 10888 7840 11253 7868
rect 10888 7812 10916 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11882 7868 11888 7880
rect 11843 7840 11888 7868
rect 11241 7831 11299 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 12526 7868 12532 7880
rect 12487 7840 12532 7868
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12710 7868 12716 7880
rect 12671 7840 12716 7868
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 13078 7868 13084 7880
rect 13039 7840 13084 7868
rect 12897 7831 12955 7837
rect 10597 7803 10655 7809
rect 10597 7769 10609 7803
rect 10643 7800 10655 7803
rect 10870 7800 10876 7812
rect 10643 7772 10876 7800
rect 10643 7769 10655 7772
rect 10597 7763 10655 7769
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 12912 7800 12940 7831
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15580 7868 15608 7908
rect 17865 7905 17877 7939
rect 17911 7905 17923 7939
rect 17865 7899 17923 7905
rect 17586 7868 17592 7880
rect 15580 7840 17592 7868
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17957 7871 18015 7877
rect 17773 7865 17831 7871
rect 17773 7831 17785 7865
rect 17819 7831 17831 7865
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 18064 7868 18092 8044
rect 26050 8032 26056 8084
rect 26108 8072 26114 8084
rect 26878 8072 26884 8084
rect 26108 8044 26884 8072
rect 26108 8032 26114 8044
rect 26878 8032 26884 8044
rect 26936 8072 26942 8084
rect 26973 8075 27031 8081
rect 26973 8072 26985 8075
rect 26936 8044 26985 8072
rect 26936 8032 26942 8044
rect 26973 8041 26985 8044
rect 27019 8072 27031 8075
rect 28534 8072 28540 8084
rect 27019 8044 28540 8072
rect 27019 8041 27031 8044
rect 26973 8035 27031 8041
rect 28534 8032 28540 8044
rect 28592 8032 28598 8084
rect 28905 8075 28963 8081
rect 28905 8041 28917 8075
rect 28951 8072 28963 8075
rect 29086 8072 29092 8084
rect 28951 8044 29092 8072
rect 28951 8041 28963 8044
rect 28905 8035 28963 8041
rect 29086 8032 29092 8044
rect 29144 8032 29150 8084
rect 31018 8032 31024 8084
rect 31076 8072 31082 8084
rect 31481 8075 31539 8081
rect 31481 8072 31493 8075
rect 31076 8044 31493 8072
rect 31076 8032 31082 8044
rect 31481 8041 31493 8044
rect 31527 8041 31539 8075
rect 31481 8035 31539 8041
rect 33413 8075 33471 8081
rect 33413 8041 33425 8075
rect 33459 8072 33471 8075
rect 33686 8072 33692 8084
rect 33459 8044 33692 8072
rect 33459 8041 33471 8044
rect 33413 8035 33471 8041
rect 33686 8032 33692 8044
rect 33744 8032 33750 8084
rect 34149 8075 34207 8081
rect 34149 8041 34161 8075
rect 34195 8072 34207 8075
rect 34514 8072 34520 8084
rect 34195 8044 34520 8072
rect 34195 8041 34207 8044
rect 34149 8035 34207 8041
rect 34514 8032 34520 8044
rect 34572 8072 34578 8084
rect 35526 8072 35532 8084
rect 34572 8044 35532 8072
rect 34572 8032 34578 8044
rect 35526 8032 35532 8044
rect 35584 8032 35590 8084
rect 36817 8075 36875 8081
rect 36188 8044 36768 8072
rect 22281 8007 22339 8013
rect 22281 7973 22293 8007
rect 22327 8004 22339 8007
rect 30466 8004 30472 8016
rect 22327 7976 30472 8004
rect 22327 7973 22339 7976
rect 22281 7967 22339 7973
rect 30466 7964 30472 7976
rect 30524 7964 30530 8016
rect 20349 7939 20407 7945
rect 20349 7905 20361 7939
rect 20395 7936 20407 7939
rect 20714 7936 20720 7948
rect 20395 7908 20720 7936
rect 20395 7905 20407 7908
rect 20349 7899 20407 7905
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 27706 7936 27712 7948
rect 25332 7908 27712 7936
rect 25332 7880 25360 7908
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 18064 7840 18153 7868
rect 17957 7831 18015 7837
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7868 20131 7871
rect 20162 7868 20168 7880
rect 20119 7840 20168 7868
rect 20119 7837 20131 7840
rect 20073 7831 20131 7837
rect 17773 7825 17831 7831
rect 13538 7800 13544 7812
rect 11204 7772 13544 7800
rect 11204 7760 11210 7772
rect 13538 7760 13544 7772
rect 13596 7760 13602 7812
rect 14645 7803 14703 7809
rect 14645 7769 14657 7803
rect 14691 7800 14703 7803
rect 14826 7800 14832 7812
rect 14691 7772 14832 7800
rect 14691 7769 14703 7772
rect 14645 7763 14703 7769
rect 14826 7760 14832 7772
rect 14884 7760 14890 7812
rect 8996 7704 10364 7732
rect 8996 7692 9002 7704
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10836 7704 11069 7732
rect 10836 7692 10842 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12250 7732 12256 7744
rect 12023 7704 12256 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12250 7692 12256 7704
rect 12308 7732 12314 7744
rect 12526 7732 12532 7744
rect 12308 7704 12532 7732
rect 12308 7692 12314 7704
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 14274 7692 14280 7744
rect 14332 7732 14338 7744
rect 15654 7732 15660 7744
rect 14332 7704 15660 7732
rect 14332 7692 14338 7704
rect 15654 7692 15660 7704
rect 15712 7732 15718 7744
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 15712 7704 16589 7732
rect 15712 7692 15718 7704
rect 16577 7701 16589 7704
rect 16623 7732 16635 7735
rect 17218 7732 17224 7744
rect 16623 7704 17224 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 17788 7732 17816 7825
rect 17972 7800 18000 7831
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 21450 7868 21456 7880
rect 21411 7840 21456 7868
rect 21450 7828 21456 7840
rect 21508 7868 21514 7880
rect 22002 7868 22008 7880
rect 21508 7840 22008 7868
rect 21508 7828 21514 7840
rect 22002 7828 22008 7840
rect 22060 7828 22066 7880
rect 22186 7868 22192 7880
rect 22147 7840 22192 7868
rect 22186 7828 22192 7840
rect 22244 7828 22250 7880
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7837 25007 7871
rect 24949 7831 25007 7837
rect 25041 7871 25099 7877
rect 25041 7837 25053 7871
rect 25087 7837 25099 7871
rect 25041 7831 25099 7837
rect 18414 7800 18420 7812
rect 17972 7772 18420 7800
rect 18414 7760 18420 7772
rect 18472 7760 18478 7812
rect 17862 7732 17868 7744
rect 17788 7704 17868 7732
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 18325 7735 18383 7741
rect 18325 7732 18337 7735
rect 18288 7704 18337 7732
rect 18288 7692 18294 7704
rect 18325 7701 18337 7704
rect 18371 7701 18383 7735
rect 24670 7732 24676 7744
rect 24631 7704 24676 7732
rect 18325 7695 18383 7701
rect 24670 7692 24676 7704
rect 24728 7692 24734 7744
rect 24964 7732 24992 7831
rect 25056 7800 25084 7831
rect 25130 7828 25136 7880
rect 25188 7868 25194 7880
rect 25188 7840 25233 7868
rect 25188 7828 25194 7840
rect 25314 7828 25320 7880
rect 25372 7868 25378 7880
rect 26050 7868 26056 7880
rect 25372 7840 25417 7868
rect 26011 7840 26056 7868
rect 25372 7828 25378 7840
rect 26050 7828 26056 7840
rect 26108 7828 26114 7880
rect 26145 7871 26203 7877
rect 26145 7837 26157 7871
rect 26191 7837 26203 7871
rect 26145 7831 26203 7837
rect 25222 7800 25228 7812
rect 25056 7772 25228 7800
rect 25222 7760 25228 7772
rect 25280 7800 25286 7812
rect 26160 7800 26188 7831
rect 26234 7828 26240 7880
rect 26292 7868 26298 7880
rect 26436 7877 26464 7908
rect 27706 7896 27712 7908
rect 27764 7936 27770 7948
rect 27764 7908 28212 7936
rect 27764 7896 27770 7908
rect 26421 7871 26479 7877
rect 26292 7840 26337 7868
rect 26292 7828 26298 7840
rect 26421 7837 26433 7871
rect 26467 7837 26479 7871
rect 27798 7868 27804 7880
rect 27759 7840 27804 7868
rect 26421 7831 26479 7837
rect 27798 7828 27804 7840
rect 27856 7828 27862 7880
rect 27893 7871 27951 7877
rect 27893 7837 27905 7871
rect 27939 7837 27951 7871
rect 27893 7831 27951 7837
rect 27908 7800 27936 7831
rect 27982 7828 27988 7880
rect 28040 7868 28046 7880
rect 28184 7877 28212 7908
rect 31018 7896 31024 7948
rect 31076 7936 31082 7948
rect 31076 7908 32076 7936
rect 31076 7896 31082 7908
rect 28169 7871 28227 7877
rect 28040 7840 28085 7868
rect 28040 7828 28046 7840
rect 28169 7837 28181 7871
rect 28215 7837 28227 7871
rect 31662 7868 31668 7880
rect 31623 7840 31668 7868
rect 28169 7831 28227 7837
rect 31662 7828 31668 7840
rect 31720 7828 31726 7880
rect 32048 7877 32076 7908
rect 32766 7896 32772 7948
rect 32824 7936 32830 7948
rect 35345 7939 35403 7945
rect 35345 7936 35357 7939
rect 32824 7908 35357 7936
rect 32824 7896 32830 7908
rect 35345 7905 35357 7908
rect 35391 7905 35403 7939
rect 35618 7936 35624 7948
rect 35579 7908 35624 7936
rect 35345 7899 35403 7905
rect 32033 7871 32091 7877
rect 32033 7837 32045 7871
rect 32079 7837 32091 7871
rect 32033 7831 32091 7837
rect 33965 7871 34023 7877
rect 33965 7837 33977 7871
rect 34011 7868 34023 7871
rect 34422 7868 34428 7880
rect 34011 7840 34428 7868
rect 34011 7837 34023 7840
rect 33965 7831 34023 7837
rect 34422 7828 34428 7840
rect 34480 7828 34486 7880
rect 28074 7800 28080 7812
rect 25280 7772 28080 7800
rect 25280 7760 25286 7772
rect 28074 7760 28080 7772
rect 28132 7760 28138 7812
rect 31757 7803 31815 7809
rect 31757 7769 31769 7803
rect 31803 7769 31815 7803
rect 31757 7763 31815 7769
rect 25038 7732 25044 7744
rect 24964 7704 25044 7732
rect 25038 7692 25044 7704
rect 25096 7692 25102 7744
rect 25682 7692 25688 7744
rect 25740 7732 25746 7744
rect 25777 7735 25835 7741
rect 25777 7732 25789 7735
rect 25740 7704 25789 7732
rect 25740 7692 25746 7704
rect 25777 7701 25789 7704
rect 25823 7701 25835 7735
rect 25777 7695 25835 7701
rect 27525 7735 27583 7741
rect 27525 7701 27537 7735
rect 27571 7732 27583 7735
rect 28350 7732 28356 7744
rect 27571 7704 28356 7732
rect 27571 7701 27583 7704
rect 27525 7695 27583 7701
rect 28350 7692 28356 7704
rect 28408 7692 28414 7744
rect 31772 7732 31800 7763
rect 31846 7760 31852 7812
rect 31904 7800 31910 7812
rect 32490 7800 32496 7812
rect 31904 7772 32496 7800
rect 31904 7760 31910 7772
rect 32490 7760 32496 7772
rect 32548 7760 32554 7812
rect 35360 7800 35388 7899
rect 35618 7896 35624 7908
rect 35676 7896 35682 7948
rect 35894 7828 35900 7880
rect 35952 7868 35958 7880
rect 36188 7877 36216 8044
rect 36354 7964 36360 8016
rect 36412 7964 36418 8016
rect 36740 8004 36768 8044
rect 36817 8041 36829 8075
rect 36863 8072 36875 8075
rect 37274 8072 37280 8084
rect 36863 8044 37280 8072
rect 36863 8041 36875 8044
rect 36817 8035 36875 8041
rect 37274 8032 37280 8044
rect 37332 8032 37338 8084
rect 40494 8004 40500 8016
rect 36740 7976 40500 8004
rect 40494 7964 40500 7976
rect 40552 7964 40558 8016
rect 36372 7936 36400 7964
rect 36372 7908 36584 7936
rect 36173 7871 36231 7877
rect 36173 7868 36185 7871
rect 35952 7840 36185 7868
rect 35952 7828 35958 7840
rect 36173 7837 36185 7840
rect 36219 7837 36231 7871
rect 36173 7831 36231 7837
rect 36262 7828 36268 7880
rect 36320 7868 36326 7880
rect 36556 7877 36584 7908
rect 36357 7871 36415 7877
rect 36541 7871 36599 7877
rect 36357 7868 36369 7871
rect 36320 7840 36369 7868
rect 36320 7828 36326 7840
rect 36357 7837 36369 7840
rect 36403 7837 36415 7871
rect 36357 7831 36415 7837
rect 36452 7865 36510 7871
rect 36452 7831 36464 7865
rect 36498 7831 36510 7865
rect 36541 7837 36553 7871
rect 36587 7837 36599 7871
rect 68094 7868 68100 7880
rect 68055 7840 68100 7868
rect 36541 7831 36599 7837
rect 36452 7825 36510 7831
rect 68094 7828 68100 7840
rect 68152 7828 68158 7880
rect 35360 7772 35894 7800
rect 33226 7732 33232 7744
rect 31772 7704 33232 7732
rect 33226 7692 33232 7704
rect 33284 7692 33290 7744
rect 35866 7732 35894 7772
rect 36170 7732 36176 7744
rect 35866 7704 36176 7732
rect 36170 7692 36176 7704
rect 36228 7732 36234 7744
rect 36473 7732 36501 7825
rect 36228 7704 36501 7732
rect 36228 7692 36234 7704
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 7374 7528 7380 7540
rect 2455 7500 2774 7528
rect 7335 7500 7380 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2746 7460 2774 7500
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 7834 7528 7840 7540
rect 7795 7500 7840 7528
rect 7834 7488 7840 7500
rect 7892 7528 7898 7540
rect 9306 7528 9312 7540
rect 7892 7500 9312 7528
rect 7892 7488 7898 7500
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 12894 7528 12900 7540
rect 10192 7500 12900 7528
rect 10192 7488 10198 7500
rect 12894 7488 12900 7500
rect 12952 7528 12958 7540
rect 14274 7528 14280 7540
rect 12952 7500 14280 7528
rect 12952 7488 12958 7500
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 18414 7528 18420 7540
rect 14884 7500 18420 7528
rect 14884 7488 14890 7500
rect 18414 7488 18420 7500
rect 18472 7528 18478 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 18472 7500 20085 7528
rect 18472 7488 18478 7500
rect 20073 7497 20085 7500
rect 20119 7497 20131 7531
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 20073 7491 20131 7497
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 26234 7488 26240 7540
rect 26292 7528 26298 7540
rect 26421 7531 26479 7537
rect 26421 7528 26433 7531
rect 26292 7500 26433 7528
rect 26292 7488 26298 7500
rect 26421 7497 26433 7500
rect 26467 7497 26479 7531
rect 26421 7491 26479 7497
rect 27801 7531 27859 7537
rect 27801 7497 27813 7531
rect 27847 7528 27859 7531
rect 27982 7528 27988 7540
rect 27847 7500 27988 7528
rect 27847 7497 27859 7500
rect 27801 7491 27859 7497
rect 27982 7488 27988 7500
rect 28040 7488 28046 7540
rect 29086 7488 29092 7540
rect 29144 7528 29150 7540
rect 36262 7528 36268 7540
rect 29144 7500 36268 7528
rect 29144 7488 29150 7500
rect 36262 7488 36268 7500
rect 36320 7488 36326 7540
rect 36354 7488 36360 7540
rect 36412 7528 36418 7540
rect 37829 7531 37887 7537
rect 37829 7528 37841 7531
rect 36412 7500 37841 7528
rect 36412 7488 36418 7500
rect 37829 7497 37841 7500
rect 37875 7497 37887 7531
rect 37829 7491 37887 7497
rect 3390 7463 3448 7469
rect 3390 7460 3402 7463
rect 2746 7432 3402 7460
rect 3390 7429 3402 7432
rect 3436 7429 3448 7463
rect 3390 7423 3448 7429
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 8294 7460 8300 7472
rect 5675 7432 8300 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 9892 7463 9950 7469
rect 9892 7429 9904 7463
rect 9938 7460 9950 7463
rect 11885 7463 11943 7469
rect 11885 7460 11897 7463
rect 9938 7432 11897 7460
rect 9938 7429 9950 7432
rect 9892 7423 9950 7429
rect 11885 7429 11897 7432
rect 11931 7429 11943 7463
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 11885 7423 11943 7429
rect 12452 7432 20729 7460
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6512 7364 6929 7392
rect 6512 7352 6518 7364
rect 6917 7361 6929 7364
rect 6963 7392 6975 7395
rect 7742 7392 7748 7404
rect 6963 7364 7748 7392
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 10134 7392 10140 7404
rect 10095 7364 10140 7392
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10781 7395 10839 7401
rect 12161 7395 12219 7401
rect 10781 7392 10793 7395
rect 10652 7364 10793 7392
rect 10652 7352 10658 7364
rect 10781 7361 10793 7364
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 12047 7367 12173 7395
rect 3142 7324 3148 7336
rect 3103 7296 3148 7324
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 4982 7324 4988 7336
rect 4943 7296 4988 7324
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7293 5411 7327
rect 5353 7287 5411 7293
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 3050 7256 3056 7268
rect 1811 7228 3056 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 3050 7216 3056 7228
rect 3108 7216 3114 7268
rect 5368 7256 5396 7287
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5500 7296 5545 7324
rect 5500 7284 5506 7296
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 7929 7327 7987 7333
rect 7929 7324 7941 7327
rect 7248 7296 7941 7324
rect 7248 7284 7254 7296
rect 7929 7293 7941 7296
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 12047 7256 12075 7367
rect 12161 7361 12173 7367
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12250 7395 12308 7401
rect 12250 7361 12262 7395
rect 12296 7361 12308 7395
rect 12250 7355 12308 7361
rect 12366 7395 12424 7401
rect 12366 7361 12378 7395
rect 12412 7392 12424 7395
rect 12452 7392 12480 7432
rect 20717 7429 20729 7432
rect 20763 7429 20775 7463
rect 21192 7460 21220 7488
rect 23934 7460 23940 7472
rect 21192 7432 21864 7460
rect 23895 7432 23940 7460
rect 20717 7423 20775 7429
rect 12412 7364 12480 7392
rect 12412 7361 12424 7364
rect 12366 7355 12424 7361
rect 12268 7324 12296 7355
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 12584 7364 12629 7392
rect 12584 7352 12590 7364
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13228 7364 14289 7392
rect 13228 7352 13234 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7392 14611 7395
rect 14826 7392 14832 7404
rect 14599 7364 14832 7392
rect 14599 7361 14611 7364
rect 14553 7355 14611 7361
rect 13538 7324 13544 7336
rect 12268 7296 13544 7324
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7324 13875 7327
rect 14568 7324 14596 7355
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 18230 7352 18236 7404
rect 18288 7401 18294 7404
rect 18288 7392 18300 7401
rect 20441 7395 20499 7401
rect 18288 7364 18333 7392
rect 18288 7355 18300 7364
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 21266 7392 21272 7404
rect 20487 7364 21272 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 18288 7352 18294 7355
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 21836 7401 21864 7432
rect 23934 7420 23940 7432
rect 23992 7420 23998 7472
rect 25593 7463 25651 7469
rect 25593 7429 25605 7463
rect 25639 7460 25651 7463
rect 26326 7460 26332 7472
rect 25639 7432 26332 7460
rect 25639 7429 25651 7432
rect 25593 7423 25651 7429
rect 26326 7420 26332 7432
rect 26384 7420 26390 7472
rect 27614 7460 27620 7472
rect 27575 7432 27620 7460
rect 27614 7420 27620 7432
rect 27672 7420 27678 7472
rect 30929 7463 30987 7469
rect 30929 7429 30941 7463
rect 30975 7460 30987 7463
rect 31018 7460 31024 7472
rect 30975 7432 31024 7460
rect 30975 7429 30987 7432
rect 30929 7423 30987 7429
rect 31018 7420 31024 7432
rect 31076 7420 31082 7472
rect 31938 7420 31944 7472
rect 31996 7460 32002 7472
rect 32398 7460 32404 7472
rect 31996 7432 32404 7460
rect 31996 7420 32002 7432
rect 32398 7420 32404 7432
rect 32456 7460 32462 7472
rect 32585 7463 32643 7469
rect 32585 7460 32597 7463
rect 32456 7432 32597 7460
rect 32456 7420 32462 7432
rect 32585 7429 32597 7432
rect 32631 7429 32643 7463
rect 32585 7423 32643 7429
rect 32769 7463 32827 7469
rect 32769 7429 32781 7463
rect 32815 7460 32827 7463
rect 34514 7460 34520 7472
rect 32815 7432 34520 7460
rect 32815 7429 32827 7432
rect 32769 7423 32827 7429
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7361 21879 7395
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21821 7355 21879 7361
rect 21928 7364 22017 7392
rect 13863 7296 14596 7324
rect 18509 7327 18567 7333
rect 13863 7293 13875 7296
rect 13817 7287 13875 7293
rect 18509 7293 18521 7327
rect 18555 7324 18567 7327
rect 18598 7324 18604 7336
rect 18555 7296 18604 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 15562 7256 15568 7268
rect 4632 7228 5396 7256
rect 10152 7228 15568 7256
rect 4632 7200 4660 7228
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 4614 7188 4620 7200
rect 4571 7160 4620 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 8757 7191 8815 7197
rect 8757 7157 8769 7191
rect 8803 7188 8815 7191
rect 10152 7188 10180 7228
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 8803 7160 10180 7188
rect 10965 7191 11023 7197
rect 8803 7157 8815 7160
rect 8757 7151 8815 7157
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11514 7188 11520 7200
rect 11011 7160 11520 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 16117 7191 16175 7197
rect 16117 7157 16129 7191
rect 16163 7188 16175 7191
rect 16390 7188 16396 7200
rect 16163 7160 16396 7188
rect 16163 7157 16175 7160
rect 16117 7151 16175 7157
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 16816 7160 17141 7188
rect 16816 7148 16822 7160
rect 17129 7157 17141 7160
rect 17175 7157 17187 7191
rect 17129 7151 17187 7157
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 18524 7188 18552 7287
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 18966 7284 18972 7336
rect 19024 7284 19030 7336
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7324 20591 7327
rect 20714 7324 20720 7336
rect 20579 7296 20720 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 18984 7256 19012 7284
rect 21928 7256 21956 7364
rect 22005 7361 22017 7364
rect 22051 7392 22063 7395
rect 22186 7392 22192 7404
rect 22051 7364 22192 7392
rect 22051 7361 22063 7364
rect 22005 7355 22063 7361
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 26053 7395 26111 7401
rect 26053 7392 26065 7395
rect 24912 7364 26065 7392
rect 24912 7352 24918 7364
rect 26053 7361 26065 7364
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 26237 7395 26295 7401
rect 26237 7361 26249 7395
rect 26283 7392 26295 7395
rect 26418 7392 26424 7404
rect 26283 7364 26424 7392
rect 26283 7361 26295 7364
rect 26237 7355 26295 7361
rect 26068 7324 26096 7355
rect 26418 7352 26424 7364
rect 26476 7352 26482 7404
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 31113 7395 31171 7401
rect 31113 7361 31125 7395
rect 31159 7392 31171 7395
rect 31386 7392 31392 7404
rect 31159 7364 31392 7392
rect 31159 7361 31171 7364
rect 31113 7355 31171 7361
rect 27246 7324 27252 7336
rect 26068 7296 27252 7324
rect 27246 7284 27252 7296
rect 27304 7324 27310 7336
rect 27448 7324 27476 7355
rect 31386 7352 31392 7364
rect 31444 7392 31450 7404
rect 32784 7392 32812 7423
rect 34514 7420 34520 7432
rect 34572 7420 34578 7472
rect 36277 7460 36305 7488
rect 36277 7432 36400 7460
rect 31444 7364 32812 7392
rect 33781 7395 33839 7401
rect 31444 7352 31450 7364
rect 33781 7361 33793 7395
rect 33827 7392 33839 7395
rect 34146 7392 34152 7404
rect 33827 7364 34152 7392
rect 33827 7361 33839 7364
rect 33781 7355 33839 7361
rect 34146 7352 34152 7364
rect 34204 7352 34210 7404
rect 34606 7352 34612 7404
rect 34664 7392 34670 7404
rect 35253 7395 35311 7401
rect 35253 7392 35265 7395
rect 34664 7364 35265 7392
rect 34664 7352 34670 7364
rect 35253 7361 35265 7364
rect 35299 7361 35311 7395
rect 35894 7392 35900 7404
rect 35855 7364 35900 7392
rect 35253 7355 35311 7361
rect 35894 7352 35900 7364
rect 35952 7352 35958 7404
rect 36078 7401 36084 7404
rect 36076 7392 36084 7401
rect 36039 7364 36084 7392
rect 36076 7355 36084 7364
rect 36078 7352 36084 7355
rect 36136 7352 36142 7404
rect 36176 7398 36234 7404
rect 36176 7364 36188 7398
rect 36222 7364 36234 7398
rect 36176 7358 36234 7364
rect 36285 7395 36343 7401
rect 36285 7361 36297 7395
rect 36331 7392 36343 7395
rect 36372 7392 36400 7432
rect 36331 7364 36400 7392
rect 37844 7392 37872 7491
rect 38657 7395 38715 7401
rect 38657 7392 38669 7395
rect 37844 7364 38669 7392
rect 36331 7361 36343 7364
rect 27304 7296 27476 7324
rect 34977 7327 35035 7333
rect 27304 7284 27310 7296
rect 34977 7293 34989 7327
rect 35023 7293 35035 7327
rect 36188 7324 36216 7358
rect 36285 7355 36343 7361
rect 38657 7361 38669 7364
rect 38703 7361 38715 7395
rect 38657 7355 38715 7361
rect 38749 7395 38807 7401
rect 38749 7361 38761 7395
rect 38795 7361 38807 7395
rect 38749 7355 38807 7361
rect 34977 7287 35035 7293
rect 36096 7296 36216 7324
rect 18984 7228 21956 7256
rect 22097 7259 22155 7265
rect 22097 7225 22109 7259
rect 22143 7256 22155 7259
rect 31846 7256 31852 7268
rect 22143 7228 31852 7256
rect 22143 7225 22155 7228
rect 22097 7219 22155 7225
rect 31846 7216 31852 7228
rect 31904 7216 31910 7268
rect 17276 7160 18552 7188
rect 17276 7148 17282 7160
rect 18782 7148 18788 7200
rect 18840 7188 18846 7200
rect 18969 7191 19027 7197
rect 18969 7188 18981 7191
rect 18840 7160 18981 7188
rect 18840 7148 18846 7160
rect 18969 7157 18981 7160
rect 19015 7157 19027 7191
rect 18969 7151 19027 7157
rect 20530 7148 20536 7200
rect 20588 7188 20594 7200
rect 22738 7188 22744 7200
rect 20588 7160 22744 7188
rect 20588 7148 20594 7160
rect 22738 7148 22744 7160
rect 22796 7188 22802 7200
rect 23293 7191 23351 7197
rect 23293 7188 23305 7191
rect 22796 7160 23305 7188
rect 22796 7148 22802 7160
rect 23293 7157 23305 7160
rect 23339 7188 23351 7191
rect 24762 7188 24768 7200
rect 23339 7160 24768 7188
rect 23339 7157 23351 7160
rect 23293 7151 23351 7157
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 27798 7148 27804 7200
rect 27856 7188 27862 7200
rect 28353 7191 28411 7197
rect 28353 7188 28365 7191
rect 27856 7160 28365 7188
rect 27856 7148 27862 7160
rect 28353 7157 28365 7160
rect 28399 7188 28411 7191
rect 28442 7188 28448 7200
rect 28399 7160 28448 7188
rect 28399 7157 28411 7160
rect 28353 7151 28411 7157
rect 28442 7148 28448 7160
rect 28500 7148 28506 7200
rect 28534 7148 28540 7200
rect 28592 7188 28598 7200
rect 30282 7188 30288 7200
rect 28592 7160 30288 7188
rect 28592 7148 28598 7160
rect 30282 7148 30288 7160
rect 30340 7148 30346 7200
rect 30745 7191 30803 7197
rect 30745 7157 30757 7191
rect 30791 7188 30803 7191
rect 31018 7188 31024 7200
rect 30791 7160 31024 7188
rect 30791 7157 30803 7160
rect 30745 7151 30803 7157
rect 31018 7148 31024 7160
rect 31076 7148 31082 7200
rect 32306 7148 32312 7200
rect 32364 7188 32370 7200
rect 32401 7191 32459 7197
rect 32401 7188 32413 7191
rect 32364 7160 32413 7188
rect 32364 7148 32370 7160
rect 32401 7157 32413 7160
rect 32447 7157 32459 7191
rect 32401 7151 32459 7157
rect 33502 7148 33508 7200
rect 33560 7188 33566 7200
rect 33965 7191 34023 7197
rect 33965 7188 33977 7191
rect 33560 7160 33977 7188
rect 33560 7148 33566 7160
rect 33965 7157 33977 7160
rect 34011 7157 34023 7191
rect 34992 7188 35020 7287
rect 36096 7268 36124 7296
rect 36078 7216 36084 7268
rect 36136 7216 36142 7268
rect 38764 7256 38792 7355
rect 38838 7352 38844 7404
rect 38896 7392 38902 7404
rect 38896 7364 38941 7392
rect 38896 7352 38902 7364
rect 39022 7352 39028 7404
rect 39080 7392 39086 7404
rect 39080 7364 39125 7392
rect 39080 7352 39086 7364
rect 36188 7228 38792 7256
rect 35618 7188 35624 7200
rect 34992 7160 35624 7188
rect 33965 7151 34023 7157
rect 35618 7148 35624 7160
rect 35676 7188 35682 7200
rect 36188 7188 36216 7228
rect 36538 7188 36544 7200
rect 35676 7160 36216 7188
rect 36499 7160 36544 7188
rect 35676 7148 35682 7160
rect 36538 7148 36544 7160
rect 36596 7148 36602 7200
rect 38378 7188 38384 7200
rect 38339 7160 38384 7188
rect 38378 7148 38384 7160
rect 38436 7148 38442 7200
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 4430 6944 4436 6996
rect 4488 6984 4494 6996
rect 10042 6984 10048 6996
rect 4488 6956 10048 6984
rect 4488 6944 4494 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10962 6984 10968 6996
rect 10520 6956 10968 6984
rect 10410 6916 10416 6928
rect 9140 6888 10416 6916
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 5166 6848 5172 6860
rect 3292 6820 5172 6848
rect 3292 6808 3298 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 5626 6848 5632 6860
rect 5587 6820 5632 6848
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 9140 6848 9168 6888
rect 10410 6876 10416 6888
rect 10468 6876 10474 6928
rect 9306 6848 9312 6860
rect 7239 6820 9168 6848
rect 9267 6820 9312 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 9824 6820 10149 6848
rect 9824 6808 9830 6820
rect 10137 6817 10149 6820
rect 10183 6848 10195 6851
rect 10226 6848 10232 6860
rect 10183 6820 10232 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 4614 6780 4620 6792
rect 2271 6752 4620 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5350 6780 5356 6792
rect 5311 6752 5356 6780
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 8202 6780 8208 6792
rect 5500 6752 5545 6780
rect 8163 6752 8208 6780
rect 5500 6740 5506 6752
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9674 6780 9680 6792
rect 9447 6752 9680 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 2133 6715 2191 6721
rect 2133 6681 2145 6715
rect 2179 6712 2191 6715
rect 2498 6712 2504 6724
rect 2179 6684 2504 6712
rect 2179 6681 2191 6684
rect 2133 6675 2191 6681
rect 2498 6672 2504 6684
rect 2556 6712 2562 6724
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2556 6684 2973 6712
rect 2556 6672 2562 6684
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 4525 6715 4583 6721
rect 4525 6681 4537 6715
rect 4571 6712 4583 6715
rect 4571 6684 5488 6712
rect 4571 6681 4583 6684
rect 4525 6675 4583 6681
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 1946 6644 1952 6656
rect 1811 6616 1952 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 4706 6644 4712 6656
rect 4019 6616 4712 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 4982 6644 4988 6656
rect 4943 6616 4988 6644
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5460 6644 5488 6684
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 9585 6715 9643 6721
rect 5592 6684 9260 6712
rect 5592 6672 5598 6684
rect 6546 6644 6552 6656
rect 5460 6616 6552 6644
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 6641 6647 6699 6653
rect 6641 6613 6653 6647
rect 6687 6644 6699 6647
rect 7466 6644 7472 6656
rect 6687 6616 7472 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 7745 6647 7803 6653
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 8294 6644 8300 6656
rect 7791 6616 8300 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8478 6644 8484 6656
rect 8435 6616 8484 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 8941 6647 8999 6653
rect 8941 6613 8953 6647
rect 8987 6644 8999 6647
rect 9122 6644 9128 6656
rect 8987 6616 9128 6644
rect 8987 6613 8999 6616
rect 8941 6607 8999 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9232 6644 9260 6684
rect 9585 6681 9597 6715
rect 9631 6712 9643 6715
rect 10520 6712 10548 6956
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 20254 6984 20260 6996
rect 12584 6956 20260 6984
rect 12584 6944 12590 6956
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 23842 6984 23848 6996
rect 23803 6956 23848 6984
rect 23842 6944 23848 6956
rect 23900 6944 23906 6996
rect 26418 6944 26424 6996
rect 26476 6984 26482 6996
rect 26789 6987 26847 6993
rect 26789 6984 26801 6987
rect 26476 6956 26801 6984
rect 26476 6944 26482 6956
rect 26789 6953 26801 6956
rect 26835 6953 26847 6987
rect 26789 6947 26847 6953
rect 30929 6987 30987 6993
rect 30929 6953 30941 6987
rect 30975 6984 30987 6987
rect 31110 6984 31116 6996
rect 30975 6956 31116 6984
rect 30975 6953 30987 6956
rect 30929 6947 30987 6953
rect 31110 6944 31116 6956
rect 31168 6944 31174 6996
rect 32398 6984 32404 6996
rect 32359 6956 32404 6984
rect 32398 6944 32404 6956
rect 32456 6944 32462 6996
rect 38838 6944 38844 6996
rect 38896 6984 38902 6996
rect 39117 6987 39175 6993
rect 39117 6984 39129 6987
rect 38896 6956 39129 6984
rect 38896 6944 38902 6956
rect 39117 6953 39129 6956
rect 39163 6953 39175 6987
rect 39117 6947 39175 6953
rect 11330 6876 11336 6928
rect 11388 6916 11394 6928
rect 12434 6916 12440 6928
rect 11388 6888 12440 6916
rect 11388 6876 11394 6888
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 14826 6876 14832 6928
rect 14884 6916 14890 6928
rect 14884 6888 14964 6916
rect 14884 6876 14890 6888
rect 10959 6851 11017 6857
rect 10959 6848 10971 6851
rect 10796 6820 10971 6848
rect 10686 6780 10692 6792
rect 10647 6752 10692 6780
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 9631 6684 10548 6712
rect 9631 6681 9643 6684
rect 9585 6675 9643 6681
rect 10796 6644 10824 6820
rect 10959 6817 10971 6820
rect 11005 6817 11017 6851
rect 10959 6811 11017 6817
rect 11146 6808 11152 6860
rect 11204 6808 11210 6860
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6848 12771 6851
rect 14274 6848 14280 6860
rect 12759 6820 14280 6848
rect 12759 6817 12771 6820
rect 12713 6811 12771 6817
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 14936 6857 14964 6888
rect 15102 6876 15108 6928
rect 15160 6876 15166 6928
rect 36262 6916 36268 6928
rect 36223 6888 36268 6916
rect 36262 6876 36268 6888
rect 36320 6876 36326 6928
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6817 14979 6851
rect 15120 6848 15148 6876
rect 17218 6848 17224 6860
rect 14921 6811 14979 6817
rect 15028 6820 15148 6848
rect 17179 6820 17224 6848
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6778 11115 6783
rect 11164 6778 11192 6808
rect 11103 6750 11192 6778
rect 11241 6783 11299 6789
rect 11103 6749 11115 6750
rect 11057 6743 11115 6749
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12618 6780 12624 6792
rect 11931 6752 12624 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 9232 6616 10824 6644
rect 10888 6644 10916 6743
rect 10962 6644 10968 6656
rect 10888 6616 10968 6644
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11256 6644 11284 6743
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13170 6780 13176 6792
rect 13131 6752 13176 6780
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 14516 6752 14565 6780
rect 14516 6740 14522 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14737 6783 14795 6789
rect 14737 6749 14749 6783
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 14752 6712 14780 6743
rect 14826 6740 14832 6792
rect 14884 6780 14890 6792
rect 14884 6752 14929 6780
rect 14884 6740 14890 6752
rect 15028 6712 15056 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 18598 6808 18604 6860
rect 18656 6848 18662 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 18656 6820 19257 6848
rect 18656 6808 18662 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 35526 6808 35532 6860
rect 35584 6808 35590 6860
rect 35713 6851 35771 6857
rect 35713 6817 35725 6851
rect 35759 6848 35771 6851
rect 35986 6848 35992 6860
rect 35759 6820 35992 6848
rect 35759 6817 35771 6820
rect 35713 6811 35771 6817
rect 35986 6808 35992 6820
rect 36044 6808 36050 6860
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 14752 6684 15056 6712
rect 11422 6644 11428 6656
rect 11204 6616 11284 6644
rect 11383 6616 11428 6644
rect 11204 6604 11210 6616
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6644 12127 6647
rect 12710 6644 12716 6656
rect 12115 6616 12716 6644
rect 12115 6613 12127 6616
rect 12069 6607 12127 6613
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 14090 6644 14096 6656
rect 13403 6616 14096 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 15120 6644 15148 6743
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 17957 6783 18015 6789
rect 17957 6780 17969 6783
rect 17644 6752 17969 6780
rect 17644 6740 17650 6752
rect 17957 6749 17969 6752
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 18104 6752 18153 6780
rect 18104 6740 18110 6752
rect 18141 6749 18153 6752
rect 18187 6749 18199 6783
rect 18233 6783 18291 6789
rect 18233 6770 18245 6783
rect 18279 6770 18291 6783
rect 18325 6783 18383 6789
rect 18141 6743 18199 6749
rect 15289 6715 15347 6721
rect 15289 6681 15301 6715
rect 15335 6712 15347 6715
rect 16954 6715 17012 6721
rect 18230 6718 18236 6770
rect 18288 6718 18294 6770
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18506 6780 18512 6792
rect 18467 6752 18512 6780
rect 18325 6743 18383 6749
rect 16954 6712 16966 6715
rect 15335 6684 16966 6712
rect 15335 6681 15347 6684
rect 15289 6675 15347 6681
rect 16954 6681 16966 6684
rect 17000 6681 17012 6715
rect 16954 6675 17012 6681
rect 15841 6647 15899 6653
rect 15841 6644 15853 6647
rect 15120 6616 15853 6644
rect 15841 6613 15853 6616
rect 15887 6644 15899 6647
rect 16022 6644 16028 6656
rect 15887 6616 16028 6644
rect 15887 6613 15899 6616
rect 15841 6607 15899 6613
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16298 6604 16304 6656
rect 16356 6644 16362 6656
rect 18340 6644 18368 6743
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 21266 6780 21272 6792
rect 21227 6752 21272 6780
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 22465 6783 22523 6789
rect 22465 6749 22477 6783
rect 22511 6780 22523 6783
rect 23474 6780 23480 6792
rect 22511 6752 23480 6780
rect 22511 6749 22523 6752
rect 22465 6743 22523 6749
rect 23474 6740 23480 6752
rect 23532 6780 23538 6792
rect 23934 6780 23940 6792
rect 23532 6752 23940 6780
rect 23532 6740 23538 6752
rect 23934 6740 23940 6752
rect 23992 6780 23998 6792
rect 25682 6789 25688 6792
rect 25409 6783 25467 6789
rect 25409 6780 25421 6783
rect 23992 6752 25421 6780
rect 23992 6740 23998 6752
rect 25409 6749 25421 6752
rect 25455 6749 25467 6783
rect 25676 6780 25688 6789
rect 25643 6752 25688 6780
rect 25409 6743 25467 6749
rect 25676 6743 25688 6752
rect 25682 6740 25688 6743
rect 25740 6740 25746 6792
rect 28350 6740 28356 6792
rect 28408 6789 28414 6792
rect 28408 6780 28420 6789
rect 28626 6780 28632 6792
rect 28408 6752 28453 6780
rect 28587 6752 28632 6780
rect 28408 6743 28420 6752
rect 28408 6740 28414 6743
rect 28626 6740 28632 6752
rect 28684 6780 28690 6792
rect 29546 6780 29552 6792
rect 28684 6752 29552 6780
rect 28684 6740 28690 6752
rect 29546 6740 29552 6752
rect 29604 6740 29610 6792
rect 30742 6780 30748 6792
rect 29748 6752 30748 6780
rect 18693 6715 18751 6721
rect 18693 6681 18705 6715
rect 18739 6712 18751 6715
rect 19490 6715 19548 6721
rect 19490 6712 19502 6715
rect 18739 6684 19502 6712
rect 18739 6681 18751 6684
rect 18693 6675 18751 6681
rect 19490 6681 19502 6684
rect 19536 6681 19548 6715
rect 19490 6675 19548 6681
rect 21453 6715 21511 6721
rect 21453 6681 21465 6715
rect 21499 6712 21511 6715
rect 21634 6712 21640 6724
rect 21499 6684 21640 6712
rect 21499 6681 21511 6684
rect 21453 6675 21511 6681
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 22732 6715 22790 6721
rect 22732 6681 22744 6715
rect 22778 6712 22790 6715
rect 24670 6712 24676 6724
rect 22778 6684 24676 6712
rect 22778 6681 22790 6684
rect 22732 6675 22790 6681
rect 24670 6672 24676 6684
rect 24728 6672 24734 6724
rect 24762 6672 24768 6724
rect 24820 6712 24826 6724
rect 24949 6715 25007 6721
rect 24820 6684 24865 6712
rect 24820 6672 24826 6684
rect 24949 6681 24961 6715
rect 24995 6712 25007 6715
rect 25038 6712 25044 6724
rect 24995 6684 25044 6712
rect 24995 6681 25007 6684
rect 24949 6675 25007 6681
rect 25038 6672 25044 6684
rect 25096 6712 25102 6724
rect 29748 6712 29776 6752
rect 30742 6740 30748 6752
rect 30800 6740 30806 6792
rect 30926 6740 30932 6792
rect 30984 6780 30990 6792
rect 33781 6783 33839 6789
rect 33781 6780 33793 6783
rect 30984 6752 33793 6780
rect 30984 6740 30990 6752
rect 33781 6749 33793 6752
rect 33827 6749 33839 6783
rect 33781 6743 33839 6749
rect 35345 6783 35403 6789
rect 35345 6749 35357 6783
rect 35391 6780 35403 6783
rect 35544 6780 35572 6808
rect 35391 6752 35572 6780
rect 36909 6783 36967 6789
rect 35391 6749 35403 6752
rect 35345 6743 35403 6749
rect 36909 6749 36921 6783
rect 36955 6780 36967 6783
rect 36955 6752 37320 6780
rect 36955 6749 36967 6752
rect 36909 6743 36967 6749
rect 37292 6724 37320 6752
rect 38654 6740 38660 6792
rect 38712 6780 38718 6792
rect 38933 6783 38991 6789
rect 38933 6780 38945 6783
rect 38712 6752 38945 6780
rect 38712 6740 38718 6752
rect 38933 6749 38945 6752
rect 38979 6749 38991 6783
rect 38933 6743 38991 6749
rect 25096 6684 29776 6712
rect 29816 6715 29874 6721
rect 25096 6672 25102 6684
rect 29816 6681 29828 6715
rect 29862 6712 29874 6715
rect 30558 6712 30564 6724
rect 29862 6684 30564 6712
rect 29862 6681 29874 6684
rect 29816 6675 29874 6681
rect 30558 6672 30564 6684
rect 30616 6672 30622 6724
rect 31386 6712 31392 6724
rect 31347 6684 31392 6712
rect 31386 6672 31392 6684
rect 31444 6672 31450 6724
rect 31570 6672 31576 6724
rect 31628 6712 31634 6724
rect 31628 6684 31721 6712
rect 31628 6672 31634 6684
rect 32950 6672 32956 6724
rect 33008 6712 33014 6724
rect 33514 6715 33572 6721
rect 33514 6712 33526 6715
rect 33008 6684 33526 6712
rect 33008 6672 33014 6684
rect 33514 6681 33526 6684
rect 33560 6681 33572 6715
rect 33514 6675 33572 6681
rect 35529 6715 35587 6721
rect 35529 6681 35541 6715
rect 35575 6681 35587 6715
rect 35529 6675 35587 6681
rect 16356 6616 18368 6644
rect 16356 6604 16362 6616
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 18564 6616 20637 6644
rect 18564 6604 18570 6616
rect 20625 6613 20637 6616
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 20864 6616 21097 6644
rect 20864 6604 20870 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 27249 6647 27307 6653
rect 27249 6613 27261 6647
rect 27295 6644 27307 6647
rect 27614 6644 27620 6656
rect 27295 6616 27620 6644
rect 27295 6613 27307 6616
rect 27249 6607 27307 6613
rect 27614 6604 27620 6616
rect 27672 6604 27678 6656
rect 30466 6604 30472 6656
rect 30524 6644 30530 6656
rect 31588 6644 31616 6672
rect 30524 6616 31616 6644
rect 31757 6647 31815 6653
rect 30524 6604 30530 6616
rect 31757 6613 31769 6647
rect 31803 6644 31815 6647
rect 31846 6644 31852 6656
rect 31803 6616 31852 6644
rect 31803 6613 31815 6616
rect 31757 6607 31815 6613
rect 31846 6604 31852 6616
rect 31904 6604 31910 6656
rect 32214 6604 32220 6656
rect 32272 6644 32278 6656
rect 35544 6644 35572 6675
rect 36538 6672 36544 6724
rect 36596 6712 36602 6724
rect 37154 6715 37212 6721
rect 37154 6712 37166 6715
rect 36596 6684 37166 6712
rect 36596 6672 36602 6684
rect 37154 6681 37166 6684
rect 37200 6681 37212 6715
rect 37154 6675 37212 6681
rect 37274 6672 37280 6724
rect 37332 6672 37338 6724
rect 38746 6712 38752 6724
rect 38707 6684 38752 6712
rect 38746 6672 38752 6684
rect 38804 6672 38810 6724
rect 38289 6647 38347 6653
rect 38289 6644 38301 6647
rect 32272 6616 38301 6644
rect 32272 6604 32278 6616
rect 38289 6613 38301 6616
rect 38335 6613 38347 6647
rect 38289 6607 38347 6613
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 2133 6443 2191 6449
rect 2133 6409 2145 6443
rect 2179 6440 2191 6443
rect 2222 6440 2228 6452
rect 2179 6412 2228 6440
rect 2179 6409 2191 6412
rect 2133 6403 2191 6409
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3970 6440 3976 6452
rect 2832 6412 3976 6440
rect 2832 6400 2838 6412
rect 3970 6400 3976 6412
rect 4028 6440 4034 6452
rect 4798 6440 4804 6452
rect 4028 6412 4804 6440
rect 4028 6400 4034 6412
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 7745 6443 7803 6449
rect 4908 6412 7696 6440
rect 3234 6332 3240 6384
rect 3292 6372 3298 6384
rect 4908 6372 4936 6412
rect 7558 6372 7564 6384
rect 3292 6344 4936 6372
rect 5828 6344 7564 6372
rect 3292 6332 3298 6344
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 5718 6304 5724 6316
rect 3375 6276 5724 6304
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5828 6313 5856 6344
rect 7558 6332 7564 6344
rect 7616 6332 7622 6384
rect 7668 6372 7696 6412
rect 7745 6409 7757 6443
rect 7791 6440 7803 6443
rect 9306 6440 9312 6452
rect 7791 6412 9312 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 12250 6440 12256 6452
rect 10152 6412 12256 6440
rect 10042 6372 10048 6384
rect 7668 6344 10048 6372
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6621 6307 6679 6313
rect 6621 6304 6633 6307
rect 6328 6276 6633 6304
rect 6328 6264 6334 6276
rect 6621 6273 6633 6276
rect 6667 6273 6679 6307
rect 6621 6267 6679 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 9122 6304 9128 6316
rect 8435 6276 9128 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9674 6304 9680 6316
rect 9635 6276 9680 6304
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 10152 6313 10180 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 14826 6440 14832 6452
rect 14783 6412 14832 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 17770 6400 17776 6452
rect 17828 6440 17834 6452
rect 17865 6443 17923 6449
rect 17865 6440 17877 6443
rect 17828 6412 17877 6440
rect 17828 6400 17834 6412
rect 17865 6409 17877 6412
rect 17911 6409 17923 6443
rect 17865 6403 17923 6409
rect 20898 6400 20904 6452
rect 20956 6400 20962 6452
rect 21358 6400 21364 6452
rect 21416 6440 21422 6452
rect 22005 6443 22063 6449
rect 22005 6440 22017 6443
rect 21416 6412 22017 6440
rect 21416 6400 21422 6412
rect 22005 6409 22017 6412
rect 22051 6409 22063 6443
rect 22005 6403 22063 6409
rect 24946 6400 24952 6452
rect 25004 6440 25010 6452
rect 25593 6443 25651 6449
rect 25593 6440 25605 6443
rect 25004 6412 25605 6440
rect 25004 6400 25010 6412
rect 25593 6409 25605 6412
rect 25639 6440 25651 6443
rect 25682 6440 25688 6452
rect 25639 6412 25688 6440
rect 25639 6409 25651 6412
rect 25593 6403 25651 6409
rect 25682 6400 25688 6412
rect 25740 6400 25746 6452
rect 26237 6443 26295 6449
rect 26237 6409 26249 6443
rect 26283 6440 26295 6443
rect 26878 6440 26884 6452
rect 26283 6412 26884 6440
rect 26283 6409 26295 6412
rect 26237 6403 26295 6409
rect 26878 6400 26884 6412
rect 26936 6400 26942 6452
rect 30558 6440 30564 6452
rect 30519 6412 30564 6440
rect 30558 6400 30564 6412
rect 30616 6400 30622 6452
rect 32306 6400 32312 6452
rect 32364 6440 32370 6452
rect 32950 6440 32956 6452
rect 32364 6412 32444 6440
rect 32911 6412 32956 6440
rect 32364 6400 32370 6412
rect 11882 6372 11888 6384
rect 10336 6344 11888 6372
rect 10336 6313 10364 6344
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 14090 6332 14096 6384
rect 14148 6372 14154 6384
rect 15381 6375 15439 6381
rect 15381 6372 15393 6375
rect 14148 6344 15393 6372
rect 14148 6332 14154 6344
rect 15381 6341 15393 6344
rect 15427 6372 15439 6375
rect 17221 6375 17279 6381
rect 17221 6372 17233 6375
rect 15427 6344 17233 6372
rect 15427 6341 15439 6344
rect 15381 6335 15439 6341
rect 17221 6341 17233 6344
rect 17267 6372 17279 6375
rect 18690 6372 18696 6384
rect 17267 6344 18696 6372
rect 17267 6341 17279 6344
rect 17221 6335 17279 6341
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 20530 6372 20536 6384
rect 18800 6344 20536 6372
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10468 6276 10793 6304
rect 10468 6264 10474 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 11422 6264 11428 6316
rect 11480 6304 11486 6316
rect 12630 6307 12688 6313
rect 12630 6304 12642 6307
rect 11480 6276 12642 6304
rect 11480 6264 11486 6276
rect 12630 6273 12642 6276
rect 12676 6273 12688 6307
rect 12894 6304 12900 6316
rect 12855 6276 12900 6304
rect 12630 6267 12688 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 14550 6304 14556 6316
rect 13771 6276 14556 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 14550 6264 14556 6276
rect 14608 6304 14614 6316
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14608 6276 14933 6304
rect 14608 6264 14614 6276
rect 14921 6273 14933 6276
rect 14967 6304 14979 6307
rect 17589 6307 17647 6313
rect 14967 6276 16436 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 1762 6236 1768 6248
rect 1723 6208 1768 6236
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 3804 6168 3832 6199
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 4120 6208 4169 6236
rect 4120 6196 4126 6208
rect 4157 6205 4169 6208
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 5442 6236 5448 6248
rect 4295 6208 5448 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5684 6208 6377 6236
rect 5684 6196 5690 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 9398 6236 9404 6248
rect 9359 6208 9404 6236
rect 6365 6199 6423 6205
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 9692 6236 9720 6264
rect 13449 6239 13507 6245
rect 9692 6208 11652 6236
rect 4982 6168 4988 6180
rect 3804 6140 4988 6168
rect 4982 6128 4988 6140
rect 5040 6168 5046 6180
rect 5040 6140 5856 6168
rect 5040 6128 5046 6140
rect 4430 6100 4436 6112
rect 4391 6072 4436 6100
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 5718 6100 5724 6112
rect 5675 6072 5724 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5828 6100 5856 6140
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 8076 6140 10977 6168
rect 8076 6128 8082 6140
rect 10965 6137 10977 6140
rect 11011 6168 11023 6171
rect 11054 6168 11060 6180
rect 11011 6140 11060 6168
rect 11011 6137 11023 6140
rect 10965 6131 11023 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 6730 6100 6736 6112
rect 5828 6072 6736 6100
rect 6730 6060 6736 6072
rect 6788 6100 6794 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 6788 6072 8217 6100
rect 6788 6060 6794 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8205 6063 8263 6069
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 10226 6100 10232 6112
rect 8352 6072 10232 6100
rect 8352 6060 8358 6072
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6100 10379 6103
rect 10410 6100 10416 6112
rect 10367 6072 10416 6100
rect 10367 6069 10379 6072
rect 10321 6063 10379 6069
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11204 6072 11529 6100
rect 11204 6060 11210 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11624 6100 11652 6208
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 11974 6100 11980 6112
rect 11624 6072 11980 6100
rect 11517 6063 11575 6069
rect 11974 6060 11980 6072
rect 12032 6100 12038 6112
rect 13464 6100 13492 6199
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 15013 6239 15071 6245
rect 15013 6236 15025 6239
rect 13872 6208 15025 6236
rect 13872 6196 13878 6208
rect 15013 6205 15025 6208
rect 15059 6205 15071 6239
rect 16408 6236 16436 6276
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 17862 6304 17868 6316
rect 17635 6276 17868 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 17862 6264 17868 6276
rect 17920 6264 17926 6316
rect 17678 6236 17684 6248
rect 16408 6208 17684 6236
rect 15013 6199 15071 6205
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18800 6236 18828 6344
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 20804 6316 20862 6319
rect 20254 6264 20260 6316
rect 20312 6304 20318 6316
rect 20625 6307 20683 6313
rect 20804 6310 20812 6316
rect 20625 6304 20637 6307
rect 20312 6276 20637 6304
rect 20312 6264 20318 6276
rect 20625 6273 20637 6276
rect 20671 6273 20683 6307
rect 20773 6282 20812 6310
rect 20804 6273 20812 6282
rect 20625 6267 20683 6273
rect 20806 6264 20812 6273
rect 20864 6264 20870 6316
rect 20916 6313 20944 6400
rect 21269 6375 21327 6381
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 23118 6375 23176 6381
rect 23118 6372 23130 6375
rect 21315 6344 23130 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 23118 6341 23130 6344
rect 23164 6341 23176 6375
rect 23118 6335 23176 6341
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 20990 6264 20996 6316
rect 21048 6304 21054 6316
rect 23385 6307 23443 6313
rect 21048 6276 21093 6304
rect 21048 6264 21054 6276
rect 23385 6273 23397 6307
rect 23431 6304 23443 6307
rect 23474 6304 23480 6316
rect 23431 6276 23480 6304
rect 23431 6273 23443 6276
rect 23385 6267 23443 6273
rect 23474 6264 23480 6276
rect 23532 6264 23538 6316
rect 24486 6313 24492 6316
rect 24480 6267 24492 6313
rect 24544 6304 24550 6316
rect 24544 6276 24580 6304
rect 24486 6264 24492 6267
rect 24544 6264 24550 6276
rect 25406 6264 25412 6316
rect 25464 6304 25470 6316
rect 26145 6307 26203 6313
rect 26145 6304 26157 6307
rect 25464 6276 26157 6304
rect 25464 6264 25470 6276
rect 26145 6273 26157 6276
rect 26191 6273 26203 6307
rect 26145 6267 26203 6273
rect 20070 6236 20076 6248
rect 17828 6208 18828 6236
rect 20031 6208 20076 6236
rect 17828 6196 17834 6208
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 24210 6236 24216 6248
rect 24171 6208 24216 6236
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 26160 6236 26188 6267
rect 26326 6264 26332 6316
rect 26384 6304 26390 6316
rect 27982 6304 27988 6316
rect 26384 6276 27988 6304
rect 26384 6264 26390 6276
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 30374 6264 30380 6316
rect 30432 6304 30438 6316
rect 30834 6304 30840 6316
rect 30432 6276 30840 6304
rect 30432 6264 30438 6276
rect 30834 6264 30840 6276
rect 30892 6264 30898 6316
rect 30929 6307 30987 6313
rect 30929 6273 30941 6307
rect 30975 6273 30987 6307
rect 30929 6267 30987 6273
rect 26973 6239 27031 6245
rect 26973 6236 26985 6239
rect 26160 6208 26985 6236
rect 26973 6205 26985 6208
rect 27019 6205 27031 6239
rect 26973 6199 27031 6205
rect 17586 6128 17592 6180
rect 17644 6168 17650 6180
rect 20254 6168 20260 6180
rect 17644 6140 20260 6168
rect 17644 6128 17650 6140
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 28626 6128 28632 6180
rect 28684 6168 28690 6180
rect 29273 6171 29331 6177
rect 29273 6168 29285 6171
rect 28684 6140 29285 6168
rect 28684 6128 28690 6140
rect 29273 6137 29285 6140
rect 29319 6137 29331 6171
rect 29273 6131 29331 6137
rect 12032 6072 13492 6100
rect 16117 6103 16175 6109
rect 12032 6060 12038 6072
rect 16117 6069 16129 6103
rect 16163 6100 16175 6103
rect 16482 6100 16488 6112
rect 16163 6072 16488 6100
rect 16163 6069 16175 6072
rect 16117 6063 16175 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 16761 6103 16819 6109
rect 16761 6069 16773 6103
rect 16807 6100 16819 6103
rect 17494 6100 17500 6112
rect 16807 6072 17500 6100
rect 16807 6069 16819 6072
rect 16761 6063 16819 6069
rect 17494 6060 17500 6072
rect 17552 6100 17558 6112
rect 17770 6100 17776 6112
rect 17552 6072 17776 6100
rect 17552 6060 17558 6072
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 18693 6103 18751 6109
rect 18693 6100 18705 6103
rect 18656 6072 18705 6100
rect 18656 6060 18662 6072
rect 18693 6069 18705 6072
rect 18739 6069 18751 6103
rect 18693 6063 18751 6069
rect 19337 6103 19395 6109
rect 19337 6069 19349 6103
rect 19383 6100 19395 6103
rect 19426 6100 19432 6112
rect 19383 6072 19432 6100
rect 19383 6069 19395 6072
rect 19337 6063 19395 6069
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 30944 6100 30972 6267
rect 31018 6264 31024 6316
rect 31076 6304 31082 6316
rect 31205 6307 31263 6313
rect 31076 6276 31121 6304
rect 31076 6264 31082 6276
rect 31205 6273 31217 6307
rect 31251 6304 31263 6307
rect 32309 6307 32367 6313
rect 32309 6304 32321 6307
rect 31251 6276 32321 6304
rect 31251 6273 31263 6276
rect 31205 6267 31263 6273
rect 32309 6273 32321 6276
rect 32355 6273 32367 6307
rect 32416 6304 32444 6412
rect 32950 6400 32956 6412
rect 33008 6400 33014 6452
rect 32766 6372 32772 6384
rect 32600 6344 32772 6372
rect 32600 6313 32628 6344
rect 32766 6332 32772 6344
rect 32824 6332 32830 6384
rect 33226 6332 33232 6384
rect 33284 6372 33290 6384
rect 33689 6375 33747 6381
rect 33689 6372 33701 6375
rect 33284 6344 33701 6372
rect 33284 6332 33290 6344
rect 33689 6341 33701 6344
rect 33735 6341 33747 6375
rect 33689 6335 33747 6341
rect 32488 6307 32546 6313
rect 32488 6304 32500 6307
rect 32416 6276 32500 6304
rect 32309 6267 32367 6273
rect 32488 6273 32500 6276
rect 32534 6273 32546 6307
rect 32488 6267 32546 6273
rect 32585 6307 32643 6313
rect 32585 6273 32597 6307
rect 32631 6273 32643 6307
rect 32585 6267 32643 6273
rect 32324 6236 32352 6267
rect 32674 6264 32680 6316
rect 32732 6304 32738 6316
rect 33502 6304 33508 6316
rect 32732 6276 33180 6304
rect 33463 6276 33508 6304
rect 32732 6264 32738 6276
rect 33152 6236 33180 6276
rect 33502 6264 33508 6276
rect 33560 6264 33566 6316
rect 35483 6307 35541 6313
rect 35483 6304 35495 6307
rect 34716 6276 35495 6304
rect 34716 6245 34744 6276
rect 35483 6273 35495 6276
rect 35529 6273 35541 6307
rect 35618 6304 35624 6316
rect 35579 6276 35624 6304
rect 35483 6267 35541 6273
rect 35618 6264 35624 6276
rect 35676 6264 35682 6316
rect 35734 6307 35792 6313
rect 35734 6273 35746 6307
rect 35780 6304 35792 6307
rect 35897 6307 35955 6313
rect 35780 6276 35857 6304
rect 35780 6273 35792 6276
rect 35734 6267 35792 6273
rect 34701 6239 34759 6245
rect 34701 6236 34713 6239
rect 32324 6208 32444 6236
rect 33152 6208 34713 6236
rect 32416 6168 32444 6208
rect 34701 6205 34713 6208
rect 34747 6205 34759 6239
rect 35829 6236 35857 6276
rect 35897 6273 35909 6307
rect 35943 6304 35955 6307
rect 35986 6304 35992 6316
rect 35943 6276 35992 6304
rect 35943 6273 35955 6276
rect 35897 6267 35955 6273
rect 35986 6264 35992 6276
rect 36044 6304 36050 6316
rect 39022 6304 39028 6316
rect 36044 6276 39028 6304
rect 36044 6264 36050 6276
rect 39022 6264 39028 6276
rect 39080 6264 39086 6316
rect 37182 6236 37188 6248
rect 35829 6208 37188 6236
rect 34701 6199 34759 6205
rect 37182 6196 37188 6208
rect 37240 6196 37246 6248
rect 33134 6168 33140 6180
rect 32416 6140 33140 6168
rect 33134 6128 33140 6140
rect 33192 6168 33198 6180
rect 34054 6168 34060 6180
rect 33192 6140 34060 6168
rect 33192 6128 33198 6140
rect 34054 6128 34060 6140
rect 34112 6128 34118 6180
rect 67634 6168 67640 6180
rect 67595 6140 67640 6168
rect 67634 6128 67640 6140
rect 67692 6128 67698 6180
rect 31662 6100 31668 6112
rect 30944 6072 31668 6100
rect 31662 6060 31668 6072
rect 31720 6100 31726 6112
rect 32766 6100 32772 6112
rect 31720 6072 32772 6100
rect 31720 6060 31726 6072
rect 32766 6060 32772 6072
rect 32824 6060 32830 6112
rect 33873 6103 33931 6109
rect 33873 6069 33885 6103
rect 33919 6100 33931 6103
rect 34606 6100 34612 6112
rect 33919 6072 34612 6100
rect 33919 6069 33931 6072
rect 33873 6063 33931 6069
rect 34606 6060 34612 6072
rect 34664 6060 34670 6112
rect 35253 6103 35311 6109
rect 35253 6069 35265 6103
rect 35299 6100 35311 6103
rect 35526 6100 35532 6112
rect 35299 6072 35532 6100
rect 35299 6069 35311 6072
rect 35253 6063 35311 6069
rect 35526 6060 35532 6072
rect 35584 6060 35590 6112
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 4890 5896 4896 5908
rect 1627 5868 4896 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 6270 5896 6276 5908
rect 6231 5868 6276 5896
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 8110 5896 8116 5908
rect 7423 5868 8116 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 12069 5899 12127 5905
rect 12069 5865 12081 5899
rect 12115 5896 12127 5899
rect 13722 5896 13728 5908
rect 12115 5868 13728 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 15194 5896 15200 5908
rect 14783 5868 15200 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15194 5856 15200 5868
rect 15252 5856 15258 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18049 5899 18107 5905
rect 18049 5896 18061 5899
rect 18012 5868 18061 5896
rect 18012 5856 18018 5868
rect 18049 5865 18061 5868
rect 18095 5865 18107 5899
rect 18049 5859 18107 5865
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 18288 5868 19257 5896
rect 18288 5856 18294 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 22281 5899 22339 5905
rect 22281 5896 22293 5899
rect 19245 5859 19303 5865
rect 21744 5868 22293 5896
rect 5442 5788 5448 5840
rect 5500 5828 5506 5840
rect 5500 5800 7236 5828
rect 5500 5788 5506 5800
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2314 5760 2320 5772
rect 1912 5732 2320 5760
rect 1912 5720 1918 5732
rect 2314 5720 2320 5732
rect 2372 5760 2378 5772
rect 2593 5763 2651 5769
rect 2593 5760 2605 5763
rect 2372 5732 2605 5760
rect 2372 5720 2378 5732
rect 2593 5729 2605 5732
rect 2639 5729 2651 5763
rect 6730 5760 6736 5772
rect 6691 5732 6736 5760
rect 2593 5723 2651 5729
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7208 5769 7236 5800
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 8294 5828 8300 5840
rect 7984 5800 8300 5828
rect 7984 5788 7990 5800
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 10928 5800 10977 5828
rect 10928 5788 10934 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 10965 5791 11023 5797
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 12526 5828 12532 5840
rect 11112 5800 12532 5828
rect 11112 5788 11118 5800
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 12710 5828 12716 5840
rect 12671 5800 12716 5828
rect 12710 5788 12716 5800
rect 12768 5828 12774 5840
rect 13538 5828 13544 5840
rect 12768 5800 13544 5828
rect 12768 5788 12774 5800
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 18322 5828 18328 5840
rect 15028 5800 18328 5828
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 9398 5760 9404 5772
rect 7239 5732 9404 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 10410 5760 10416 5772
rect 10371 5732 10416 5760
rect 10410 5720 10416 5732
rect 10468 5760 10474 5772
rect 11514 5760 11520 5772
rect 10468 5732 11520 5760
rect 10468 5720 10474 5732
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 12406 5732 14473 5760
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 3200 5664 5181 5692
rect 3200 5652 3206 5664
rect 5169 5661 5181 5664
rect 5215 5692 5227 5695
rect 5626 5692 5632 5704
rect 5215 5664 5632 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 7098 5692 7104 5704
rect 7059 5664 7104 5692
rect 6089 5655 6147 5661
rect 2409 5627 2467 5633
rect 2409 5593 2421 5627
rect 2455 5624 2467 5627
rect 2774 5624 2780 5636
rect 2455 5596 2780 5624
rect 2455 5593 2467 5596
rect 2409 5587 2467 5593
rect 2774 5584 2780 5596
rect 2832 5584 2838 5636
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4902 5627 4960 5633
rect 4902 5624 4914 5627
rect 4212 5596 4914 5624
rect 4212 5584 4218 5596
rect 4902 5593 4914 5596
rect 4948 5593 4960 5627
rect 6104 5624 6132 5655
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8294 5692 8300 5704
rect 8255 5664 8300 5692
rect 8113 5655 8171 5661
rect 7929 5627 7987 5633
rect 7929 5624 7941 5627
rect 6104 5596 7941 5624
rect 4902 5587 4960 5593
rect 7929 5593 7941 5596
rect 7975 5593 7987 5627
rect 8128 5624 8156 5655
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8938 5692 8944 5704
rect 8899 5664 8944 5692
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 9048 5664 9229 5692
rect 8662 5624 8668 5636
rect 8128 5596 8668 5624
rect 7929 5587 7987 5593
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 2004 5528 2053 5556
rect 2004 5516 2010 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 2547 5528 3801 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 3789 5525 3801 5528
rect 3835 5556 3847 5559
rect 4062 5556 4068 5568
rect 3835 5528 4068 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 7006 5556 7012 5568
rect 5224 5528 7012 5556
rect 5224 5516 5230 5528
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 9048 5556 9076 5664
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 12406 5692 12434 5732
rect 14461 5729 14473 5732
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 14608 5732 14653 5760
rect 14608 5720 14614 5732
rect 9364 5664 12434 5692
rect 12805 5695 12863 5701
rect 9364 5652 9370 5664
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 13262 5692 13268 5704
rect 12851 5664 13268 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5661 13599 5695
rect 14090 5692 14096 5704
rect 14051 5664 14096 5692
rect 13541 5655 13599 5661
rect 9122 5584 9128 5636
rect 9180 5624 9186 5636
rect 10229 5627 10287 5633
rect 10229 5624 10241 5627
rect 9180 5596 10241 5624
rect 9180 5584 9186 5596
rect 10229 5593 10241 5596
rect 10275 5624 10287 5627
rect 10965 5627 11023 5633
rect 10275 5596 10824 5624
rect 10275 5593 10287 5596
rect 10229 5587 10287 5593
rect 8352 5528 9076 5556
rect 10505 5559 10563 5565
rect 8352 5516 8358 5528
rect 10505 5525 10517 5559
rect 10551 5556 10563 5559
rect 10686 5556 10692 5568
rect 10551 5528 10692 5556
rect 10551 5525 10563 5528
rect 10505 5519 10563 5525
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10796 5556 10824 5596
rect 10965 5593 10977 5627
rect 11011 5624 11023 5627
rect 11606 5624 11612 5636
rect 11011 5596 11612 5624
rect 11011 5593 11023 5596
rect 10965 5587 11023 5593
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 12066 5584 12072 5636
rect 12124 5624 12130 5636
rect 12529 5627 12587 5633
rect 12529 5624 12541 5627
rect 12124 5596 12541 5624
rect 12124 5584 12130 5596
rect 12529 5593 12541 5596
rect 12575 5593 12587 5627
rect 13170 5624 13176 5636
rect 12529 5587 12587 5593
rect 12636 5596 13176 5624
rect 12636 5556 12664 5596
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 13556 5624 13584 5655
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 15028 5624 15056 5800
rect 18322 5788 18328 5800
rect 18380 5788 18386 5840
rect 19150 5788 19156 5840
rect 19208 5828 19214 5840
rect 21744 5828 21772 5868
rect 22281 5865 22293 5868
rect 22327 5896 22339 5899
rect 23658 5896 23664 5908
rect 22327 5868 23664 5896
rect 22327 5865 22339 5868
rect 22281 5859 22339 5865
rect 23658 5856 23664 5868
rect 23716 5856 23722 5908
rect 24397 5899 24455 5905
rect 24397 5865 24409 5899
rect 24443 5896 24455 5899
rect 24486 5896 24492 5908
rect 24443 5868 24492 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 26326 5896 26332 5908
rect 26287 5868 26332 5896
rect 26326 5856 26332 5868
rect 26384 5856 26390 5908
rect 26694 5856 26700 5908
rect 26752 5896 26758 5908
rect 26881 5899 26939 5905
rect 26881 5896 26893 5899
rect 26752 5868 26893 5896
rect 26752 5856 26758 5868
rect 26881 5865 26893 5868
rect 26927 5896 26939 5899
rect 27338 5896 27344 5908
rect 26927 5868 27344 5896
rect 26927 5865 26939 5868
rect 26881 5859 26939 5865
rect 27338 5856 27344 5868
rect 27396 5856 27402 5908
rect 27525 5899 27583 5905
rect 27525 5865 27537 5899
rect 27571 5896 27583 5899
rect 27890 5896 27896 5908
rect 27571 5868 27896 5896
rect 27571 5865 27583 5868
rect 27525 5859 27583 5865
rect 27890 5856 27896 5868
rect 27948 5856 27954 5908
rect 29454 5856 29460 5908
rect 29512 5896 29518 5908
rect 29549 5899 29607 5905
rect 29549 5896 29561 5899
rect 29512 5868 29561 5896
rect 29512 5856 29518 5868
rect 29549 5865 29561 5868
rect 29595 5865 29607 5899
rect 29549 5859 29607 5865
rect 30742 5856 30748 5908
rect 30800 5896 30806 5908
rect 32953 5899 33011 5905
rect 32953 5896 32965 5899
rect 30800 5868 32965 5896
rect 30800 5856 30806 5868
rect 19208 5800 21772 5828
rect 19208 5788 19214 5800
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 16485 5763 16543 5769
rect 16485 5760 16497 5763
rect 15335 5732 16497 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 16485 5729 16497 5732
rect 16531 5760 16543 5763
rect 17126 5760 17132 5772
rect 16531 5732 17132 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 17678 5720 17684 5772
rect 17736 5760 17742 5772
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 17736 5732 18245 5760
rect 17736 5720 17742 5732
rect 18233 5729 18245 5732
rect 18279 5760 18291 5763
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 18279 5732 19441 5760
rect 18279 5729 18291 5732
rect 18233 5723 18291 5729
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 19521 5763 19579 5769
rect 19521 5729 19533 5763
rect 19567 5760 19579 5763
rect 20070 5760 20076 5772
rect 19567 5732 20076 5760
rect 19567 5729 19579 5732
rect 19521 5723 19579 5729
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 20364 5769 20392 5800
rect 24210 5788 24216 5840
rect 24268 5828 24274 5840
rect 28350 5828 28356 5840
rect 24268 5800 28356 5828
rect 24268 5788 24274 5800
rect 28350 5788 28356 5800
rect 28408 5828 28414 5840
rect 28626 5828 28632 5840
rect 28408 5800 28632 5828
rect 28408 5788 28414 5800
rect 28626 5788 28632 5800
rect 28684 5788 28690 5840
rect 20349 5763 20407 5769
rect 20349 5729 20361 5763
rect 20395 5729 20407 5763
rect 20349 5723 20407 5729
rect 20898 5720 20904 5772
rect 20956 5760 20962 5772
rect 22925 5763 22983 5769
rect 22925 5760 22937 5763
rect 20956 5732 22937 5760
rect 20956 5720 20962 5732
rect 22925 5729 22937 5732
rect 22971 5729 22983 5763
rect 22925 5723 22983 5729
rect 23201 5763 23259 5769
rect 23201 5729 23213 5763
rect 23247 5760 23259 5763
rect 25590 5760 25596 5772
rect 23247 5732 25596 5760
rect 23247 5729 23259 5732
rect 23201 5723 23259 5729
rect 15194 5692 15200 5704
rect 15155 5664 15200 5692
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15378 5692 15384 5704
rect 15339 5664 15384 5692
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5692 17647 5695
rect 18046 5692 18052 5704
rect 17635 5664 18052 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5692 18383 5695
rect 19334 5692 19340 5704
rect 18371 5664 19340 5692
rect 18371 5661 18383 5664
rect 18325 5655 18383 5661
rect 19306 5660 19340 5664
rect 19334 5652 19340 5660
rect 19392 5652 19398 5704
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5661 20683 5695
rect 21634 5692 21640 5704
rect 21595 5664 21640 5692
rect 20625 5655 20683 5661
rect 13556 5596 15056 5624
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 16117 5627 16175 5633
rect 16117 5624 16129 5627
rect 15344 5596 16129 5624
rect 15344 5584 15350 5596
rect 16117 5593 16129 5596
rect 16163 5624 16175 5627
rect 16298 5624 16304 5636
rect 16163 5596 16304 5624
rect 16163 5593 16175 5596
rect 16117 5587 16175 5593
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 16577 5627 16635 5633
rect 16577 5593 16589 5627
rect 16623 5624 16635 5627
rect 16850 5624 16856 5636
rect 16623 5596 16856 5624
rect 16623 5593 16635 5596
rect 16577 5587 16635 5593
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 18690 5624 18696 5636
rect 18651 5596 18696 5624
rect 18690 5584 18696 5596
rect 18748 5624 18754 5636
rect 19889 5627 19947 5633
rect 19889 5624 19901 5627
rect 18748 5596 19901 5624
rect 18748 5584 18754 5596
rect 19889 5593 19901 5596
rect 19935 5593 19947 5627
rect 19889 5587 19947 5593
rect 20254 5584 20260 5636
rect 20312 5624 20318 5636
rect 20640 5624 20668 5655
rect 21634 5652 21640 5664
rect 21692 5652 21698 5704
rect 24578 5652 24584 5704
rect 24636 5701 24642 5704
rect 24780 5701 24808 5732
rect 25590 5720 25596 5732
rect 25648 5720 25654 5772
rect 27890 5720 27896 5772
rect 27948 5760 27954 5772
rect 30926 5760 30932 5772
rect 27948 5732 28396 5760
rect 30887 5732 30932 5760
rect 27948 5720 27954 5732
rect 24636 5695 24685 5701
rect 24636 5661 24639 5695
rect 24673 5661 24685 5695
rect 24636 5655 24685 5661
rect 24765 5695 24823 5701
rect 24765 5661 24777 5695
rect 24811 5661 24823 5695
rect 24765 5655 24823 5661
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5668 24915 5695
rect 25041 5695 25099 5701
rect 24903 5661 24992 5668
rect 24857 5655 24992 5661
rect 25041 5661 25053 5695
rect 25087 5692 25099 5695
rect 25130 5692 25136 5704
rect 25087 5664 25136 5692
rect 25087 5661 25099 5664
rect 25041 5655 25099 5661
rect 24636 5652 24642 5655
rect 24872 5640 24992 5655
rect 25130 5652 25136 5664
rect 25188 5652 25194 5704
rect 25682 5692 25688 5704
rect 25643 5664 25688 5692
rect 25682 5652 25688 5664
rect 25740 5652 25746 5704
rect 28166 5701 28172 5704
rect 27985 5695 28043 5701
rect 27985 5692 27997 5695
rect 27908 5664 27997 5692
rect 20312 5596 20668 5624
rect 24964 5624 24992 5640
rect 27908 5636 27936 5664
rect 27985 5661 27997 5664
rect 28031 5661 28043 5695
rect 28164 5692 28172 5701
rect 28127 5664 28172 5692
rect 27985 5655 28043 5661
rect 28164 5655 28172 5664
rect 28166 5652 28172 5655
rect 28224 5652 28230 5704
rect 28368 5701 28396 5732
rect 30926 5720 30932 5732
rect 30984 5720 30990 5772
rect 28353 5695 28411 5701
rect 28264 5689 28322 5695
rect 28264 5655 28276 5689
rect 28310 5655 28322 5689
rect 28353 5661 28365 5695
rect 28399 5661 28411 5695
rect 28353 5655 28411 5661
rect 31588 5686 31616 5868
rect 32953 5865 32965 5868
rect 32999 5896 33011 5899
rect 32999 5868 33824 5896
rect 32999 5865 33011 5868
rect 32953 5859 33011 5865
rect 31665 5695 31723 5701
rect 31665 5686 31677 5695
rect 31588 5661 31677 5686
rect 31711 5661 31723 5695
rect 31588 5658 31723 5661
rect 31665 5655 31723 5658
rect 31754 5692 31812 5698
rect 31754 5658 31766 5692
rect 31800 5658 31812 5692
rect 28264 5649 28322 5655
rect 31754 5652 31812 5658
rect 31846 5652 31852 5704
rect 31904 5701 31910 5704
rect 31904 5692 31912 5701
rect 32033 5695 32091 5701
rect 31904 5664 31949 5692
rect 31904 5655 31912 5664
rect 32033 5661 32045 5695
rect 32079 5692 32091 5695
rect 33134 5692 33140 5704
rect 32079 5664 33140 5692
rect 32079 5661 32091 5664
rect 32033 5655 32091 5661
rect 31904 5652 31910 5655
rect 33134 5652 33140 5664
rect 33192 5652 33198 5704
rect 33796 5701 33824 5868
rect 38654 5856 38660 5908
rect 38712 5896 38718 5908
rect 38749 5899 38807 5905
rect 38749 5896 38761 5899
rect 38712 5868 38761 5896
rect 38712 5856 38718 5868
rect 38749 5865 38761 5868
rect 38795 5865 38807 5899
rect 38749 5859 38807 5865
rect 35618 5760 35624 5772
rect 33888 5732 35624 5760
rect 33888 5701 33916 5732
rect 35618 5720 35624 5732
rect 35676 5720 35682 5772
rect 33781 5695 33839 5701
rect 33781 5661 33793 5695
rect 33827 5661 33839 5695
rect 33781 5655 33839 5661
rect 33873 5695 33931 5701
rect 33873 5661 33885 5695
rect 33919 5661 33931 5695
rect 33873 5655 33931 5661
rect 33965 5695 34023 5701
rect 33965 5661 33977 5695
rect 34011 5692 34023 5695
rect 34054 5692 34060 5704
rect 34011 5664 34060 5692
rect 34011 5661 34023 5664
rect 33965 5655 34023 5661
rect 34054 5652 34060 5664
rect 34112 5652 34118 5704
rect 34149 5695 34207 5701
rect 34149 5661 34161 5695
rect 34195 5692 34207 5695
rect 34238 5692 34244 5704
rect 34195 5664 34244 5692
rect 34195 5661 34207 5664
rect 34149 5655 34207 5661
rect 34238 5652 34244 5664
rect 34296 5652 34302 5704
rect 37369 5695 37427 5701
rect 37369 5692 37381 5695
rect 37292 5664 37381 5692
rect 25501 5627 25559 5633
rect 25501 5624 25513 5627
rect 24964 5596 25513 5624
rect 20312 5584 20318 5596
rect 25501 5593 25513 5596
rect 25547 5593 25559 5627
rect 25866 5624 25872 5636
rect 25827 5596 25872 5624
rect 25501 5587 25559 5593
rect 25866 5584 25872 5596
rect 25924 5584 25930 5636
rect 26970 5584 26976 5636
rect 27028 5624 27034 5636
rect 27890 5624 27896 5636
rect 27028 5596 27896 5624
rect 27028 5584 27034 5596
rect 27890 5584 27896 5596
rect 27948 5584 27954 5636
rect 28276 5568 28304 5649
rect 28629 5627 28687 5633
rect 28629 5593 28641 5627
rect 28675 5624 28687 5627
rect 30662 5627 30720 5633
rect 30662 5624 30674 5627
rect 28675 5596 30674 5624
rect 28675 5593 28687 5596
rect 28629 5587 28687 5593
rect 30662 5593 30674 5596
rect 30708 5593 30720 5627
rect 31772 5624 31800 5652
rect 37292 5636 37320 5664
rect 37369 5661 37381 5664
rect 37415 5661 37427 5695
rect 37369 5655 37427 5661
rect 37636 5695 37694 5701
rect 37636 5661 37648 5695
rect 37682 5692 37694 5695
rect 38378 5692 38384 5704
rect 37682 5664 38384 5692
rect 37682 5661 37694 5664
rect 37636 5655 37694 5661
rect 38378 5652 38384 5664
rect 38436 5652 38442 5704
rect 35066 5624 35072 5636
rect 30662 5587 30720 5593
rect 31680 5596 31800 5624
rect 35027 5596 35072 5624
rect 31680 5568 31708 5596
rect 35066 5584 35072 5596
rect 35124 5624 35130 5636
rect 35342 5624 35348 5636
rect 35124 5596 35348 5624
rect 35124 5584 35130 5596
rect 35342 5584 35348 5596
rect 35400 5584 35406 5636
rect 36817 5627 36875 5633
rect 36817 5593 36829 5627
rect 36863 5624 36875 5627
rect 37274 5624 37280 5636
rect 36863 5596 37280 5624
rect 36863 5593 36875 5596
rect 36817 5587 36875 5593
rect 37274 5584 37280 5596
rect 37332 5584 37338 5636
rect 12802 5556 12808 5568
rect 10796 5528 12664 5556
rect 12763 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 16666 5556 16672 5568
rect 16439 5528 16672 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 16761 5559 16819 5565
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 19978 5556 19984 5568
rect 16807 5528 19984 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 20070 5516 20076 5568
rect 20128 5556 20134 5568
rect 20806 5556 20812 5568
rect 20128 5528 20812 5556
rect 20128 5516 20134 5528
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 21821 5559 21879 5565
rect 21821 5525 21833 5559
rect 21867 5556 21879 5559
rect 23014 5556 23020 5568
rect 21867 5528 23020 5556
rect 21867 5525 21879 5528
rect 21821 5519 21879 5525
rect 23014 5516 23020 5528
rect 23072 5516 23078 5568
rect 27246 5516 27252 5568
rect 27304 5556 27310 5568
rect 28258 5556 28264 5568
rect 27304 5528 28264 5556
rect 27304 5516 27310 5528
rect 28258 5516 28264 5528
rect 28316 5516 28322 5568
rect 31294 5516 31300 5568
rect 31352 5556 31358 5568
rect 31389 5559 31447 5565
rect 31389 5556 31401 5559
rect 31352 5528 31401 5556
rect 31352 5516 31358 5528
rect 31389 5525 31401 5528
rect 31435 5525 31447 5559
rect 31389 5519 31447 5525
rect 31662 5516 31668 5568
rect 31720 5516 31726 5568
rect 33505 5559 33563 5565
rect 33505 5525 33517 5559
rect 33551 5556 33563 5559
rect 34514 5556 34520 5568
rect 33551 5528 34520 5556
rect 33551 5525 33563 5528
rect 33505 5519 33563 5525
rect 34514 5516 34520 5528
rect 34572 5516 34578 5568
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 4154 5352 4160 5364
rect 2823 5324 4160 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4982 5352 4988 5364
rect 4479 5324 4988 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5534 5352 5540 5364
rect 5123 5324 5540 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 7469 5355 7527 5361
rect 7469 5321 7481 5355
rect 7515 5321 7527 5355
rect 8662 5352 8668 5364
rect 8623 5324 8668 5352
rect 7469 5315 7527 5321
rect 7484 5284 7512 5315
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9030 5352 9036 5364
rect 8991 5324 9036 5352
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9306 5352 9312 5364
rect 9171 5324 9312 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 10965 5355 11023 5361
rect 10965 5321 10977 5355
rect 11011 5352 11023 5355
rect 14918 5352 14924 5364
rect 11011 5324 14924 5352
rect 11011 5321 11023 5324
rect 10965 5315 11023 5321
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15010 5312 15016 5364
rect 15068 5352 15074 5364
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 15068 5324 15117 5352
rect 15068 5312 15074 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15105 5315 15163 5321
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 16945 5355 17003 5361
rect 16945 5352 16957 5355
rect 16356 5324 16957 5352
rect 16356 5312 16362 5324
rect 16945 5321 16957 5324
rect 16991 5321 17003 5355
rect 16945 5315 17003 5321
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 19392 5324 20729 5352
rect 19392 5312 19398 5324
rect 20717 5321 20729 5324
rect 20763 5352 20775 5355
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 20763 5324 21833 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 23014 5312 23020 5364
rect 23072 5352 23078 5364
rect 23072 5324 24716 5352
rect 23072 5312 23078 5324
rect 10870 5284 10876 5296
rect 7484 5256 10876 5284
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 11514 5284 11520 5296
rect 11475 5256 11520 5284
rect 11514 5244 11520 5256
rect 11572 5244 11578 5296
rect 11606 5244 11612 5296
rect 11664 5284 11670 5296
rect 12342 5284 12348 5296
rect 11664 5256 12348 5284
rect 11664 5244 11670 5256
rect 12342 5244 12348 5256
rect 12400 5244 12406 5296
rect 13538 5244 13544 5296
rect 13596 5284 13602 5296
rect 15378 5284 15384 5296
rect 13596 5256 15384 5284
rect 13596 5244 13602 5256
rect 1762 5216 1768 5228
rect 1723 5188 1768 5216
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2179 5188 2605 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5442 5216 5448 5228
rect 4939 5188 5448 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 5810 5216 5816 5228
rect 5675 5188 5816 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 5810 5176 5816 5188
rect 5868 5216 5874 5228
rect 6362 5216 6368 5228
rect 5868 5188 6368 5216
rect 5868 5176 5874 5188
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 6638 5216 6644 5228
rect 6599 5188 6644 5216
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 8018 5216 8024 5228
rect 7331 5188 8024 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 9766 5216 9772 5228
rect 8168 5188 9772 5216
rect 8168 5176 8174 5188
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 10134 5216 10140 5228
rect 10095 5188 10140 5216
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10888 5216 10916 5244
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 10888 5188 11989 5216
rect 10781 5179 10839 5185
rect 11977 5185 11989 5188
rect 12023 5216 12035 5219
rect 12894 5216 12900 5228
rect 12023 5188 12900 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 4798 5148 4804 5160
rect 4759 5120 4804 5148
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 9306 5148 9312 5160
rect 6748 5120 9168 5148
rect 9267 5120 9312 5148
rect 3973 5083 4031 5089
rect 3973 5049 3985 5083
rect 4019 5080 4031 5083
rect 6748 5080 6776 5120
rect 4019 5052 6776 5080
rect 6825 5083 6883 5089
rect 4019 5049 4031 5052
rect 3973 5043 4031 5049
rect 6825 5049 6837 5083
rect 6871 5080 6883 5083
rect 8846 5080 8852 5092
rect 6871 5052 8852 5080
rect 6871 5049 6883 5052
rect 6825 5043 6883 5049
rect 8846 5040 8852 5052
rect 8904 5040 8910 5092
rect 3418 5012 3424 5024
rect 3379 4984 3424 5012
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 7374 5012 7380 5024
rect 5859 4984 7380 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7524 4984 8033 5012
rect 7524 4972 7530 4984
rect 8021 4981 8033 4984
rect 8067 5012 8079 5015
rect 8938 5012 8944 5024
rect 8067 4984 8944 5012
rect 8067 4981 8079 4984
rect 8021 4975 8079 4981
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 9140 5012 9168 5120
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10796 5148 10824 5179
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13262 5216 13268 5228
rect 13223 5188 13268 5216
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 14660 5225 14688 5256
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 17126 5284 17132 5296
rect 17087 5256 17132 5284
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 17405 5287 17463 5293
rect 17405 5253 17417 5287
rect 17451 5284 17463 5287
rect 20438 5284 20444 5296
rect 17451 5256 20444 5284
rect 17451 5253 17463 5256
rect 17405 5247 17463 5253
rect 20438 5244 20444 5256
rect 20496 5244 20502 5296
rect 24688 5284 24716 5324
rect 24762 5312 24768 5364
rect 24820 5352 24826 5364
rect 24949 5355 25007 5361
rect 24949 5352 24961 5355
rect 24820 5324 24961 5352
rect 24820 5312 24826 5324
rect 24949 5321 24961 5324
rect 24995 5321 25007 5355
rect 24949 5315 25007 5321
rect 25590 5312 25596 5364
rect 25648 5352 25654 5364
rect 27246 5352 27252 5364
rect 25648 5324 27252 5352
rect 25648 5312 25654 5324
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 27982 5312 27988 5364
rect 28040 5352 28046 5364
rect 29641 5355 29699 5361
rect 29641 5352 29653 5355
rect 28040 5324 29653 5352
rect 28040 5312 28046 5324
rect 29641 5321 29653 5324
rect 29687 5352 29699 5355
rect 34790 5352 34796 5364
rect 29687 5324 34796 5352
rect 29687 5321 29699 5324
rect 29641 5315 29699 5321
rect 34790 5312 34796 5324
rect 34848 5352 34854 5364
rect 35066 5352 35072 5364
rect 34848 5324 35072 5352
rect 34848 5312 34854 5324
rect 35066 5312 35072 5324
rect 35124 5312 35130 5364
rect 37182 5312 37188 5364
rect 37240 5352 37246 5364
rect 37277 5355 37335 5361
rect 37277 5352 37289 5355
rect 37240 5324 37289 5352
rect 37240 5312 37246 5324
rect 37277 5321 37289 5324
rect 37323 5321 37335 5355
rect 37277 5315 37335 5321
rect 25866 5284 25872 5296
rect 20640 5256 23888 5284
rect 24688 5256 25872 5284
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 13372 5188 13921 5216
rect 10100 5120 10824 5148
rect 11885 5151 11943 5157
rect 10100 5108 10106 5120
rect 11885 5117 11897 5151
rect 11931 5148 11943 5151
rect 12802 5148 12808 5160
rect 11931 5120 12808 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 13170 5108 13176 5160
rect 13228 5148 13234 5160
rect 13372 5148 13400 5188
rect 13909 5185 13921 5188
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 13228 5120 13400 5148
rect 13449 5151 13507 5157
rect 13228 5108 13234 5120
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 13538 5148 13544 5160
rect 13495 5120 13544 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 14936 5148 14964 5179
rect 15010 5176 15016 5228
rect 15068 5216 15074 5228
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 15068 5188 15301 5216
rect 15068 5176 15074 5188
rect 15289 5185 15301 5188
rect 15335 5216 15347 5219
rect 15335 5188 15424 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15396 5148 15424 5188
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16632 5188 17049 5216
rect 16632 5176 16638 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5216 19027 5219
rect 19242 5216 19248 5228
rect 19015 5188 19248 5216
rect 19015 5185 19027 5188
rect 18969 5179 19027 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 19610 5216 19616 5228
rect 19571 5188 19616 5216
rect 19610 5176 19616 5188
rect 19668 5176 19674 5228
rect 20070 5176 20076 5228
rect 20128 5216 20134 5228
rect 20640 5225 20668 5256
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 20128 5188 20637 5216
rect 20128 5176 20134 5188
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 21174 5176 21180 5228
rect 21232 5216 21238 5228
rect 22934 5219 22992 5225
rect 22934 5216 22946 5219
rect 21232 5188 22946 5216
rect 21232 5176 21238 5188
rect 22934 5185 22946 5188
rect 22980 5185 22992 5219
rect 22934 5179 22992 5185
rect 23201 5219 23259 5225
rect 23201 5185 23213 5219
rect 23247 5216 23259 5219
rect 23474 5216 23480 5228
rect 23247 5188 23480 5216
rect 23247 5185 23259 5188
rect 23201 5179 23259 5185
rect 23474 5176 23480 5188
rect 23532 5176 23538 5228
rect 23658 5216 23664 5228
rect 23619 5188 23664 5216
rect 23658 5176 23664 5188
rect 23716 5176 23722 5228
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 14016 5120 15332 5148
rect 15396 5120 16681 5148
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5080 10379 5083
rect 10367 5052 12296 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 10226 5012 10232 5024
rect 9140 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 11606 5012 11612 5024
rect 11567 4984 11612 5012
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 12032 4984 12173 5012
rect 12032 4972 12038 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12268 5012 12296 5052
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 13081 5083 13139 5089
rect 13081 5080 13093 5083
rect 12400 5052 13093 5080
rect 12400 5040 12406 5052
rect 13081 5049 13093 5052
rect 13127 5049 13139 5083
rect 13081 5043 13139 5049
rect 14016 5012 14044 5120
rect 15304 5092 15332 5120
rect 16669 5117 16681 5120
rect 16715 5148 16727 5151
rect 16850 5148 16856 5160
rect 16715 5120 16856 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5148 18567 5151
rect 19150 5148 19156 5160
rect 18555 5120 19156 5148
rect 18555 5117 18567 5120
rect 18509 5111 18567 5117
rect 19150 5108 19156 5120
rect 19208 5108 19214 5160
rect 20530 5148 20536 5160
rect 19260 5120 20536 5148
rect 14642 5040 14648 5092
rect 14700 5080 14706 5092
rect 15194 5080 15200 5092
rect 14700 5052 15200 5080
rect 14700 5040 14706 5052
rect 12268 4984 14044 5012
rect 14093 5015 14151 5021
rect 12161 4975 12219 4981
rect 14093 4981 14105 5015
rect 14139 5012 14151 5015
rect 14734 5012 14740 5024
rect 14139 4984 14740 5012
rect 14139 4981 14151 4984
rect 14093 4975 14151 4981
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 14844 5021 14872 5052
rect 15194 5040 15200 5052
rect 15252 5040 15258 5092
rect 15286 5040 15292 5092
rect 15344 5040 15350 5092
rect 16117 5083 16175 5089
rect 16117 5049 16129 5083
rect 16163 5080 16175 5083
rect 17770 5080 17776 5092
rect 16163 5052 17776 5080
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 17770 5040 17776 5052
rect 17828 5040 17834 5092
rect 19260 5080 19288 5120
rect 20530 5108 20536 5120
rect 20588 5148 20594 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20588 5120 20821 5148
rect 20588 5108 20594 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20809 5111 20867 5117
rect 19076 5052 19288 5080
rect 23860 5080 23888 5256
rect 25866 5244 25872 5256
rect 25924 5284 25930 5296
rect 26053 5287 26111 5293
rect 26053 5284 26065 5287
rect 25924 5256 26065 5284
rect 25924 5244 25930 5256
rect 26053 5253 26065 5256
rect 26099 5253 26111 5287
rect 26053 5247 26111 5253
rect 26237 5287 26295 5293
rect 26237 5253 26249 5287
rect 26283 5284 26295 5287
rect 26602 5284 26608 5296
rect 26283 5256 26608 5284
rect 26283 5253 26295 5256
rect 26237 5247 26295 5253
rect 26602 5244 26608 5256
rect 26660 5244 26666 5296
rect 23937 5219 23995 5225
rect 23937 5185 23949 5219
rect 23983 5216 23995 5219
rect 25130 5216 25136 5228
rect 23983 5188 25136 5216
rect 23983 5185 23995 5188
rect 23937 5179 23995 5185
rect 25130 5176 25136 5188
rect 25188 5216 25194 5228
rect 26970 5216 26976 5228
rect 25188 5188 26976 5216
rect 25188 5176 25194 5188
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 27264 5225 27292 5312
rect 28261 5287 28319 5293
rect 28261 5253 28273 5287
rect 28307 5284 28319 5287
rect 29454 5284 29460 5296
rect 28307 5256 29460 5284
rect 28307 5253 28319 5256
rect 28261 5247 28319 5253
rect 29454 5244 29460 5256
rect 29512 5244 29518 5296
rect 30926 5244 30932 5296
rect 30984 5284 30990 5296
rect 32217 5287 32275 5293
rect 30984 5256 31616 5284
rect 30984 5244 30990 5256
rect 31588 5228 31616 5256
rect 32217 5253 32229 5287
rect 32263 5284 32275 5287
rect 32674 5284 32680 5296
rect 32263 5256 32680 5284
rect 32263 5253 32275 5256
rect 32217 5247 32275 5253
rect 32674 5244 32680 5256
rect 32732 5244 32738 5296
rect 33502 5244 33508 5296
rect 33560 5284 33566 5296
rect 33781 5287 33839 5293
rect 33781 5284 33793 5287
rect 33560 5256 33793 5284
rect 33560 5244 33566 5256
rect 33781 5253 33793 5256
rect 33827 5253 33839 5287
rect 33962 5284 33968 5296
rect 33923 5256 33968 5284
rect 33781 5247 33839 5253
rect 27136 5219 27194 5225
rect 27136 5216 27148 5219
rect 27080 5188 27148 5216
rect 26421 5151 26479 5157
rect 26421 5117 26433 5151
rect 26467 5148 26479 5151
rect 27080 5148 27108 5188
rect 27136 5185 27148 5188
rect 27182 5185 27194 5219
rect 27136 5179 27194 5185
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 27338 5176 27344 5228
rect 27396 5216 27402 5228
rect 28074 5216 28080 5228
rect 27396 5188 27441 5216
rect 28035 5188 28080 5216
rect 27396 5176 27402 5188
rect 28074 5176 28080 5188
rect 28132 5176 28138 5228
rect 28166 5176 28172 5228
rect 28224 5216 28230 5228
rect 28445 5219 28503 5225
rect 28445 5216 28457 5219
rect 28224 5188 28457 5216
rect 28224 5176 28230 5188
rect 28445 5185 28457 5188
rect 28491 5185 28503 5219
rect 28445 5179 28503 5185
rect 31294 5176 31300 5228
rect 31352 5225 31358 5228
rect 31352 5216 31364 5225
rect 31570 5216 31576 5228
rect 31352 5188 31397 5216
rect 31483 5188 31576 5216
rect 31352 5179 31364 5188
rect 31352 5176 31358 5179
rect 31570 5176 31576 5188
rect 31628 5176 31634 5228
rect 26467 5120 27108 5148
rect 26467 5117 26479 5120
rect 26421 5111 26479 5117
rect 28718 5080 28724 5092
rect 23860 5052 28724 5080
rect 14829 5015 14887 5021
rect 14829 4981 14841 5015
rect 14875 4981 14887 5015
rect 14829 4975 14887 4981
rect 17678 4972 17684 5024
rect 17736 5012 17742 5024
rect 19076 5012 19104 5052
rect 28718 5040 28724 5052
rect 28776 5040 28782 5092
rect 30193 5083 30251 5089
rect 30193 5049 30205 5083
rect 30239 5080 30251 5083
rect 30466 5080 30472 5092
rect 30239 5052 30472 5080
rect 30239 5049 30251 5052
rect 30193 5043 30251 5049
rect 30466 5040 30472 5052
rect 30524 5040 30530 5092
rect 33796 5080 33824 5247
rect 33962 5244 33968 5256
rect 34020 5244 34026 5296
rect 34054 5244 34060 5296
rect 34112 5284 34118 5296
rect 34149 5287 34207 5293
rect 34149 5284 34161 5287
rect 34112 5256 34161 5284
rect 34112 5244 34118 5256
rect 34149 5253 34161 5256
rect 34195 5253 34207 5287
rect 34149 5247 34207 5253
rect 34606 5244 34612 5296
rect 34664 5284 34670 5296
rect 35618 5284 35624 5296
rect 34664 5256 34928 5284
rect 34664 5244 34670 5256
rect 34238 5176 34244 5228
rect 34296 5216 34302 5228
rect 34900 5225 34928 5256
rect 34992 5256 35624 5284
rect 34992 5225 35020 5256
rect 35618 5244 35624 5256
rect 35676 5244 35682 5296
rect 38105 5287 38163 5293
rect 38105 5284 38117 5287
rect 36188 5256 38117 5284
rect 34701 5219 34759 5225
rect 34701 5216 34713 5219
rect 34296 5188 34713 5216
rect 34296 5176 34302 5188
rect 34701 5185 34713 5188
rect 34747 5185 34759 5219
rect 34701 5179 34759 5185
rect 34885 5219 34943 5225
rect 34885 5185 34897 5219
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 34977 5219 35035 5225
rect 34977 5185 34989 5219
rect 35023 5185 35035 5219
rect 34977 5179 35035 5185
rect 35069 5219 35127 5225
rect 35069 5185 35081 5219
rect 35115 5185 35127 5219
rect 35986 5216 35992 5228
rect 35947 5188 35992 5216
rect 35069 5179 35127 5185
rect 34054 5108 34060 5160
rect 34112 5148 34118 5160
rect 35084 5148 35112 5179
rect 35986 5176 35992 5188
rect 36044 5176 36050 5228
rect 36188 5225 36216 5256
rect 38105 5253 38117 5256
rect 38151 5253 38163 5287
rect 38286 5284 38292 5296
rect 38247 5256 38292 5284
rect 38105 5247 38163 5253
rect 38286 5244 38292 5256
rect 38344 5244 38350 5296
rect 36173 5219 36231 5225
rect 36173 5185 36185 5219
rect 36219 5185 36231 5219
rect 36173 5179 36231 5185
rect 36265 5219 36323 5225
rect 36265 5185 36277 5219
rect 36311 5185 36323 5219
rect 36265 5179 36323 5185
rect 34112 5120 35112 5148
rect 34112 5108 34118 5120
rect 35618 5108 35624 5160
rect 35676 5148 35682 5160
rect 36280 5148 36308 5179
rect 36354 5176 36360 5228
rect 36412 5216 36418 5228
rect 36412 5188 36457 5216
rect 36412 5176 36418 5188
rect 36814 5176 36820 5228
rect 36872 5216 36878 5228
rect 37461 5219 37519 5225
rect 37461 5216 37473 5219
rect 36872 5188 37473 5216
rect 36872 5176 36878 5188
rect 37461 5185 37473 5188
rect 37507 5185 37519 5219
rect 37461 5179 37519 5185
rect 37645 5219 37703 5225
rect 37645 5185 37657 5219
rect 37691 5185 37703 5219
rect 37645 5179 37703 5185
rect 38473 5219 38531 5225
rect 38473 5185 38485 5219
rect 38519 5216 38531 5219
rect 38746 5216 38752 5228
rect 38519 5188 38752 5216
rect 38519 5185 38531 5188
rect 38473 5179 38531 5185
rect 35676 5120 36308 5148
rect 37660 5148 37688 5179
rect 38488 5148 38516 5179
rect 38746 5176 38752 5188
rect 38804 5176 38810 5228
rect 37660 5120 38516 5148
rect 35676 5108 35682 5120
rect 37660 5080 37688 5120
rect 58802 5108 58808 5160
rect 58860 5148 58866 5160
rect 59449 5151 59507 5157
rect 59449 5148 59461 5151
rect 58860 5120 59461 5148
rect 58860 5108 58866 5120
rect 59449 5117 59461 5120
rect 59495 5117 59507 5151
rect 59449 5111 59507 5117
rect 33796 5052 37688 5080
rect 59262 5040 59268 5092
rect 59320 5080 59326 5092
rect 60093 5083 60151 5089
rect 60093 5080 60105 5083
rect 59320 5052 60105 5080
rect 59320 5040 59326 5052
rect 60093 5049 60105 5052
rect 60139 5049 60151 5083
rect 60093 5043 60151 5049
rect 17736 4984 19104 5012
rect 19153 5015 19211 5021
rect 17736 4972 17742 4984
rect 19153 4981 19165 5015
rect 19199 5012 19211 5015
rect 19426 5012 19432 5024
rect 19199 4984 19432 5012
rect 19199 4981 19211 4984
rect 19153 4975 19211 4981
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 19797 5015 19855 5021
rect 19797 4981 19809 5015
rect 19843 5012 19855 5015
rect 19978 5012 19984 5024
rect 19843 4984 19984 5012
rect 19843 4981 19855 4984
rect 19797 4975 19855 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20257 5015 20315 5021
rect 20257 4981 20269 5015
rect 20303 5012 20315 5015
rect 20346 5012 20352 5024
rect 20303 4984 20352 5012
rect 20303 4981 20315 4984
rect 20257 4975 20315 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 27338 5012 27344 5024
rect 20956 4984 27344 5012
rect 20956 4972 20962 4984
rect 27338 4972 27344 4984
rect 27396 4972 27402 5024
rect 27614 5012 27620 5024
rect 27575 4984 27620 5012
rect 27614 4972 27620 4984
rect 27672 4972 27678 5024
rect 35342 5012 35348 5024
rect 35303 4984 35348 5012
rect 35342 4972 35348 4984
rect 35400 4972 35406 5024
rect 36630 5012 36636 5024
rect 36591 4984 36636 5012
rect 36630 4972 36636 4984
rect 36688 4972 36694 5024
rect 58710 4972 58716 5024
rect 58768 5012 58774 5024
rect 58805 5015 58863 5021
rect 58805 5012 58817 5015
rect 58768 4984 58817 5012
rect 58768 4972 58774 4984
rect 58805 4981 58817 4984
rect 58851 4981 58863 5015
rect 67634 5012 67640 5024
rect 67595 4984 67640 5012
rect 58805 4975 58863 4981
rect 67634 4972 67640 4984
rect 67692 4972 67698 5024
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 5626 4808 5632 4820
rect 5587 4780 5632 4808
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10410 4808 10416 4820
rect 10008 4780 10416 4808
rect 10008 4768 10014 4780
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 14642 4808 14648 4820
rect 12952 4780 14648 4808
rect 12952 4768 12958 4780
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 21174 4808 21180 4820
rect 21135 4780 21180 4808
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 23569 4811 23627 4817
rect 23569 4777 23581 4811
rect 23615 4808 23627 4811
rect 23658 4808 23664 4820
rect 23615 4780 23664 4808
rect 23615 4777 23627 4780
rect 23569 4771 23627 4777
rect 23658 4768 23664 4780
rect 23716 4768 23722 4820
rect 30742 4768 30748 4820
rect 30800 4808 30806 4820
rect 31205 4811 31263 4817
rect 31205 4808 31217 4811
rect 30800 4780 31217 4808
rect 30800 4768 30806 4780
rect 31205 4777 31217 4780
rect 31251 4777 31263 4811
rect 31205 4771 31263 4777
rect 32125 4811 32183 4817
rect 32125 4777 32137 4811
rect 32171 4808 32183 4811
rect 33226 4808 33232 4820
rect 32171 4780 33232 4808
rect 32171 4777 32183 4780
rect 32125 4771 32183 4777
rect 33226 4768 33232 4780
rect 33284 4768 33290 4820
rect 34790 4768 34796 4820
rect 34848 4808 34854 4820
rect 34885 4811 34943 4817
rect 34885 4808 34897 4811
rect 34848 4780 34897 4808
rect 34848 4768 34854 4780
rect 34885 4777 34897 4780
rect 34931 4777 34943 4811
rect 34885 4771 34943 4777
rect 38286 4768 38292 4820
rect 38344 4808 38350 4820
rect 38657 4811 38715 4817
rect 38657 4808 38669 4811
rect 38344 4780 38669 4808
rect 38344 4768 38350 4780
rect 38657 4777 38669 4780
rect 38703 4777 38715 4811
rect 38657 4771 38715 4777
rect 4249 4743 4307 4749
rect 4249 4709 4261 4743
rect 4295 4740 4307 4743
rect 6454 4740 6460 4752
rect 4295 4712 6460 4740
rect 4295 4709 4307 4712
rect 4249 4703 4307 4709
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 9033 4743 9091 4749
rect 9033 4709 9045 4743
rect 9079 4740 9091 4743
rect 11974 4740 11980 4752
rect 9079 4712 11980 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 12161 4743 12219 4749
rect 12161 4709 12173 4743
rect 12207 4709 12219 4743
rect 12161 4703 12219 4709
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4672 1639 4675
rect 6914 4672 6920 4684
rect 1627 4644 6920 4672
rect 1627 4641 1639 4644
rect 1581 4635 1639 4641
rect 6914 4632 6920 4644
rect 6972 4672 6978 4684
rect 6972 4644 7144 4672
rect 6972 4632 6978 4644
rect 2590 4604 2596 4616
rect 2551 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4604 4123 4607
rect 4614 4604 4620 4616
rect 4111 4576 4620 4604
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 7116 4613 7144 4644
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9582 4672 9588 4684
rect 8904 4644 9588 4672
rect 8904 4632 8910 4644
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4672 10471 4675
rect 10502 4672 10508 4684
rect 10459 4644 10508 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 10870 4672 10876 4684
rect 10704 4644 10876 4672
rect 7101 4607 7159 4613
rect 4764 4576 4809 4604
rect 4764 4564 4770 4576
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 8110 4604 8116 4616
rect 8071 4576 8116 4604
rect 7101 4567 7159 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 9674 4604 9680 4616
rect 9635 4576 9680 4604
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 10704 4613 10732 4644
rect 10870 4632 10876 4644
rect 10928 4672 10934 4684
rect 11330 4672 11336 4684
rect 10928 4644 11336 4672
rect 10928 4632 10934 4644
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11422 4632 11428 4684
rect 11480 4632 11486 4684
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 12176 4672 12204 4703
rect 13538 4700 13544 4752
rect 13596 4700 13602 4752
rect 14918 4700 14924 4752
rect 14976 4740 14982 4752
rect 18601 4743 18659 4749
rect 18601 4740 18613 4743
rect 14976 4712 18613 4740
rect 14976 4700 14982 4712
rect 18601 4709 18613 4712
rect 18647 4740 18659 4743
rect 20070 4740 20076 4752
rect 18647 4712 20076 4740
rect 18647 4709 18659 4712
rect 18601 4703 18659 4709
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 25777 4743 25835 4749
rect 25777 4709 25789 4743
rect 25823 4740 25835 4743
rect 25823 4712 26464 4740
rect 25823 4709 25835 4712
rect 25777 4703 25835 4709
rect 11940 4644 12204 4672
rect 11940 4632 11946 4644
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 13556 4672 13584 4700
rect 12308 4644 12353 4672
rect 13556 4644 14504 4672
rect 12308 4632 12314 4644
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4573 10747 4607
rect 11146 4604 11152 4616
rect 11107 4576 11152 4604
rect 10689 4567 10747 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11440 4604 11468 4632
rect 11974 4604 11980 4616
rect 11440 4576 11980 4604
rect 11974 4564 11980 4576
rect 12032 4613 12038 4616
rect 12032 4607 12090 4613
rect 12032 4573 12044 4607
rect 12078 4573 12090 4607
rect 12032 4567 12090 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13630 4604 13636 4616
rect 13587 4576 13636 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 12032 4564 12038 4567
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 14476 4613 14504 4644
rect 17678 4632 17684 4684
rect 17736 4672 17742 4684
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17736 4644 17969 4672
rect 17736 4632 17742 4644
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 20254 4672 20260 4684
rect 17957 4635 18015 4641
rect 20180 4644 20260 4672
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 15010 4604 15016 4616
rect 14783 4576 15016 4604
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 15010 4564 15016 4576
rect 15068 4564 15074 4616
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4604 15163 4607
rect 15286 4604 15292 4616
rect 15151 4576 15292 4604
rect 15151 4573 15163 4576
rect 15105 4567 15163 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 15562 4604 15568 4616
rect 15523 4576 15568 4604
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 16850 4604 16856 4616
rect 16811 4576 16856 4604
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 17494 4604 17500 4616
rect 17184 4576 17500 4604
rect 17184 4564 17190 4576
rect 17494 4564 17500 4576
rect 17552 4604 17558 4616
rect 17773 4607 17831 4613
rect 17773 4604 17785 4607
rect 17552 4576 17785 4604
rect 17552 4564 17558 4576
rect 17773 4573 17785 4576
rect 17819 4573 17831 4607
rect 17773 4567 17831 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 20070 4604 20076 4616
rect 19751 4576 20076 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20180 4613 20208 4644
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 21634 4672 21640 4684
rect 21595 4644 21640 4672
rect 21634 4632 21640 4644
rect 21692 4632 21698 4684
rect 24210 4632 24216 4684
rect 24268 4672 24274 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 24268 4644 24409 4672
rect 24268 4632 24274 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4573 20223 4607
rect 20346 4604 20352 4616
rect 20307 4576 20352 4604
rect 20165 4567 20223 4573
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 26436 4613 26464 4712
rect 57238 4700 57244 4752
rect 57296 4740 57302 4752
rect 57885 4743 57943 4749
rect 57885 4740 57897 4743
rect 57296 4712 57897 4740
rect 57296 4700 57302 4712
rect 57885 4709 57897 4712
rect 57931 4709 57943 4743
rect 57885 4703 57943 4709
rect 58250 4700 58256 4752
rect 58308 4740 58314 4752
rect 59173 4743 59231 4749
rect 59173 4740 59185 4743
rect 58308 4712 59185 4740
rect 58308 4700 58314 4712
rect 59173 4709 59185 4712
rect 59219 4709 59231 4743
rect 59173 4703 59231 4709
rect 36630 4632 36636 4684
rect 36688 4672 36694 4684
rect 36688 4644 37412 4672
rect 36688 4632 36694 4644
rect 20533 4607 20591 4613
rect 20533 4573 20545 4607
rect 20579 4604 20591 4607
rect 20993 4607 21051 4613
rect 20993 4604 21005 4607
rect 20579 4576 21005 4604
rect 20579 4573 20591 4576
rect 20533 4567 20591 4573
rect 20993 4573 21005 4576
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 26421 4607 26479 4613
rect 26421 4573 26433 4607
rect 26467 4604 26479 4607
rect 26510 4604 26516 4616
rect 26467 4576 26516 4604
rect 26467 4573 26479 4576
rect 26421 4567 26479 4573
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 28445 4607 28503 4613
rect 28445 4573 28457 4607
rect 28491 4604 28503 4607
rect 28994 4604 29000 4616
rect 28491 4576 29000 4604
rect 28491 4573 28503 4576
rect 28445 4567 28503 4573
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 31570 4564 31576 4616
rect 31628 4604 31634 4616
rect 33505 4607 33563 4613
rect 33505 4604 33517 4607
rect 31628 4576 33517 4604
rect 31628 4564 31634 4576
rect 33505 4573 33517 4576
rect 33551 4604 33563 4607
rect 35158 4604 35164 4616
rect 33551 4576 35164 4604
rect 33551 4573 33563 4576
rect 33505 4567 33563 4573
rect 35158 4564 35164 4576
rect 35216 4604 35222 4616
rect 35437 4607 35495 4613
rect 35437 4604 35449 4607
rect 35216 4576 35449 4604
rect 35216 4564 35222 4576
rect 35437 4573 35449 4576
rect 35483 4573 35495 4607
rect 35437 4567 35495 4573
rect 11422 4536 11428 4548
rect 4908 4508 11428 4536
rect 2133 4471 2191 4477
rect 2133 4437 2145 4471
rect 2179 4468 2191 4471
rect 2498 4468 2504 4480
rect 2179 4440 2504 4468
rect 2179 4437 2191 4440
rect 2133 4431 2191 4437
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 4908 4477 4936 4508
rect 11422 4496 11428 4508
rect 11480 4536 11486 4548
rect 11885 4539 11943 4545
rect 11885 4536 11897 4539
rect 11480 4508 11897 4536
rect 11480 4496 11486 4508
rect 11885 4505 11897 4508
rect 11931 4505 11943 4539
rect 11885 4499 11943 4505
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 12621 4539 12679 4545
rect 12621 4536 12633 4539
rect 12400 4508 12633 4536
rect 12400 4496 12406 4508
rect 12621 4505 12633 4508
rect 12667 4536 12679 4539
rect 13998 4536 14004 4548
rect 12667 4508 14004 4536
rect 12667 4505 12679 4508
rect 12621 4499 12679 4505
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 18966 4536 18972 4548
rect 14936 4508 18972 4536
rect 4893 4471 4951 4477
rect 2832 4440 2877 4468
rect 2832 4428 2838 4440
rect 4893 4437 4905 4471
rect 4939 4437 4951 4471
rect 4893 4431 4951 4437
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7064 4440 8033 4468
rect 7064 4428 7070 4440
rect 8021 4437 8033 4440
rect 8067 4468 8079 4471
rect 8110 4468 8116 4480
rect 8067 4440 8116 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 8754 4428 8760 4480
rect 8812 4468 8818 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 8812 4440 10149 4468
rect 8812 4428 8818 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 11333 4471 11391 4477
rect 11333 4437 11345 4471
rect 11379 4468 11391 4471
rect 11698 4468 11704 4480
rect 11379 4440 11704 4468
rect 11379 4437 11391 4440
rect 11333 4431 11391 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 13354 4468 13360 4480
rect 13315 4440 13360 4468
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 14936 4477 14964 4508
rect 18966 4496 18972 4508
rect 19024 4496 19030 4548
rect 19242 4496 19248 4548
rect 19300 4536 19306 4548
rect 22833 4539 22891 4545
rect 22833 4536 22845 4539
rect 19300 4508 22845 4536
rect 19300 4496 19306 4508
rect 22833 4505 22845 4508
rect 22879 4505 22891 4539
rect 22833 4499 22891 4505
rect 24664 4539 24722 4545
rect 24664 4505 24676 4539
rect 24710 4536 24722 4539
rect 25222 4536 25228 4548
rect 24710 4508 25228 4536
rect 24710 4505 24722 4508
rect 24664 4499 24722 4505
rect 25222 4496 25228 4508
rect 25280 4496 25286 4548
rect 25866 4496 25872 4548
rect 25924 4536 25930 4548
rect 26605 4539 26663 4545
rect 26605 4536 26617 4539
rect 25924 4508 26617 4536
rect 25924 4496 25930 4508
rect 26605 4505 26617 4508
rect 26651 4536 26663 4539
rect 28166 4536 28172 4548
rect 26651 4508 28172 4536
rect 26651 4505 26663 4508
rect 26605 4499 26663 4505
rect 28166 4496 28172 4508
rect 28224 4536 28230 4548
rect 28261 4539 28319 4545
rect 28261 4536 28273 4539
rect 28224 4508 28273 4536
rect 28224 4496 28230 4508
rect 28261 4505 28273 4508
rect 28307 4505 28319 4539
rect 28261 4499 28319 4505
rect 30834 4496 30840 4548
rect 30892 4536 30898 4548
rect 33260 4539 33318 4545
rect 30892 4508 33180 4536
rect 30892 4496 30898 4508
rect 14921 4471 14979 4477
rect 14921 4437 14933 4471
rect 14967 4437 14979 4471
rect 15746 4468 15752 4480
rect 15707 4440 15752 4468
rect 14921 4431 14979 4437
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 16666 4468 16672 4480
rect 16627 4440 16672 4468
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17405 4471 17463 4477
rect 17405 4437 17417 4471
rect 17451 4468 17463 4471
rect 17494 4468 17500 4480
rect 17451 4440 17500 4468
rect 17451 4437 17463 4440
rect 17405 4431 17463 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 17920 4440 17965 4468
rect 17920 4428 17926 4440
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 20346 4468 20352 4480
rect 19668 4440 20352 4468
rect 19668 4428 19674 4440
rect 20346 4428 20352 4440
rect 20404 4468 20410 4480
rect 22281 4471 22339 4477
rect 22281 4468 22293 4471
rect 20404 4440 22293 4468
rect 20404 4428 20410 4440
rect 22281 4437 22293 4440
rect 22327 4437 22339 4471
rect 22281 4431 22339 4437
rect 25682 4428 25688 4480
rect 25740 4468 25746 4480
rect 26237 4471 26295 4477
rect 26237 4468 26249 4471
rect 25740 4440 26249 4468
rect 25740 4428 25746 4440
rect 26237 4437 26249 4440
rect 26283 4437 26295 4471
rect 26237 4431 26295 4437
rect 28534 4428 28540 4480
rect 28592 4468 28598 4480
rect 28629 4471 28687 4477
rect 28629 4468 28641 4471
rect 28592 4440 28641 4468
rect 28592 4428 28598 4440
rect 28629 4437 28641 4440
rect 28675 4437 28687 4471
rect 33152 4468 33180 4508
rect 33260 4505 33272 4539
rect 33306 4536 33318 4539
rect 35342 4536 35348 4548
rect 33306 4508 35348 4536
rect 33306 4505 33318 4508
rect 33260 4499 33318 4505
rect 35342 4496 35348 4508
rect 35400 4496 35406 4548
rect 34054 4468 34060 4480
rect 33152 4440 34060 4468
rect 28629 4431 28687 4437
rect 34054 4428 34060 4440
rect 34112 4428 34118 4480
rect 35452 4468 35480 4567
rect 35526 4564 35532 4616
rect 35584 4604 35590 4616
rect 35704 4607 35762 4613
rect 35704 4604 35716 4607
rect 35584 4576 35716 4604
rect 35584 4564 35590 4576
rect 35704 4573 35716 4576
rect 35750 4573 35762 4607
rect 37274 4604 37280 4616
rect 35704 4567 35762 4573
rect 35820 4576 37280 4604
rect 35820 4468 35848 4576
rect 37274 4564 37280 4576
rect 37332 4564 37338 4616
rect 37384 4604 37412 4644
rect 58894 4632 58900 4684
rect 58952 4672 58958 4684
rect 60461 4675 60519 4681
rect 60461 4672 60473 4675
rect 58952 4644 60473 4672
rect 58952 4632 58958 4644
rect 60461 4641 60473 4644
rect 60507 4641 60519 4675
rect 60461 4635 60519 4641
rect 37533 4607 37591 4613
rect 37533 4604 37545 4607
rect 37384 4576 37545 4604
rect 37533 4573 37545 4576
rect 37579 4573 37591 4607
rect 37533 4567 37591 4573
rect 57146 4564 57152 4616
rect 57204 4604 57210 4616
rect 57241 4607 57299 4613
rect 57241 4604 57253 4607
rect 57204 4576 57253 4604
rect 57204 4564 57210 4576
rect 57241 4573 57253 4576
rect 57287 4573 57299 4607
rect 57241 4567 57299 4573
rect 57606 4564 57612 4616
rect 57664 4604 57670 4616
rect 58529 4607 58587 4613
rect 58529 4604 58541 4607
rect 57664 4576 58541 4604
rect 57664 4564 57670 4576
rect 58529 4573 58541 4576
rect 58575 4573 58587 4607
rect 58529 4567 58587 4573
rect 36814 4468 36820 4480
rect 35452 4440 35848 4468
rect 36775 4440 36820 4468
rect 36814 4428 36820 4440
rect 36872 4428 36878 4480
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 2041 4267 2099 4273
rect 2041 4233 2053 4267
rect 2087 4264 2099 4267
rect 2130 4264 2136 4276
rect 2087 4236 2136 4264
rect 2087 4233 2099 4236
rect 2041 4227 2099 4233
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 7800 4236 8493 4264
rect 7800 4224 7806 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8846 4264 8852 4276
rect 8807 4236 8852 4264
rect 8481 4227 8539 4233
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 8996 4236 9041 4264
rect 8996 4224 9002 4236
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 10410 4264 10416 4276
rect 9916 4236 10416 4264
rect 9916 4224 9922 4236
rect 10410 4224 10416 4236
rect 10468 4264 10474 4276
rect 10686 4264 10692 4276
rect 10744 4273 10750 4276
rect 10744 4267 10763 4273
rect 10468 4236 10692 4264
rect 10468 4224 10474 4236
rect 10686 4224 10692 4236
rect 10751 4233 10763 4267
rect 10870 4264 10876 4276
rect 10831 4236 10876 4264
rect 10744 4227 10763 4233
rect 10744 4224 10750 4227
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 12066 4264 12072 4276
rect 11480 4236 12072 4264
rect 11480 4224 11486 4236
rect 12066 4224 12072 4236
rect 12124 4264 12130 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 12124 4236 12173 4264
rect 12124 4224 12130 4236
rect 12161 4233 12173 4236
rect 12207 4264 12219 4267
rect 12342 4264 12348 4276
rect 12207 4236 12348 4264
rect 12207 4233 12219 4236
rect 12161 4227 12219 4233
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 14461 4267 14519 4273
rect 14461 4264 14473 4267
rect 13320 4236 14473 4264
rect 13320 4224 13326 4236
rect 14461 4233 14473 4236
rect 14507 4233 14519 4267
rect 14461 4227 14519 4233
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 17313 4267 17371 4273
rect 17313 4264 17325 4267
rect 16908 4236 17325 4264
rect 16908 4224 16914 4236
rect 17313 4233 17325 4236
rect 17359 4233 17371 4267
rect 17313 4227 17371 4233
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 21634 4264 21640 4276
rect 18012 4236 21640 4264
rect 18012 4224 18018 4236
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 26602 4224 26608 4276
rect 26660 4264 26666 4276
rect 26973 4267 27031 4273
rect 26973 4264 26985 4267
rect 26660 4236 26985 4264
rect 26660 4224 26666 4236
rect 26973 4233 26985 4236
rect 27019 4233 27031 4267
rect 26973 4227 27031 4233
rect 28994 4224 29000 4276
rect 29052 4264 29058 4276
rect 29457 4267 29515 4273
rect 29457 4264 29469 4267
rect 29052 4236 29469 4264
rect 29052 4224 29058 4236
rect 29457 4233 29469 4236
rect 29503 4233 29515 4267
rect 29457 4227 29515 4233
rect 33781 4267 33839 4273
rect 33781 4233 33793 4267
rect 33827 4264 33839 4267
rect 33962 4264 33968 4276
rect 33827 4236 33968 4264
rect 33827 4233 33839 4236
rect 33781 4227 33839 4233
rect 33962 4224 33968 4236
rect 34020 4224 34026 4276
rect 35897 4267 35955 4273
rect 35897 4233 35909 4267
rect 35943 4264 35955 4267
rect 36262 4264 36268 4276
rect 35943 4236 36268 4264
rect 35943 4233 35955 4236
rect 35897 4227 35955 4233
rect 36262 4224 36268 4236
rect 36320 4224 36326 4276
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 3574 4199 3632 4205
rect 3574 4196 3586 4199
rect 2832 4168 3586 4196
rect 2832 4156 2838 4168
rect 3574 4165 3586 4168
rect 3620 4165 3632 4199
rect 3574 4159 3632 4165
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 7009 4199 7067 4205
rect 7009 4196 7021 4199
rect 5675 4168 7021 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 7009 4165 7021 4168
rect 7055 4196 7067 4199
rect 8754 4196 8760 4208
rect 7055 4168 8760 4196
rect 7055 4165 7067 4168
rect 7009 4159 7067 4165
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 10502 4196 10508 4208
rect 9646 4168 10180 4196
rect 10463 4168 10508 4196
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3200 4100 3341 4128
rect 3200 4088 3206 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 7190 4128 7196 4140
rect 4764 4100 7196 4128
rect 4764 4088 4770 4100
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7616 4100 7665 4128
rect 7616 4088 7622 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7800 4100 7849 4128
rect 7800 4088 7806 4100
rect 7837 4097 7849 4100
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 7984 4100 8029 4128
rect 7984 4088 7990 4100
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 9646 4128 9674 4168
rect 8168 4100 9674 4128
rect 8168 4088 8174 4100
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 9916 4100 9961 4128
rect 9916 4088 9922 4100
rect 1854 4060 1860 4072
rect 1815 4032 1860 4060
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4060 2007 4063
rect 1995 4032 2774 4060
rect 1995 4029 2007 4032
rect 1949 4023 2007 4029
rect 2130 3884 2136 3936
rect 2188 3924 2194 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2188 3896 2421 3924
rect 2188 3884 2194 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2746 3924 2774 4032
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 9033 4063 9091 4069
rect 9033 4060 9045 4063
rect 8812 4032 9045 4060
rect 8812 4020 8818 4032
rect 9033 4029 9045 4032
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 9674 4060 9680 4072
rect 9180 4032 9680 4060
rect 9180 4020 9186 4032
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4060 10103 4063
rect 10152 4060 10180 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 11609 4199 11667 4205
rect 11609 4165 11621 4199
rect 11655 4196 11667 4199
rect 11882 4196 11888 4208
rect 11655 4168 11888 4196
rect 11655 4165 11667 4168
rect 11609 4159 11667 4165
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 20806 4196 20812 4208
rect 18288 4168 19472 4196
rect 20767 4168 20812 4196
rect 18288 4156 18294 4168
rect 10594 4088 10600 4140
rect 10652 4128 10658 4140
rect 12342 4128 12348 4140
rect 10652 4100 12348 4128
rect 10652 4088 10658 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13446 4128 13452 4140
rect 13311 4100 13452 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 14642 4128 14648 4140
rect 14047 4100 14648 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 14829 4131 14887 4137
rect 14829 4097 14841 4131
rect 14875 4128 14887 4131
rect 15286 4128 15292 4140
rect 14875 4100 15292 4128
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4128 15623 4131
rect 16114 4128 16120 4140
rect 15611 4100 16120 4128
rect 15611 4097 15623 4100
rect 15565 4091 15623 4097
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 17494 4128 17500 4140
rect 17455 4100 17500 4128
rect 17494 4088 17500 4100
rect 17552 4088 17558 4140
rect 17678 4128 17684 4140
rect 17639 4100 17684 4128
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 18782 4128 18788 4140
rect 17788 4100 18788 4128
rect 10091 4032 10180 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 12032 4032 12081 4060
rect 12032 4020 12038 4032
rect 12069 4029 12081 4032
rect 12115 4060 12127 4063
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 12115 4032 14749 4060
rect 12115 4029 12127 4032
rect 12069 4023 12127 4029
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4060 16083 4063
rect 17788 4060 17816 4100
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 19444 4137 19472 4168
rect 20806 4156 20812 4168
rect 20864 4156 20870 4208
rect 20898 4156 20904 4208
rect 20956 4196 20962 4208
rect 20956 4168 21001 4196
rect 20956 4156 20962 4168
rect 23474 4156 23480 4208
rect 23532 4196 23538 4208
rect 23532 4168 23888 4196
rect 23532 4156 23538 4168
rect 19429 4131 19487 4137
rect 19429 4097 19441 4131
rect 19475 4097 19487 4131
rect 19610 4128 19616 4140
rect 19571 4100 19616 4128
rect 19429 4091 19487 4097
rect 19334 4060 19340 4072
rect 16071 4032 17816 4060
rect 17880 4032 19340 4060
rect 16071 4029 16083 4032
rect 16025 4023 16083 4029
rect 5813 3995 5871 4001
rect 5813 3961 5825 3995
rect 5859 3992 5871 3995
rect 7742 3992 7748 4004
rect 5859 3964 7748 3992
rect 5859 3961 5871 3964
rect 5813 3955 5871 3961
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 11609 3995 11667 4001
rect 9640 3964 10732 3992
rect 9640 3952 9646 3964
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 2746 3896 4721 3924
rect 2409 3887 2467 3893
rect 4709 3893 4721 3896
rect 4755 3924 4767 3927
rect 4798 3924 4804 3936
rect 4755 3896 4804 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6822 3924 6828 3936
rect 6503 3896 6828 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 10704 3933 10732 3964
rect 11609 3961 11621 3995
rect 11655 3992 11667 3995
rect 12250 3992 12256 4004
rect 11655 3964 12256 3992
rect 11655 3961 11667 3964
rect 11609 3955 11667 3961
rect 12250 3952 12256 3964
rect 12308 3952 12314 4004
rect 12894 3952 12900 4004
rect 12952 3992 12958 4004
rect 15381 3995 15439 4001
rect 15381 3992 15393 3995
rect 12952 3964 15393 3992
rect 12952 3952 12958 3964
rect 15381 3961 15393 3964
rect 15427 3961 15439 3995
rect 15381 3955 15439 3961
rect 17494 3952 17500 4004
rect 17552 3992 17558 4004
rect 17880 3992 17908 4032
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 19444 4060 19472 4091
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 21174 4088 21180 4140
rect 21232 4128 21238 4140
rect 23860 4137 23888 4168
rect 27614 4156 27620 4208
rect 27672 4196 27678 4208
rect 28086 4199 28144 4205
rect 28086 4196 28098 4199
rect 27672 4168 28098 4196
rect 27672 4156 27678 4168
rect 28086 4165 28098 4168
rect 28132 4165 28144 4199
rect 28086 4159 28144 4165
rect 31478 4156 31484 4208
rect 31536 4196 31542 4208
rect 36814 4196 36820 4208
rect 31536 4168 36820 4196
rect 31536 4156 31542 4168
rect 36814 4156 36820 4168
rect 36872 4156 36878 4208
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21232 4100 21833 4128
rect 21232 4088 21238 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 23578 4131 23636 4137
rect 23578 4128 23590 4131
rect 21821 4091 21879 4097
rect 22020 4100 23590 4128
rect 19794 4060 19800 4072
rect 19444 4032 19800 4060
rect 19794 4020 19800 4032
rect 19852 4060 19858 4072
rect 20438 4060 20444 4072
rect 19852 4032 20444 4060
rect 19852 4020 19858 4032
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 20588 4032 20729 4060
rect 20588 4020 20594 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 17552 3964 17908 3992
rect 18325 3995 18383 4001
rect 17552 3952 17558 3964
rect 18325 3961 18337 3995
rect 18371 3992 18383 3995
rect 19518 3992 19524 4004
rect 18371 3964 19524 3992
rect 18371 3961 18383 3964
rect 18325 3955 18383 3961
rect 19518 3952 19524 3964
rect 19576 3952 19582 4004
rect 19613 3995 19671 4001
rect 19613 3961 19625 3995
rect 19659 3992 19671 3995
rect 20162 3992 20168 4004
rect 19659 3964 20168 3992
rect 19659 3961 19671 3964
rect 19613 3955 19671 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 20806 3952 20812 4004
rect 20864 3992 20870 4004
rect 22020 4001 22048 4100
rect 23578 4097 23590 4100
rect 23624 4097 23636 4131
rect 23578 4091 23636 4097
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 24670 4088 24676 4140
rect 24728 4128 24734 4140
rect 25406 4128 25412 4140
rect 24728 4100 25412 4128
rect 24728 4088 24734 4100
rect 25406 4088 25412 4100
rect 25464 4137 25470 4140
rect 25464 4131 25513 4137
rect 25464 4097 25467 4131
rect 25501 4097 25513 4131
rect 25590 4128 25596 4140
rect 25551 4100 25596 4128
rect 25464 4091 25513 4097
rect 25464 4088 25470 4091
rect 25590 4088 25596 4100
rect 25648 4088 25654 4140
rect 25682 4088 25688 4140
rect 25740 4131 25746 4140
rect 25869 4131 25927 4137
rect 25740 4103 25782 4131
rect 25740 4088 25746 4103
rect 25869 4097 25881 4131
rect 25915 4128 25927 4131
rect 26970 4128 26976 4140
rect 25915 4100 26976 4128
rect 25915 4097 25927 4100
rect 25869 4091 25927 4097
rect 26970 4088 26976 4100
rect 27028 4088 27034 4140
rect 28350 4128 28356 4140
rect 28311 4100 28356 4128
rect 28350 4088 28356 4100
rect 28408 4088 28414 4140
rect 28718 4088 28724 4140
rect 28776 4128 28782 4140
rect 28813 4131 28871 4137
rect 28813 4128 28825 4131
rect 28776 4100 28825 4128
rect 28776 4088 28782 4100
rect 28813 4097 28825 4100
rect 28859 4097 28871 4131
rect 28813 4091 28871 4097
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 30570 4131 30628 4137
rect 30570 4128 30582 4131
rect 29052 4100 30582 4128
rect 29052 4088 29058 4100
rect 30570 4097 30582 4100
rect 30616 4097 30628 4131
rect 30570 4091 30628 4097
rect 30837 4131 30895 4137
rect 30837 4097 30849 4131
rect 30883 4128 30895 4131
rect 31570 4128 31576 4140
rect 30883 4100 31576 4128
rect 30883 4097 30895 4100
rect 30837 4091 30895 4097
rect 31570 4088 31576 4100
rect 31628 4088 31634 4140
rect 34514 4088 34520 4140
rect 34572 4128 34578 4140
rect 34894 4131 34952 4137
rect 34894 4128 34906 4131
rect 34572 4100 34906 4128
rect 34572 4088 34578 4100
rect 34894 4097 34906 4100
rect 34940 4097 34952 4131
rect 35158 4128 35164 4140
rect 35119 4100 35164 4128
rect 34894 4091 34952 4097
rect 35158 4088 35164 4100
rect 35216 4088 35222 4140
rect 57974 4088 57980 4140
rect 58032 4128 58038 4140
rect 59817 4131 59875 4137
rect 59817 4128 59829 4131
rect 58032 4100 59829 4128
rect 58032 4088 58038 4100
rect 59817 4097 59829 4100
rect 59863 4097 59875 4131
rect 59817 4091 59875 4097
rect 25222 4060 25228 4072
rect 25183 4032 25228 4060
rect 25222 4020 25228 4032
rect 25280 4020 25286 4072
rect 59170 4020 59176 4072
rect 59228 4060 59234 4072
rect 61105 4063 61163 4069
rect 61105 4060 61117 4063
rect 59228 4032 61117 4060
rect 59228 4020 59234 4032
rect 61105 4029 61117 4032
rect 61151 4029 61163 4063
rect 61105 4023 61163 4029
rect 22005 3995 22063 4001
rect 20864 3964 21404 3992
rect 20864 3952 20870 3964
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 8260 3896 9689 3924
rect 8260 3884 8266 3896
rect 9677 3893 9689 3896
rect 9723 3893 9735 3927
rect 9677 3887 9735 3893
rect 10689 3927 10747 3933
rect 10689 3893 10701 3927
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 11848 3896 12357 3924
rect 11848 3884 11854 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 13081 3927 13139 3933
rect 13081 3893 13093 3927
rect 13127 3924 13139 3927
rect 13262 3924 13268 3936
rect 13127 3896 13268 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13688 3896 13829 3924
rect 13688 3884 13694 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 13817 3887 13875 3893
rect 14829 3927 14887 3933
rect 14829 3893 14841 3927
rect 14875 3924 14887 3927
rect 15010 3924 15016 3936
rect 14875 3896 15016 3924
rect 14875 3893 14887 3896
rect 14829 3887 14887 3893
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 18874 3924 18880 3936
rect 16899 3896 18880 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 18969 3927 19027 3933
rect 18969 3893 18981 3927
rect 19015 3924 19027 3927
rect 19334 3924 19340 3936
rect 19015 3896 19340 3924
rect 19015 3893 19027 3896
rect 18969 3887 19027 3893
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 20990 3884 20996 3936
rect 21048 3924 21054 3936
rect 21269 3927 21327 3933
rect 21269 3924 21281 3927
rect 21048 3896 21281 3924
rect 21048 3884 21054 3896
rect 21269 3893 21281 3896
rect 21315 3893 21327 3927
rect 21376 3924 21404 3964
rect 22005 3961 22017 3995
rect 22051 3961 22063 3995
rect 22005 3955 22063 3961
rect 57514 3952 57520 4004
rect 57572 3992 57578 4004
rect 58529 3995 58587 4001
rect 58529 3992 58541 3995
rect 57572 3964 58541 3992
rect 57572 3952 57578 3964
rect 58529 3961 58541 3964
rect 58575 3961 58587 3995
rect 58529 3955 58587 3961
rect 58618 3952 58624 4004
rect 58676 3992 58682 4004
rect 60461 3995 60519 4001
rect 60461 3992 60473 3995
rect 58676 3964 60473 3992
rect 58676 3952 58682 3964
rect 60461 3961 60473 3964
rect 60507 3961 60519 3995
rect 60461 3955 60519 3961
rect 22465 3927 22523 3933
rect 22465 3924 22477 3927
rect 21376 3896 22477 3924
rect 21269 3887 21327 3893
rect 22465 3893 22477 3896
rect 22511 3893 22523 3927
rect 24670 3924 24676 3936
rect 24631 3896 24676 3924
rect 22465 3887 22523 3893
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 56134 3884 56140 3936
rect 56192 3924 56198 3936
rect 56229 3927 56287 3933
rect 56229 3924 56241 3927
rect 56192 3896 56241 3924
rect 56192 3884 56198 3896
rect 56229 3893 56241 3896
rect 56275 3893 56287 3927
rect 56229 3887 56287 3893
rect 56318 3884 56324 3936
rect 56376 3924 56382 3936
rect 56873 3927 56931 3933
rect 56873 3924 56885 3927
rect 56376 3896 56885 3924
rect 56376 3884 56382 3896
rect 56873 3893 56885 3896
rect 56919 3893 56931 3927
rect 56873 3887 56931 3893
rect 56962 3884 56968 3936
rect 57020 3924 57026 3936
rect 57885 3927 57943 3933
rect 57885 3924 57897 3927
rect 57020 3896 57897 3924
rect 57020 3884 57026 3896
rect 57885 3893 57897 3896
rect 57931 3893 57943 3927
rect 57885 3887 57943 3893
rect 58066 3884 58072 3936
rect 58124 3924 58130 3936
rect 59173 3927 59231 3933
rect 59173 3924 59185 3927
rect 58124 3896 59185 3924
rect 58124 3884 58130 3896
rect 59173 3893 59185 3896
rect 59219 3893 59231 3927
rect 59173 3887 59231 3893
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2590 3720 2596 3732
rect 2363 3692 2596 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2590 3680 2596 3692
rect 2648 3680 2654 3732
rect 4706 3720 4712 3732
rect 2746 3692 4712 3720
rect 1854 3612 1860 3664
rect 1912 3652 1918 3664
rect 2746 3652 2774 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 6730 3720 6736 3732
rect 6691 3692 6736 3720
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 7432 3692 10609 3720
rect 7432 3680 7438 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 13078 3720 13084 3732
rect 10597 3683 10655 3689
rect 12084 3692 13084 3720
rect 3234 3652 3240 3664
rect 1912 3624 2774 3652
rect 3195 3624 3240 3652
rect 1912 3612 1918 3624
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 4798 3652 4804 3664
rect 4632 3624 4804 3652
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 4632 3593 4660 3624
rect 4798 3612 4804 3624
rect 4856 3652 4862 3664
rect 5350 3652 5356 3664
rect 4856 3624 5356 3652
rect 4856 3612 4862 3624
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 6362 3612 6368 3664
rect 6420 3652 6426 3664
rect 9674 3652 9680 3664
rect 6420 3624 9680 3652
rect 6420 3612 6426 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 9769 3655 9827 3661
rect 9769 3621 9781 3655
rect 9815 3621 9827 3655
rect 9769 3615 9827 3621
rect 1949 3587 2007 3593
rect 1949 3584 1961 3587
rect 1820 3556 1961 3584
rect 1820 3544 1826 3556
rect 1949 3553 1961 3556
rect 1995 3553 2007 3587
rect 1949 3547 2007 3553
rect 4617 3587 4675 3593
rect 4617 3553 4629 3587
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 4764 3556 4809 3584
rect 4764 3544 4770 3556
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7650 3584 7656 3596
rect 7156 3556 7656 3584
rect 7156 3544 7162 3556
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 7742 3544 7748 3596
rect 7800 3584 7806 3596
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 7800 3556 7849 3584
rect 7800 3544 7806 3556
rect 7837 3553 7849 3556
rect 7883 3584 7895 3587
rect 9306 3584 9312 3596
rect 7883 3556 9312 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9784 3584 9812 3615
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 12084 3652 12112 3692
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 14550 3720 14556 3732
rect 13587 3692 14556 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 17037 3723 17095 3729
rect 14700 3692 16988 3720
rect 14700 3680 14706 3692
rect 10008 3624 12112 3652
rect 10008 3612 10014 3624
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 12805 3655 12863 3661
rect 12805 3652 12817 3655
rect 12584 3624 12817 3652
rect 12584 3612 12590 3624
rect 12805 3621 12817 3624
rect 12851 3621 12863 3655
rect 16960 3652 16988 3692
rect 17037 3689 17049 3723
rect 17083 3720 17095 3723
rect 17862 3720 17868 3732
rect 17083 3692 17868 3720
rect 17083 3689 17095 3692
rect 17037 3683 17095 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 19610 3720 19616 3732
rect 18616 3692 19616 3720
rect 18506 3652 18512 3664
rect 16960 3624 18512 3652
rect 12805 3615 12863 3621
rect 18506 3612 18512 3624
rect 18564 3612 18570 3664
rect 12066 3584 12072 3596
rect 9784 3556 12072 3584
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 12768 3556 13369 3584
rect 12768 3544 12774 3556
rect 13357 3553 13369 3556
rect 13403 3584 13415 3587
rect 14182 3584 14188 3596
rect 13403 3556 14188 3584
rect 13403 3553 13415 3556
rect 13357 3547 13415 3553
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 15654 3584 15660 3596
rect 15615 3556 15660 3584
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 18616 3584 18644 3692
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 20073 3723 20131 3729
rect 20073 3720 20085 3723
rect 19944 3692 20085 3720
rect 19944 3680 19950 3692
rect 20073 3689 20085 3692
rect 20119 3689 20131 3723
rect 21174 3720 21180 3732
rect 21135 3692 21180 3720
rect 20073 3683 20131 3689
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 28994 3720 29000 3732
rect 28955 3692 29000 3720
rect 28994 3680 29000 3692
rect 29052 3680 29058 3732
rect 57790 3680 57796 3732
rect 57848 3720 57854 3732
rect 58066 3720 58072 3732
rect 57848 3692 58072 3720
rect 57848 3680 57854 3692
rect 58066 3680 58072 3692
rect 58124 3680 58130 3732
rect 18693 3655 18751 3661
rect 18693 3621 18705 3655
rect 18739 3652 18751 3655
rect 19337 3655 19395 3661
rect 19337 3652 19349 3655
rect 18739 3624 19349 3652
rect 18739 3621 18751 3624
rect 18693 3615 18751 3621
rect 19337 3621 19349 3624
rect 19383 3621 19395 3655
rect 19337 3615 19395 3621
rect 41138 3612 41144 3664
rect 41196 3652 41202 3664
rect 41785 3655 41843 3661
rect 41785 3652 41797 3655
rect 41196 3624 41797 3652
rect 41196 3612 41202 3624
rect 41785 3621 41797 3624
rect 41831 3621 41843 3655
rect 41785 3615 41843 3621
rect 56502 3612 56508 3664
rect 56560 3652 56566 3664
rect 57885 3655 57943 3661
rect 57885 3652 57897 3655
rect 56560 3624 57897 3652
rect 56560 3612 56566 3624
rect 57885 3621 57897 3624
rect 57931 3621 57943 3655
rect 57885 3615 57943 3621
rect 58342 3612 58348 3664
rect 58400 3652 58406 3664
rect 61105 3655 61163 3661
rect 61105 3652 61117 3655
rect 58400 3624 61117 3652
rect 58400 3612 58406 3624
rect 61105 3621 61117 3624
rect 61151 3621 61163 3655
rect 61105 3615 61163 3621
rect 16868 3556 18644 3584
rect 2130 3516 2136 3528
rect 2091 3488 2136 3516
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 3016 3488 3065 3516
rect 3016 3476 3022 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3142 3476 3148 3528
rect 3200 3516 3206 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 3200 3488 5365 3516
rect 3200 3476 3206 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5620 3519 5678 3525
rect 5620 3485 5632 3519
rect 5666 3485 5678 3519
rect 7558 3516 7564 3528
rect 7519 3488 7564 3516
rect 5620 3479 5678 3485
rect 1489 3451 1547 3457
rect 1489 3417 1501 3451
rect 1535 3448 1547 3451
rect 4525 3451 4583 3457
rect 1535 3420 4476 3448
rect 1535 3417 1547 3420
rect 1489 3411 1547 3417
rect 4154 3380 4160 3392
rect 4115 3352 4160 3380
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4448 3380 4476 3420
rect 4525 3417 4537 3451
rect 4571 3448 4583 3451
rect 4890 3448 4896 3460
rect 4571 3420 4896 3448
rect 4571 3417 4583 3420
rect 4525 3411 4583 3417
rect 4890 3408 4896 3420
rect 4948 3448 4954 3460
rect 5258 3448 5264 3460
rect 4948 3420 5264 3448
rect 4948 3408 4954 3420
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 5368 3448 5396 3479
rect 5534 3448 5540 3460
rect 5368 3420 5540 3448
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 5644 3448 5672 3479
rect 7558 3476 7564 3488
rect 7616 3516 7622 3528
rect 8202 3516 8208 3528
rect 7616 3488 8208 3516
rect 7616 3476 7622 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9950 3516 9956 3528
rect 9911 3488 9956 3516
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 11238 3516 11244 3528
rect 10376 3488 11008 3516
rect 11199 3488 11244 3516
rect 10376 3476 10382 3488
rect 5718 3448 5724 3460
rect 5644 3420 5724 3448
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 7834 3448 7840 3460
rect 6696 3420 7840 3448
rect 6696 3408 6702 3420
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 10581 3451 10639 3457
rect 9048 3420 10548 3448
rect 6270 3380 6276 3392
rect 4448 3352 6276 3380
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 7190 3380 7196 3392
rect 7151 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 9048 3389 9076 3420
rect 9033 3383 9091 3389
rect 9033 3349 9045 3383
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 10134 3380 10140 3392
rect 9732 3352 10140 3380
rect 9732 3340 9738 3352
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10410 3380 10416 3392
rect 10371 3352 10416 3380
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10520 3380 10548 3420
rect 10581 3417 10593 3451
rect 10627 3448 10639 3451
rect 10686 3448 10692 3460
rect 10627 3420 10692 3448
rect 10627 3417 10639 3420
rect 10581 3411 10639 3417
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 10778 3408 10784 3460
rect 10836 3448 10842 3460
rect 10980 3448 11008 3488
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 11882 3516 11888 3528
rect 11563 3488 11888 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 13262 3516 13268 3528
rect 12406 3488 13268 3516
rect 12406 3448 12434 3488
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 15746 3516 15752 3528
rect 14792 3488 15752 3516
rect 14792 3476 14798 3488
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 15924 3519 15982 3525
rect 15924 3485 15936 3519
rect 15970 3516 15982 3519
rect 16666 3516 16672 3528
rect 15970 3488 16672 3516
rect 15970 3485 15982 3488
rect 15924 3479 15982 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 10836 3420 10881 3448
rect 10980 3420 12434 3448
rect 10836 3408 10842 3420
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 12805 3451 12863 3457
rect 12805 3448 12817 3451
rect 12676 3420 12817 3448
rect 12676 3408 12682 3420
rect 12805 3417 12817 3420
rect 12851 3417 12863 3451
rect 12805 3411 12863 3417
rect 13998 3408 14004 3460
rect 14056 3448 14062 3460
rect 16868 3448 16896 3556
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 19797 3587 19855 3593
rect 19797 3584 19809 3587
rect 19484 3556 19809 3584
rect 19484 3544 19490 3556
rect 19797 3553 19809 3556
rect 19843 3553 19855 3587
rect 19797 3547 19855 3553
rect 19889 3587 19947 3593
rect 19889 3553 19901 3587
rect 19935 3584 19947 3587
rect 19978 3584 19984 3596
rect 19935 3556 19984 3584
rect 19935 3553 19947 3556
rect 19889 3547 19947 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20254 3544 20260 3596
rect 20312 3584 20318 3596
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20312 3556 20821 3584
rect 20312 3544 20318 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 28258 3544 28264 3596
rect 28316 3584 28322 3596
rect 28316 3556 28672 3584
rect 28316 3544 28322 3556
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3516 18567 3519
rect 20162 3516 20168 3528
rect 18555 3488 20168 3516
rect 18555 3485 18567 3488
rect 18509 3479 18567 3485
rect 14056 3420 16896 3448
rect 14056 3408 14062 3420
rect 11330 3380 11336 3392
rect 10520 3352 11336 3380
rect 11330 3340 11336 3352
rect 11388 3340 11394 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 11790 3380 11796 3392
rect 11664 3352 11796 3380
rect 11664 3340 11670 3352
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 13078 3340 13084 3392
rect 13136 3380 13142 3392
rect 13265 3383 13323 3389
rect 13265 3380 13277 3383
rect 13136 3352 13277 3380
rect 13136 3340 13142 3352
rect 13265 3349 13277 3352
rect 13311 3380 13323 3383
rect 13722 3380 13728 3392
rect 13311 3352 13728 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 13722 3340 13728 3352
rect 13780 3380 13786 3392
rect 14550 3380 14556 3392
rect 13780 3352 14556 3380
rect 13780 3340 13786 3352
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 14700 3352 14745 3380
rect 14700 3340 14706 3352
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17954 3380 17960 3392
rect 17276 3352 17960 3380
rect 17276 3340 17282 3352
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18064 3380 18092 3479
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 20990 3516 20996 3528
rect 20951 3488 20996 3516
rect 20990 3476 20996 3488
rect 21048 3476 21054 3528
rect 21818 3476 21824 3528
rect 21876 3516 21882 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21876 3488 21925 3516
rect 21876 3476 21882 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 22646 3476 22652 3528
rect 22704 3516 22710 3528
rect 22741 3519 22799 3525
rect 22741 3516 22753 3519
rect 22704 3488 22753 3516
rect 22704 3476 22710 3488
rect 22741 3485 22753 3488
rect 22787 3485 22799 3519
rect 22741 3479 22799 3485
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 23569 3519 23627 3525
rect 23569 3516 23581 3519
rect 23532 3488 23581 3516
rect 23532 3476 23538 3488
rect 23569 3485 23581 3488
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 24360 3488 24409 3516
rect 24360 3476 24366 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 25130 3476 25136 3528
rect 25188 3516 25194 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 25188 3488 25237 3516
rect 25188 3476 25194 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25958 3476 25964 3528
rect 26016 3516 26022 3528
rect 26053 3519 26111 3525
rect 26053 3516 26065 3519
rect 26016 3488 26065 3516
rect 26016 3476 26022 3488
rect 26053 3485 26065 3488
rect 26099 3485 26111 3519
rect 26053 3479 26111 3485
rect 26786 3476 26792 3528
rect 26844 3516 26850 3528
rect 26881 3519 26939 3525
rect 26881 3516 26893 3519
rect 26844 3488 26893 3516
rect 26844 3476 26850 3488
rect 26881 3485 26893 3488
rect 26927 3485 26939 3519
rect 26881 3479 26939 3485
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 27709 3519 27767 3525
rect 27709 3516 27721 3519
rect 27672 3488 27721 3516
rect 27672 3476 27678 3488
rect 27709 3485 27721 3488
rect 27755 3485 27767 3519
rect 27709 3479 27767 3485
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 28353 3519 28411 3525
rect 28353 3516 28365 3519
rect 27948 3488 28365 3516
rect 27948 3476 27954 3488
rect 28353 3485 28365 3488
rect 28399 3485 28411 3519
rect 28534 3516 28540 3528
rect 28495 3488 28540 3516
rect 28353 3479 28411 3485
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 28644 3525 28672 3556
rect 55766 3544 55772 3596
rect 55824 3584 55830 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 55824 3556 56609 3584
rect 55824 3544 55830 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 56778 3544 56784 3596
rect 56836 3584 56842 3596
rect 58529 3587 58587 3593
rect 58529 3584 58541 3587
rect 56836 3556 58541 3584
rect 56836 3544 56842 3556
rect 58529 3553 58541 3556
rect 58575 3553 58587 3587
rect 58529 3547 58587 3553
rect 58986 3544 58992 3596
rect 59044 3584 59050 3596
rect 61749 3587 61807 3593
rect 61749 3584 61761 3587
rect 59044 3556 61761 3584
rect 59044 3544 59050 3556
rect 61749 3553 61761 3556
rect 61795 3553 61807 3587
rect 61749 3547 61807 3553
rect 28629 3519 28687 3525
rect 28629 3485 28641 3519
rect 28675 3485 28687 3519
rect 28629 3479 28687 3485
rect 28718 3476 28724 3528
rect 28776 3516 28782 3528
rect 28776 3488 28821 3516
rect 28776 3476 28782 3488
rect 29822 3476 29828 3528
rect 29880 3516 29886 3528
rect 29917 3519 29975 3525
rect 29917 3516 29929 3519
rect 29880 3488 29929 3516
rect 29880 3476 29886 3488
rect 29917 3485 29929 3488
rect 29963 3485 29975 3519
rect 29917 3479 29975 3485
rect 30650 3476 30656 3528
rect 30708 3516 30714 3528
rect 30745 3519 30803 3525
rect 30745 3516 30757 3519
rect 30708 3488 30757 3516
rect 30708 3476 30714 3488
rect 30745 3485 30757 3488
rect 30791 3485 30803 3519
rect 30745 3479 30803 3485
rect 31478 3476 31484 3528
rect 31536 3516 31542 3528
rect 31573 3519 31631 3525
rect 31573 3516 31585 3519
rect 31536 3488 31585 3516
rect 31536 3476 31542 3488
rect 31573 3485 31585 3488
rect 31619 3485 31631 3519
rect 31573 3479 31631 3485
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 32401 3519 32459 3525
rect 32401 3516 32413 3519
rect 32364 3488 32413 3516
rect 32364 3476 32370 3488
rect 32401 3485 32413 3488
rect 32447 3485 32459 3519
rect 32401 3479 32459 3485
rect 33134 3476 33140 3528
rect 33192 3516 33198 3528
rect 33229 3519 33287 3525
rect 33229 3516 33241 3519
rect 33192 3488 33241 3516
rect 33192 3476 33198 3488
rect 33229 3485 33241 3488
rect 33275 3485 33287 3519
rect 33229 3479 33287 3485
rect 39206 3476 39212 3528
rect 39264 3516 39270 3528
rect 39853 3519 39911 3525
rect 39853 3516 39865 3519
rect 39264 3488 39865 3516
rect 39264 3476 39270 3488
rect 39853 3485 39865 3488
rect 39899 3485 39911 3519
rect 39853 3479 39911 3485
rect 40034 3476 40040 3528
rect 40092 3516 40098 3528
rect 40497 3519 40555 3525
rect 40497 3516 40509 3519
rect 40092 3488 40509 3516
rect 40092 3476 40098 3488
rect 40497 3485 40509 3488
rect 40543 3485 40555 3519
rect 40497 3479 40555 3485
rect 40862 3476 40868 3528
rect 40920 3516 40926 3528
rect 41141 3519 41199 3525
rect 41141 3516 41153 3519
rect 40920 3488 41153 3516
rect 40920 3476 40926 3488
rect 41141 3485 41153 3488
rect 41187 3485 41199 3519
rect 41141 3479 41199 3485
rect 42518 3476 42524 3528
rect 42576 3516 42582 3528
rect 42613 3519 42671 3525
rect 42613 3516 42625 3519
rect 42576 3488 42625 3516
rect 42576 3476 42582 3488
rect 42613 3485 42625 3488
rect 42659 3485 42671 3519
rect 42613 3479 42671 3485
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 43128 3488 43269 3516
rect 43128 3476 43134 3488
rect 43257 3485 43269 3488
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 45002 3476 45008 3528
rect 45060 3516 45066 3528
rect 45097 3519 45155 3525
rect 45097 3516 45109 3519
rect 45060 3488 45109 3516
rect 45060 3476 45066 3488
rect 45097 3485 45109 3488
rect 45143 3485 45155 3519
rect 45097 3479 45155 3485
rect 45278 3476 45284 3528
rect 45336 3516 45342 3528
rect 45741 3519 45799 3525
rect 45741 3516 45753 3519
rect 45336 3488 45753 3516
rect 45336 3476 45342 3488
rect 45741 3485 45753 3488
rect 45787 3485 45799 3519
rect 45741 3479 45799 3485
rect 46106 3476 46112 3528
rect 46164 3516 46170 3528
rect 46385 3519 46443 3525
rect 46385 3516 46397 3519
rect 46164 3488 46397 3516
rect 46164 3476 46170 3488
rect 46385 3485 46397 3488
rect 46431 3485 46443 3519
rect 46385 3479 46443 3485
rect 46934 3476 46940 3528
rect 46992 3516 46998 3528
rect 47029 3519 47087 3525
rect 47029 3516 47041 3519
rect 46992 3488 47041 3516
rect 46992 3476 46998 3488
rect 47029 3485 47041 3488
rect 47075 3485 47087 3519
rect 47029 3479 47087 3485
rect 47762 3476 47768 3528
rect 47820 3516 47826 3528
rect 47857 3519 47915 3525
rect 47857 3516 47869 3519
rect 47820 3488 47869 3516
rect 47820 3476 47826 3488
rect 47857 3485 47869 3488
rect 47903 3485 47915 3519
rect 47857 3479 47915 3485
rect 48866 3476 48872 3528
rect 48924 3516 48930 3528
rect 48961 3519 49019 3525
rect 48961 3516 48973 3519
rect 48924 3488 48973 3516
rect 48924 3476 48930 3488
rect 48961 3485 48973 3488
rect 49007 3485 49019 3519
rect 48961 3479 49019 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50341 3519 50399 3525
rect 50341 3516 50353 3519
rect 50212 3488 50353 3516
rect 50212 3476 50218 3488
rect 50341 3485 50353 3488
rect 50387 3485 50399 3519
rect 50341 3479 50399 3485
rect 50798 3476 50804 3528
rect 50856 3516 50862 3528
rect 50985 3519 51043 3525
rect 50985 3516 50997 3519
rect 50856 3488 50997 3516
rect 50856 3476 50862 3488
rect 50985 3485 50997 3488
rect 51031 3485 51043 3519
rect 50985 3479 51043 3485
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 51629 3519 51687 3525
rect 51629 3516 51641 3519
rect 51408 3488 51641 3516
rect 51408 3476 51414 3488
rect 51629 3485 51641 3488
rect 51675 3485 51687 3519
rect 51629 3479 51687 3485
rect 52730 3476 52736 3528
rect 52788 3516 52794 3528
rect 52825 3519 52883 3525
rect 52825 3516 52837 3519
rect 52788 3488 52837 3516
rect 52788 3476 52794 3488
rect 52825 3485 52837 3488
rect 52871 3485 52883 3519
rect 52825 3479 52883 3485
rect 53006 3476 53012 3528
rect 53064 3516 53070 3528
rect 53469 3519 53527 3525
rect 53469 3516 53481 3519
rect 53064 3488 53481 3516
rect 53064 3476 53070 3488
rect 53469 3485 53481 3488
rect 53515 3485 53527 3519
rect 53469 3479 53527 3485
rect 54662 3476 54668 3528
rect 54720 3516 54726 3528
rect 55309 3519 55367 3525
rect 55309 3516 55321 3519
rect 54720 3488 55321 3516
rect 54720 3476 54726 3488
rect 55309 3485 55321 3488
rect 55355 3485 55367 3519
rect 55309 3479 55367 3485
rect 55490 3476 55496 3528
rect 55548 3516 55554 3528
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 55548 3488 55965 3516
rect 55548 3476 55554 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 55953 3479 56011 3485
rect 56226 3476 56232 3528
rect 56284 3516 56290 3528
rect 57241 3519 57299 3525
rect 57241 3516 57253 3519
rect 56284 3488 57253 3516
rect 56284 3476 56290 3488
rect 57241 3485 57253 3488
rect 57287 3485 57299 3519
rect 57241 3479 57299 3485
rect 57330 3476 57336 3528
rect 57388 3516 57394 3528
rect 59173 3519 59231 3525
rect 59173 3516 59185 3519
rect 57388 3488 59185 3516
rect 57388 3476 57394 3488
rect 59173 3485 59185 3488
rect 59219 3485 59231 3519
rect 60458 3516 60464 3528
rect 60419 3488 60464 3516
rect 59173 3479 59231 3485
rect 60458 3476 60464 3488
rect 60516 3476 60522 3528
rect 68094 3516 68100 3528
rect 68055 3488 68100 3516
rect 68094 3476 68100 3488
rect 68152 3476 68158 3528
rect 19334 3448 19340 3460
rect 19295 3420 19340 3448
rect 19334 3408 19340 3420
rect 19392 3408 19398 3460
rect 19426 3380 19432 3392
rect 18064 3352 19432 3380
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 4672 3148 5457 3176
rect 4672 3136 4678 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 7190 3176 7196 3188
rect 5445 3139 5503 3145
rect 5644 3148 7196 3176
rect 4154 3108 4160 3120
rect 2746 3080 4160 3108
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3040 1547 3043
rect 2133 3043 2191 3049
rect 2133 3040 2145 3043
rect 1535 3012 2145 3040
rect 1535 3009 1547 3012
rect 1489 3003 1547 3009
rect 2133 3009 2145 3012
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2746 3040 2774 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 2363 3012 2774 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 5644 3049 5672 3148
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7708 3148 7757 3176
rect 7708 3136 7714 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 11422 3176 11428 3188
rect 7892 3148 11428 3176
rect 7892 3136 7898 3148
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12158 3176 12164 3188
rect 11931 3148 12164 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 13372 3148 14053 3176
rect 6380 3080 8248 3108
rect 6380 3049 6408 3080
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3200 3012 3433 3040
rect 3200 3000 3206 3012
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 3677 3043 3735 3049
rect 3677 3040 3689 3043
rect 3421 3003 3479 3009
rect 3528 3012 3689 3040
rect 1762 2932 1768 2984
rect 1820 2972 1826 2984
rect 2501 2975 2559 2981
rect 2501 2972 2513 2975
rect 1820 2944 2513 2972
rect 1820 2932 1826 2944
rect 2501 2941 2513 2944
rect 2547 2972 2559 2975
rect 2590 2972 2596 2984
rect 2547 2944 2596 2972
rect 2547 2941 2559 2944
rect 2501 2935 2559 2941
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 3528 2972 3556 3012
rect 3677 3009 3689 3012
rect 3723 3009 3735 3043
rect 3677 3003 3735 3009
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3009 5687 3043
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5629 3003 5687 3009
rect 5736 3012 6377 3040
rect 2746 2944 3556 2972
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 2746 2904 2774 2944
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 5736 2972 5764 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 8220 3049 8248 3080
rect 10226 3068 10232 3120
rect 10284 3108 10290 3120
rect 10873 3111 10931 3117
rect 10873 3108 10885 3111
rect 10284 3080 10885 3108
rect 10284 3068 10290 3080
rect 10873 3077 10885 3080
rect 10919 3108 10931 3111
rect 11606 3108 11612 3120
rect 10919 3080 11612 3108
rect 10919 3077 10931 3080
rect 10873 3071 10931 3077
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 12618 3068 12624 3120
rect 12676 3108 12682 3120
rect 13372 3117 13400 3148
rect 13357 3111 13415 3117
rect 13357 3108 13369 3111
rect 12676 3080 13369 3108
rect 12676 3068 12682 3080
rect 13357 3077 13369 3080
rect 13403 3077 13415 3111
rect 13357 3071 13415 3077
rect 13722 3068 13728 3120
rect 13780 3068 13786 3120
rect 6621 3043 6679 3049
rect 6621 3040 6633 3043
rect 6512 3012 6633 3040
rect 6512 3000 6518 3012
rect 6621 3009 6633 3012
rect 6667 3009 6679 3043
rect 6621 3003 6679 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 8478 3049 8484 3052
rect 8472 3040 8484 3049
rect 8439 3012 8484 3040
rect 8472 3003 8484 3012
rect 8478 3000 8484 3003
rect 8536 3000 8542 3052
rect 12250 3040 12256 3052
rect 12176 3012 12256 3040
rect 5592 2944 5764 2972
rect 5813 2975 5871 2981
rect 5592 2932 5598 2944
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 8312 2972 8340 3000
rect 12176 2984 12204 3012
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12492 3012 12725 3040
rect 12492 3000 12498 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 13740 3040 13768 3068
rect 13814 3043 13872 3049
rect 13814 3040 13826 3043
rect 13740 3012 13826 3040
rect 12713 3003 12771 3009
rect 13814 3009 13826 3012
rect 13860 3009 13872 3043
rect 14025 3040 14053 3148
rect 14090 3136 14096 3188
rect 14148 3176 14154 3188
rect 16761 3179 16819 3185
rect 16761 3176 16773 3179
rect 14148 3148 16773 3176
rect 14148 3136 14154 3148
rect 16761 3145 16773 3148
rect 16807 3145 16819 3179
rect 16761 3139 16819 3145
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 20956 3148 21833 3176
rect 20956 3136 20962 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 55950 3136 55956 3188
rect 56008 3176 56014 3188
rect 58066 3176 58072 3188
rect 56008 3148 58072 3176
rect 56008 3136 56014 3148
rect 58066 3136 58072 3148
rect 58124 3136 58130 3188
rect 14550 3068 14556 3120
rect 14608 3068 14614 3120
rect 15930 3068 15936 3120
rect 15988 3108 15994 3120
rect 15988 3080 17448 3108
rect 15988 3068 15994 3080
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 14025 3012 14473 3040
rect 13814 3003 13872 3009
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 14568 3040 14596 3068
rect 14737 3043 14795 3049
rect 14737 3040 14749 3043
rect 14568 3012 14749 3040
rect 14461 3003 14519 3009
rect 14737 3009 14749 3012
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3040 15807 3043
rect 16758 3040 16764 3052
rect 15795 3012 16764 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17310 3040 17316 3052
rect 16991 3012 17316 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17420 3049 17448 3080
rect 57698 3068 57704 3120
rect 57756 3108 57762 3120
rect 60458 3108 60464 3120
rect 57756 3080 60464 3108
rect 57756 3068 57762 3080
rect 60458 3068 60464 3080
rect 60516 3068 60522 3120
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 20162 3000 20168 3052
rect 20220 3040 20226 3052
rect 21726 3040 21732 3052
rect 20220 3012 21732 3040
rect 20220 3000 20226 3012
rect 21726 3000 21732 3012
rect 21784 3000 21790 3052
rect 58158 3000 58164 3052
rect 58216 3040 58222 3052
rect 61105 3043 61163 3049
rect 61105 3040 61117 3043
rect 58216 3012 61117 3040
rect 58216 3000 58222 3012
rect 61105 3009 61117 3012
rect 61151 3009 61163 3043
rect 61105 3003 61163 3009
rect 10594 2972 10600 2984
rect 5859 2944 5948 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 4798 2904 4804 2916
rect 1719 2876 2774 2904
rect 4759 2876 4804 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 4798 2864 4804 2876
rect 4856 2864 4862 2916
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 5920 2836 5948 2944
rect 7392 2944 8340 2972
rect 10555 2944 10600 2972
rect 7392 2836 7420 2944
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 12158 2972 12164 2984
rect 12071 2944 12164 2972
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 13633 2975 13691 2981
rect 13633 2941 13645 2975
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 11882 2864 11888 2916
rect 11940 2904 11946 2916
rect 12250 2904 12256 2916
rect 11940 2876 12256 2904
rect 11940 2864 11946 2876
rect 12250 2864 12256 2876
rect 12308 2864 12314 2916
rect 12526 2864 12532 2916
rect 12584 2904 12590 2916
rect 13446 2904 13452 2916
rect 12584 2876 13452 2904
rect 12584 2864 12590 2876
rect 13446 2864 13452 2876
rect 13504 2904 13510 2916
rect 13648 2904 13676 2935
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 18693 2975 18751 2981
rect 14608 2944 14653 2972
rect 14608 2932 14614 2944
rect 18693 2941 18705 2975
rect 18739 2972 18751 2975
rect 20254 2972 20260 2984
rect 18739 2944 20260 2972
rect 18739 2941 18751 2944
rect 18693 2935 18751 2941
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 20625 2975 20683 2981
rect 20625 2941 20637 2975
rect 20671 2972 20683 2975
rect 21266 2972 21272 2984
rect 20671 2944 21272 2972
rect 20671 2941 20683 2944
rect 20625 2935 20683 2941
rect 21266 2932 21272 2944
rect 21324 2932 21330 2984
rect 37274 2932 37280 2984
rect 37332 2972 37338 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37332 2944 37933 2972
rect 37332 2932 37338 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 44726 2932 44732 2984
rect 44784 2972 44790 2984
rect 45649 2975 45707 2981
rect 45649 2972 45661 2975
rect 44784 2944 45661 2972
rect 44784 2932 44790 2944
rect 45649 2941 45661 2944
rect 45695 2941 45707 2975
rect 45649 2935 45707 2941
rect 48590 2932 48596 2984
rect 48648 2972 48654 2984
rect 49513 2975 49571 2981
rect 49513 2972 49525 2975
rect 48648 2944 49525 2972
rect 48648 2932 48654 2944
rect 49513 2941 49525 2944
rect 49559 2941 49571 2975
rect 49513 2935 49571 2941
rect 52454 2932 52460 2984
rect 52512 2972 52518 2984
rect 53377 2975 53435 2981
rect 53377 2972 53389 2975
rect 52512 2944 53389 2972
rect 52512 2932 52518 2944
rect 53377 2941 53389 2944
rect 53423 2941 53435 2975
rect 53377 2935 53435 2941
rect 53558 2932 53564 2984
rect 53616 2972 53622 2984
rect 55214 2972 55220 2984
rect 53616 2944 55220 2972
rect 53616 2932 53622 2944
rect 55214 2932 55220 2944
rect 55272 2932 55278 2984
rect 56686 2932 56692 2984
rect 56744 2972 56750 2984
rect 56744 2944 58204 2972
rect 56744 2932 56750 2944
rect 13504 2876 13676 2904
rect 13740 2876 14228 2904
rect 13504 2864 13510 2876
rect 2648 2808 7420 2836
rect 2648 2796 2654 2808
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 9585 2839 9643 2845
rect 9585 2836 9597 2839
rect 8444 2808 9597 2836
rect 8444 2796 8450 2808
rect 9585 2805 9597 2808
rect 9631 2805 9643 2839
rect 9585 2799 9643 2805
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 13740 2845 13768 2876
rect 14200 2848 14228 2876
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15565 2907 15623 2913
rect 15565 2904 15577 2907
rect 14884 2876 15577 2904
rect 14884 2864 14890 2876
rect 15565 2873 15577 2876
rect 15611 2873 15623 2907
rect 15565 2867 15623 2873
rect 15654 2864 15660 2916
rect 15712 2904 15718 2916
rect 17589 2907 17647 2913
rect 17589 2904 17601 2907
rect 15712 2876 17601 2904
rect 15712 2864 15718 2876
rect 17589 2873 17601 2876
rect 17635 2873 17647 2907
rect 17589 2867 17647 2873
rect 19337 2907 19395 2913
rect 19337 2873 19349 2907
rect 19383 2904 19395 2907
rect 20438 2904 20444 2916
rect 19383 2876 20444 2904
rect 19383 2873 19395 2876
rect 19337 2867 19395 2873
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 38378 2864 38384 2916
rect 38436 2904 38442 2916
rect 39209 2907 39267 2913
rect 39209 2904 39221 2907
rect 38436 2876 39221 2904
rect 38436 2864 38442 2876
rect 39209 2873 39221 2876
rect 39255 2873 39267 2907
rect 39209 2867 39267 2873
rect 39758 2864 39764 2916
rect 39816 2904 39822 2916
rect 40497 2907 40555 2913
rect 40497 2904 40509 2907
rect 39816 2876 40509 2904
rect 39816 2864 39822 2876
rect 40497 2873 40509 2876
rect 40543 2873 40555 2907
rect 40497 2867 40555 2873
rect 42242 2864 42248 2916
rect 42300 2904 42306 2916
rect 43073 2907 43131 2913
rect 43073 2904 43085 2907
rect 42300 2876 43085 2904
rect 42300 2864 42306 2876
rect 43073 2873 43085 2876
rect 43119 2873 43131 2907
rect 43073 2867 43131 2873
rect 43622 2864 43628 2916
rect 43680 2904 43686 2916
rect 44361 2907 44419 2913
rect 44361 2904 44373 2907
rect 43680 2876 44373 2904
rect 43680 2864 43686 2876
rect 44361 2873 44373 2876
rect 44407 2873 44419 2907
rect 44361 2867 44419 2873
rect 47486 2864 47492 2916
rect 47544 2904 47550 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 47544 2876 48237 2904
rect 47544 2864 47550 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 49418 2864 49424 2916
rect 49476 2904 49482 2916
rect 50157 2907 50215 2913
rect 50157 2904 50169 2907
rect 49476 2876 50169 2904
rect 49476 2864 49482 2876
rect 50157 2873 50169 2876
rect 50203 2873 50215 2907
rect 50157 2867 50215 2873
rect 50614 2864 50620 2916
rect 50672 2904 50678 2916
rect 51445 2907 51503 2913
rect 51445 2904 51457 2907
rect 50672 2876 51457 2904
rect 50672 2864 50678 2876
rect 51445 2873 51457 2876
rect 51491 2873 51503 2907
rect 51445 2867 51503 2873
rect 53282 2864 53288 2916
rect 53340 2904 53346 2916
rect 54021 2907 54079 2913
rect 54021 2904 54033 2907
rect 53340 2876 54033 2904
rect 53340 2864 53346 2876
rect 54021 2873 54033 2876
rect 54067 2873 54079 2907
rect 54021 2867 54079 2873
rect 54386 2864 54392 2916
rect 54444 2904 54450 2916
rect 55309 2907 55367 2913
rect 55309 2904 55321 2907
rect 54444 2876 55321 2904
rect 54444 2864 54450 2876
rect 55309 2873 55321 2876
rect 55355 2873 55367 2907
rect 55309 2867 55367 2873
rect 55674 2864 55680 2916
rect 55732 2904 55738 2916
rect 56597 2907 56655 2913
rect 56597 2904 56609 2907
rect 55732 2876 56609 2904
rect 55732 2864 55738 2876
rect 56597 2873 56609 2876
rect 56643 2873 56655 2907
rect 56597 2867 56655 2873
rect 57054 2864 57060 2916
rect 57112 2904 57118 2916
rect 58176 2904 58204 2944
rect 58434 2932 58440 2984
rect 58492 2972 58498 2984
rect 61749 2975 61807 2981
rect 61749 2972 61761 2975
rect 58492 2944 61761 2972
rect 58492 2932 58498 2944
rect 61749 2941 61761 2944
rect 61795 2941 61807 2975
rect 61749 2935 61807 2941
rect 58529 2907 58587 2913
rect 58529 2904 58541 2907
rect 57112 2876 58020 2904
rect 58176 2876 58541 2904
rect 57112 2864 57118 2876
rect 12345 2839 12403 2845
rect 12345 2836 12357 2839
rect 12032 2808 12357 2836
rect 12032 2796 12038 2808
rect 12345 2805 12357 2808
rect 12391 2805 12403 2839
rect 12345 2799 12403 2805
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2805 13783 2839
rect 13998 2836 14004 2848
rect 13959 2808 14004 2836
rect 13725 2799 13783 2805
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 14240 2808 14473 2836
rect 14240 2796 14246 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14918 2836 14924 2848
rect 14879 2808 14924 2836
rect 14461 2799 14519 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 15838 2796 15844 2848
rect 15896 2836 15902 2848
rect 18690 2836 18696 2848
rect 15896 2808 18696 2836
rect 15896 2796 15902 2808
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 19981 2839 20039 2845
rect 19981 2805 19993 2839
rect 20027 2836 20039 2839
rect 20714 2836 20720 2848
rect 20027 2808 20720 2836
rect 20027 2805 20039 2808
rect 19981 2799 20039 2805
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 21269 2839 21327 2845
rect 21269 2805 21281 2839
rect 21315 2836 21327 2839
rect 21542 2836 21548 2848
rect 21315 2808 21548 2836
rect 21315 2805 21327 2808
rect 21269 2799 21327 2805
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 22557 2839 22615 2845
rect 22557 2805 22569 2839
rect 22603 2836 22615 2839
rect 22922 2836 22928 2848
rect 22603 2808 22928 2836
rect 22603 2805 22615 2808
rect 22557 2799 22615 2805
rect 22922 2796 22928 2808
rect 22980 2796 22986 2848
rect 23201 2839 23259 2845
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 23750 2836 23756 2848
rect 23247 2808 23756 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 23750 2796 23756 2808
rect 23808 2796 23814 2848
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 24026 2836 24032 2848
rect 23891 2808 24032 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 24854 2836 24860 2848
rect 24535 2808 24860 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2836 25191 2839
rect 25682 2836 25688 2848
rect 25179 2808 25688 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 25682 2796 25688 2808
rect 25740 2796 25746 2848
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 26234 2836 26240 2848
rect 25823 2808 26240 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 26234 2796 26240 2808
rect 26292 2796 26298 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 27062 2836 27068 2848
rect 26467 2808 27068 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 27062 2796 27068 2808
rect 27120 2796 27126 2848
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2836 27767 2839
rect 28166 2836 28172 2848
rect 27755 2808 28172 2836
rect 27755 2805 27767 2808
rect 27709 2799 27767 2805
rect 28166 2796 28172 2808
rect 28224 2796 28230 2848
rect 28353 2839 28411 2845
rect 28353 2805 28365 2839
rect 28399 2836 28411 2839
rect 28718 2836 28724 2848
rect 28399 2808 28724 2836
rect 28399 2805 28411 2808
rect 28353 2799 28411 2805
rect 28718 2796 28724 2808
rect 28776 2796 28782 2848
rect 28997 2839 29055 2845
rect 28997 2805 29009 2839
rect 29043 2836 29055 2839
rect 29270 2836 29276 2848
rect 29043 2808 29276 2836
rect 29043 2805 29055 2808
rect 28997 2799 29055 2805
rect 29270 2796 29276 2808
rect 29328 2796 29334 2848
rect 29641 2839 29699 2845
rect 29641 2805 29653 2839
rect 29687 2836 29699 2839
rect 30098 2836 30104 2848
rect 29687 2808 30104 2836
rect 29687 2805 29699 2808
rect 29641 2799 29699 2805
rect 30098 2796 30104 2808
rect 30156 2796 30162 2848
rect 30285 2839 30343 2845
rect 30285 2805 30297 2839
rect 30331 2836 30343 2839
rect 30374 2836 30380 2848
rect 30331 2808 30380 2836
rect 30331 2805 30343 2808
rect 30285 2799 30343 2805
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 30929 2839 30987 2845
rect 30929 2805 30941 2839
rect 30975 2836 30987 2839
rect 31202 2836 31208 2848
rect 30975 2808 31208 2836
rect 30975 2805 30987 2808
rect 30929 2799 30987 2805
rect 31202 2796 31208 2808
rect 31260 2796 31266 2848
rect 31573 2839 31631 2845
rect 31573 2805 31585 2839
rect 31619 2836 31631 2839
rect 32030 2836 32036 2848
rect 31619 2808 32036 2836
rect 31619 2805 31631 2808
rect 31573 2799 31631 2805
rect 32030 2796 32036 2808
rect 32088 2796 32094 2848
rect 32858 2836 32864 2848
rect 32819 2808 32864 2836
rect 32858 2796 32864 2808
rect 32916 2796 32922 2848
rect 33505 2839 33563 2845
rect 33505 2805 33517 2839
rect 33551 2836 33563 2839
rect 33686 2836 33692 2848
rect 33551 2808 33692 2836
rect 33551 2805 33563 2808
rect 33505 2799 33563 2805
rect 33686 2796 33692 2808
rect 33744 2796 33750 2848
rect 34149 2839 34207 2845
rect 34149 2805 34161 2839
rect 34195 2836 34207 2839
rect 34238 2836 34244 2848
rect 34195 2808 34244 2836
rect 34195 2805 34207 2808
rect 34149 2799 34207 2805
rect 34238 2796 34244 2808
rect 34296 2796 34302 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34609 2839 34667 2845
rect 34609 2836 34621 2839
rect 34572 2808 34621 2836
rect 34572 2796 34578 2808
rect 34609 2805 34621 2808
rect 34655 2805 34667 2839
rect 34609 2799 34667 2805
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35437 2839 35495 2845
rect 35437 2836 35449 2839
rect 35400 2808 35449 2836
rect 35400 2796 35406 2808
rect 35437 2805 35449 2808
rect 35483 2805 35495 2839
rect 35437 2799 35495 2805
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 36265 2839 36323 2845
rect 36265 2836 36277 2839
rect 36228 2808 36277 2836
rect 36228 2796 36234 2808
rect 36265 2805 36277 2808
rect 36311 2805 36323 2839
rect 36265 2799 36323 2805
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36780 2808 37289 2836
rect 36780 2796 36786 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37826 2796 37832 2848
rect 37884 2836 37890 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 37884 2808 38577 2836
rect 37884 2796 37890 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 38930 2796 38936 2848
rect 38988 2836 38994 2848
rect 39853 2839 39911 2845
rect 39853 2836 39865 2839
rect 38988 2808 39865 2836
rect 38988 2796 38994 2808
rect 39853 2805 39865 2808
rect 39899 2805 39911 2839
rect 39853 2799 39911 2805
rect 40310 2796 40316 2848
rect 40368 2836 40374 2848
rect 41141 2839 41199 2845
rect 41141 2836 41153 2839
rect 40368 2808 41153 2836
rect 40368 2796 40374 2808
rect 41141 2805 41153 2808
rect 41187 2805 41199 2839
rect 41141 2799 41199 2805
rect 41690 2796 41696 2848
rect 41748 2836 41754 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41748 2808 42441 2836
rect 41748 2796 41754 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 42794 2796 42800 2848
rect 42852 2836 42858 2848
rect 43717 2839 43775 2845
rect 43717 2836 43729 2839
rect 42852 2808 43729 2836
rect 42852 2796 42858 2808
rect 43717 2805 43729 2808
rect 43763 2805 43775 2839
rect 43717 2799 43775 2805
rect 44174 2796 44180 2848
rect 44232 2836 44238 2848
rect 45005 2839 45063 2845
rect 45005 2836 45017 2839
rect 44232 2808 45017 2836
rect 44232 2796 44238 2808
rect 45005 2805 45017 2808
rect 45051 2805 45063 2839
rect 45005 2799 45063 2805
rect 45554 2796 45560 2848
rect 45612 2836 45618 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45612 2808 46305 2836
rect 45612 2796 45618 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 46658 2796 46664 2848
rect 46716 2836 46722 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46716 2808 47593 2836
rect 46716 2796 46722 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 48038 2796 48044 2848
rect 48096 2836 48102 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48096 2808 48881 2836
rect 48096 2796 48102 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49970 2796 49976 2848
rect 50028 2836 50034 2848
rect 50801 2839 50859 2845
rect 50801 2836 50813 2839
rect 50028 2808 50813 2836
rect 50028 2796 50034 2808
rect 50801 2805 50813 2808
rect 50847 2805 50859 2839
rect 50801 2799 50859 2805
rect 51902 2796 51908 2848
rect 51960 2836 51966 2848
rect 52733 2839 52791 2845
rect 52733 2836 52745 2839
rect 51960 2808 52745 2836
rect 51960 2796 51966 2808
rect 52733 2805 52745 2808
rect 52779 2805 52791 2839
rect 52733 2799 52791 2805
rect 53834 2796 53840 2848
rect 53892 2836 53898 2848
rect 54665 2839 54723 2845
rect 54665 2836 54677 2839
rect 53892 2808 54677 2836
rect 53892 2796 53898 2808
rect 54665 2805 54677 2808
rect 54711 2805 54723 2839
rect 54665 2799 54723 2805
rect 55398 2796 55404 2848
rect 55456 2836 55462 2848
rect 55953 2839 56011 2845
rect 55953 2836 55965 2839
rect 55456 2808 55965 2836
rect 55456 2796 55462 2808
rect 55953 2805 55965 2808
rect 55999 2805 56011 2839
rect 55953 2799 56011 2805
rect 56042 2796 56048 2848
rect 56100 2836 56106 2848
rect 57885 2839 57943 2845
rect 57885 2836 57897 2839
rect 56100 2808 57897 2836
rect 56100 2796 56106 2808
rect 57885 2805 57897 2808
rect 57931 2805 57943 2839
rect 57992 2836 58020 2876
rect 58529 2873 58541 2876
rect 58575 2873 58587 2907
rect 58529 2867 58587 2873
rect 59354 2864 59360 2916
rect 59412 2904 59418 2916
rect 63037 2907 63095 2913
rect 63037 2904 63049 2907
rect 59412 2876 63049 2904
rect 59412 2864 59418 2876
rect 63037 2873 63049 2876
rect 63083 2873 63095 2907
rect 63037 2867 63095 2873
rect 59173 2839 59231 2845
rect 59173 2836 59185 2839
rect 57992 2808 59185 2836
rect 57885 2799 57943 2805
rect 59173 2805 59185 2808
rect 59219 2805 59231 2839
rect 59173 2799 59231 2805
rect 59446 2796 59452 2848
rect 59504 2836 59510 2848
rect 59817 2839 59875 2845
rect 59817 2836 59829 2839
rect 59504 2808 59829 2836
rect 59504 2796 59510 2808
rect 59817 2805 59829 2808
rect 59863 2805 59875 2839
rect 60458 2836 60464 2848
rect 60419 2808 60464 2836
rect 59817 2799 59875 2805
rect 60458 2796 60464 2808
rect 60516 2796 60522 2848
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 4614 2632 4620 2644
rect 4571 2604 4620 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 6825 2635 6883 2641
rect 6825 2632 6837 2635
rect 6696 2604 6837 2632
rect 6696 2592 6702 2604
rect 6825 2601 6837 2604
rect 6871 2601 6883 2635
rect 6825 2595 6883 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 8352 2604 9505 2632
rect 8352 2592 8358 2604
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 9493 2595 9551 2601
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11296 2604 11621 2632
rect 11296 2592 11302 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 11977 2635 12035 2641
rect 11977 2601 11989 2635
rect 12023 2632 12035 2635
rect 12250 2632 12256 2644
rect 12023 2604 12256 2632
rect 12023 2601 12035 2604
rect 11977 2595 12035 2601
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 14829 2635 14887 2641
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 15010 2632 15016 2644
rect 14875 2604 15016 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 15010 2592 15016 2604
rect 15068 2592 15074 2644
rect 16761 2635 16819 2641
rect 16761 2601 16773 2635
rect 16807 2632 16819 2635
rect 17126 2632 17132 2644
rect 16807 2604 17132 2632
rect 16807 2601 16819 2604
rect 16761 2595 16819 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 19337 2635 19395 2641
rect 17236 2604 18368 2632
rect 2593 2567 2651 2573
rect 2593 2533 2605 2567
rect 2639 2564 2651 2567
rect 8110 2564 8116 2576
rect 2639 2536 8116 2564
rect 2639 2533 2651 2536
rect 2593 2527 2651 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 8205 2567 8263 2573
rect 8205 2533 8217 2567
rect 8251 2564 8263 2567
rect 10778 2564 10784 2576
rect 8251 2536 10784 2564
rect 8251 2533 8263 2536
rect 8205 2527 8263 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12434 2564 12440 2576
rect 12115 2536 12440 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 14458 2524 14464 2576
rect 14516 2564 14522 2576
rect 15841 2567 15899 2573
rect 15841 2564 15853 2567
rect 14516 2536 15853 2564
rect 14516 2524 14522 2536
rect 15841 2533 15853 2536
rect 15887 2533 15899 2567
rect 15841 2527 15899 2533
rect 2498 2456 2504 2508
rect 2556 2496 2562 2508
rect 10689 2499 10747 2505
rect 2556 2468 9720 2496
rect 2556 2456 2562 2468
rect 9692 2440 9720 2468
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 10735 2468 11897 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 11885 2465 11897 2468
rect 11931 2496 11943 2499
rect 12158 2496 12164 2508
rect 11931 2468 12164 2496
rect 11931 2465 11943 2468
rect 11885 2459 11943 2465
rect 12158 2456 12164 2468
rect 12216 2456 12222 2508
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 14550 2496 14556 2508
rect 14148 2468 14556 2496
rect 14148 2456 14154 2468
rect 14550 2456 14556 2468
rect 14608 2496 14614 2508
rect 14608 2468 16896 2496
rect 14608 2456 14614 2468
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1544 2400 1777 2428
rect 1544 2388 1550 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 1765 2391 1823 2397
rect 1780 2360 1808 2391
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4982 2428 4988 2440
rect 4387 2400 4988 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5626 2428 5632 2440
rect 5587 2400 5632 2428
rect 5626 2388 5632 2400
rect 5684 2428 5690 2440
rect 5902 2428 5908 2440
rect 5684 2400 5908 2428
rect 5684 2388 5690 2400
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 6178 2388 6184 2440
rect 6236 2428 6242 2440
rect 6638 2428 6644 2440
rect 6236 2400 6644 2428
rect 6236 2388 6242 2400
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 8018 2428 8024 2440
rect 7699 2400 8024 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 9674 2428 9680 2440
rect 9587 2400 9680 2428
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10560 2400 10977 2428
rect 10560 2388 10566 2400
rect 10965 2397 10977 2400
rect 11011 2428 11023 2431
rect 11514 2428 11520 2440
rect 11011 2400 11520 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 11974 2388 11980 2440
rect 12032 2428 12038 2440
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12032 2400 12449 2428
rect 12032 2388 12038 2400
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 12986 2428 12992 2440
rect 12947 2400 12992 2428
rect 12437 2391 12495 2397
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 13136 2400 13369 2428
rect 13136 2388 13142 2400
rect 13357 2397 13369 2400
rect 13403 2428 13415 2431
rect 16022 2428 16028 2440
rect 13403 2400 15424 2428
rect 15983 2400 16028 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 11054 2360 11060 2372
rect 1780 2332 11060 2360
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 12158 2320 12164 2372
rect 12216 2360 12222 2372
rect 13004 2360 13032 2388
rect 14550 2360 14556 2372
rect 12216 2332 13032 2360
rect 14511 2332 14556 2360
rect 12216 2320 12222 2332
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 15396 2360 15424 2400
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16868 2437 16896 2468
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17236 2360 17264 2604
rect 18230 2564 18236 2576
rect 18191 2536 18236 2564
rect 18230 2524 18236 2536
rect 18288 2524 18294 2576
rect 18340 2564 18368 2604
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 19978 2632 19984 2644
rect 19383 2604 19984 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 21726 2592 21732 2644
rect 21784 2632 21790 2644
rect 21821 2635 21879 2641
rect 21821 2632 21833 2635
rect 21784 2604 21833 2632
rect 21784 2592 21790 2604
rect 21821 2601 21833 2604
rect 21867 2601 21879 2635
rect 21821 2595 21879 2601
rect 21910 2592 21916 2644
rect 21968 2632 21974 2644
rect 26973 2635 27031 2641
rect 26973 2632 26985 2635
rect 21968 2604 26985 2632
rect 21968 2592 21974 2604
rect 26973 2601 26985 2604
rect 27019 2601 27031 2635
rect 26973 2595 27031 2601
rect 55214 2592 55220 2644
rect 55272 2632 55278 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 55272 2604 55321 2632
rect 55272 2592 55278 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 57422 2592 57428 2644
rect 57480 2632 57486 2644
rect 61105 2635 61163 2641
rect 61105 2632 61117 2635
rect 57480 2604 61117 2632
rect 57480 2592 57486 2604
rect 61105 2601 61117 2604
rect 61151 2601 61163 2635
rect 61105 2595 61163 2601
rect 20530 2564 20536 2576
rect 18340 2536 20536 2564
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 22094 2564 22100 2576
rect 20671 2536 22100 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 22094 2524 22100 2536
rect 22152 2524 22158 2576
rect 22557 2567 22615 2573
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 23198 2564 23204 2576
rect 22603 2536 23204 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 23198 2524 23204 2536
rect 23256 2524 23262 2576
rect 25777 2567 25835 2573
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 27338 2564 27344 2576
rect 25823 2536 27344 2564
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 27338 2524 27344 2536
rect 27396 2524 27402 2576
rect 28353 2567 28411 2573
rect 28353 2533 28365 2567
rect 28399 2564 28411 2567
rect 28994 2564 29000 2576
rect 28399 2536 29000 2564
rect 28399 2533 28411 2536
rect 28353 2527 28411 2533
rect 28994 2524 29000 2536
rect 29052 2524 29058 2576
rect 30285 2567 30343 2573
rect 30285 2533 30297 2567
rect 30331 2564 30343 2567
rect 30926 2564 30932 2576
rect 30331 2536 30932 2564
rect 30331 2533 30343 2536
rect 30285 2527 30343 2533
rect 30926 2524 30932 2536
rect 30984 2524 30990 2576
rect 40586 2524 40592 2576
rect 40644 2564 40650 2576
rect 42429 2567 42487 2573
rect 42429 2564 42441 2567
rect 40644 2536 42441 2564
rect 40644 2524 40650 2536
rect 42429 2533 42441 2536
rect 42475 2533 42487 2567
rect 42429 2527 42487 2533
rect 44450 2524 44456 2576
rect 44508 2564 44514 2576
rect 46293 2567 46351 2573
rect 46293 2564 46305 2567
rect 44508 2536 46305 2564
rect 44508 2524 44514 2536
rect 46293 2533 46305 2536
rect 46339 2533 46351 2567
rect 46293 2527 46351 2533
rect 48314 2524 48320 2576
rect 48372 2564 48378 2576
rect 50157 2567 50215 2573
rect 50157 2564 50169 2567
rect 48372 2536 50169 2564
rect 48372 2524 48378 2536
rect 50157 2533 50169 2536
rect 50203 2533 50215 2567
rect 50157 2527 50215 2533
rect 52178 2524 52184 2576
rect 52236 2564 52242 2576
rect 54021 2567 54079 2573
rect 54021 2564 54033 2567
rect 52236 2536 54033 2564
rect 52236 2524 52242 2536
rect 54021 2533 54033 2536
rect 54067 2533 54079 2567
rect 54021 2527 54079 2533
rect 55858 2524 55864 2576
rect 55916 2564 55922 2576
rect 57885 2567 57943 2573
rect 57885 2564 57897 2567
rect 55916 2536 57897 2564
rect 55916 2524 55922 2536
rect 57885 2533 57897 2536
rect 57931 2533 57943 2567
rect 57885 2527 57943 2533
rect 58066 2524 58072 2576
rect 58124 2564 58130 2576
rect 58529 2567 58587 2573
rect 58529 2564 58541 2567
rect 58124 2536 58541 2564
rect 58124 2524 58130 2536
rect 58529 2533 58541 2536
rect 58575 2533 58587 2567
rect 58529 2527 58587 2533
rect 60461 2567 60519 2573
rect 60461 2533 60473 2567
rect 60507 2533 60519 2567
rect 60461 2527 60519 2533
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 21910 2496 21916 2508
rect 17920 2468 21916 2496
rect 17920 2456 17926 2468
rect 21910 2456 21916 2468
rect 21968 2456 21974 2508
rect 22002 2456 22008 2508
rect 22060 2496 22066 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 22060 2468 24409 2496
rect 22060 2456 22066 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 25133 2499 25191 2505
rect 25133 2465 25145 2499
rect 25179 2496 25191 2499
rect 26510 2496 26516 2508
rect 25179 2468 26516 2496
rect 25179 2465 25191 2468
rect 25133 2459 25191 2465
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 36998 2456 37004 2508
rect 37056 2496 37062 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 37056 2468 37933 2496
rect 37056 2456 37062 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 38102 2456 38108 2508
rect 38160 2496 38166 2508
rect 39853 2499 39911 2505
rect 39853 2496 39865 2499
rect 38160 2468 39865 2496
rect 38160 2456 38166 2468
rect 39853 2465 39865 2468
rect 39899 2465 39911 2499
rect 39853 2459 39911 2465
rect 41414 2456 41420 2508
rect 41472 2496 41478 2508
rect 43073 2499 43131 2505
rect 43073 2496 43085 2499
rect 41472 2468 43085 2496
rect 41472 2456 41478 2468
rect 43073 2465 43085 2468
rect 43119 2465 43131 2499
rect 43073 2459 43131 2465
rect 43346 2456 43352 2508
rect 43404 2496 43410 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 43404 2468 45017 2496
rect 43404 2456 43410 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45005 2459 45063 2465
rect 46382 2456 46388 2508
rect 46440 2496 46446 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 46440 2468 48237 2496
rect 46440 2456 46446 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 49142 2456 49148 2508
rect 49200 2496 49206 2508
rect 50801 2499 50859 2505
rect 50801 2496 50813 2499
rect 49200 2468 50813 2496
rect 49200 2456 49206 2468
rect 50801 2465 50813 2468
rect 50847 2465 50859 2499
rect 50801 2459 50859 2465
rect 51074 2456 51080 2508
rect 51132 2496 51138 2508
rect 52733 2499 52791 2505
rect 52733 2496 52745 2499
rect 51132 2468 52745 2496
rect 51132 2456 51138 2468
rect 52733 2465 52745 2468
rect 52779 2465 52791 2499
rect 52733 2459 52791 2465
rect 54938 2456 54944 2508
rect 54996 2496 55002 2508
rect 56597 2499 56655 2505
rect 56597 2496 56609 2499
rect 54996 2468 56609 2496
rect 54996 2456 55002 2468
rect 56597 2465 56609 2468
rect 56643 2465 56655 2499
rect 60476 2496 60504 2527
rect 63678 2496 63684 2508
rect 60476 2468 60596 2496
rect 63639 2468 63684 2496
rect 56597 2459 56655 2465
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2428 17739 2431
rect 17880 2428 17908 2456
rect 17727 2400 17908 2428
rect 18417 2431 18475 2437
rect 17727 2397 17739 2400
rect 17681 2391 17739 2397
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2428 20039 2431
rect 20990 2428 20996 2440
rect 20027 2400 20996 2428
rect 20027 2397 20039 2400
rect 19981 2391 20039 2397
rect 18432 2360 18460 2391
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22370 2428 22376 2440
rect 21315 2400 22376 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22370 2388 22376 2400
rect 22428 2388 22434 2440
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 25406 2428 25412 2440
rect 23891 2400 25412 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 22002 2360 22008 2372
rect 15396 2332 17264 2360
rect 17420 2332 22008 2360
rect 1946 2292 1952 2304
rect 1907 2264 1952 2292
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 3234 2292 3240 2304
rect 3195 2264 3240 2292
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 3878 2292 3884 2304
rect 3839 2264 3884 2292
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 7469 2295 7527 2301
rect 7469 2261 7481 2295
rect 7515 2292 7527 2295
rect 10318 2292 10324 2304
rect 7515 2264 10324 2292
rect 7515 2261 7527 2264
rect 7469 2255 7527 2261
rect 10318 2252 10324 2264
rect 10376 2252 10382 2304
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 17420 2292 17448 2332
rect 22002 2320 22008 2332
rect 22060 2320 22066 2372
rect 23216 2360 23244 2391
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2397 26479 2431
rect 26421 2391 26479 2397
rect 27709 2431 27767 2437
rect 27709 2397 27721 2431
rect 27755 2428 27767 2431
rect 28442 2428 28448 2440
rect 27755 2400 28448 2428
rect 27755 2397 27767 2400
rect 27709 2391 27767 2397
rect 24578 2360 24584 2372
rect 23216 2332 24584 2360
rect 24578 2320 24584 2332
rect 24636 2320 24642 2372
rect 26436 2360 26464 2391
rect 28442 2388 28448 2400
rect 28500 2388 28506 2440
rect 28997 2431 29055 2437
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 29546 2428 29552 2440
rect 29043 2400 29552 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 30929 2431 30987 2437
rect 30929 2397 30941 2431
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 31573 2431 31631 2437
rect 31573 2397 31585 2431
rect 31619 2428 31631 2431
rect 32582 2428 32588 2440
rect 31619 2400 32588 2428
rect 31619 2397 31631 2400
rect 31573 2391 31631 2397
rect 27890 2360 27896 2372
rect 26436 2332 27896 2360
rect 27890 2320 27896 2332
rect 27948 2320 27954 2372
rect 30944 2360 30972 2391
rect 32582 2388 32588 2400
rect 32640 2388 32646 2440
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 33410 2428 33416 2440
rect 32907 2400 33416 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 33410 2388 33416 2400
rect 33468 2388 33474 2440
rect 33505 2431 33563 2437
rect 33505 2397 33517 2431
rect 33551 2428 33563 2431
rect 33962 2428 33968 2440
rect 33551 2400 33968 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 33962 2388 33968 2400
rect 34020 2388 34026 2440
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34790 2428 34796 2440
rect 34195 2400 34796 2428
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 34790 2388 34796 2400
rect 34848 2388 34854 2440
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2428 34943 2431
rect 35066 2428 35072 2440
rect 34931 2400 35072 2428
rect 34931 2397 34943 2400
rect 34885 2391 34943 2397
rect 35066 2388 35072 2400
rect 35124 2388 35130 2440
rect 35529 2431 35587 2437
rect 35529 2397 35541 2431
rect 35575 2428 35587 2431
rect 35618 2428 35624 2440
rect 35575 2400 35624 2428
rect 35575 2397 35587 2400
rect 35529 2391 35587 2397
rect 35618 2388 35624 2400
rect 35676 2388 35682 2440
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35952 2400 36001 2428
rect 35952 2388 35958 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36446 2388 36452 2440
rect 36504 2428 36510 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36504 2400 37289 2428
rect 36504 2388 36510 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37550 2388 37556 2440
rect 37608 2428 37614 2440
rect 38565 2431 38623 2437
rect 38565 2428 38577 2431
rect 37608 2400 38577 2428
rect 37608 2388 37614 2400
rect 38565 2397 38577 2400
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 40497 2431 40555 2437
rect 40497 2428 40509 2431
rect 38712 2400 40509 2428
rect 38712 2388 38718 2400
rect 40497 2397 40509 2400
rect 40543 2397 40555 2431
rect 40497 2391 40555 2397
rect 41141 2431 41199 2437
rect 41141 2397 41153 2431
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 31754 2360 31760 2372
rect 30944 2332 31760 2360
rect 31754 2320 31760 2332
rect 31812 2320 31818 2372
rect 39482 2320 39488 2372
rect 39540 2360 39546 2372
rect 41156 2360 41184 2391
rect 41966 2388 41972 2440
rect 42024 2428 42030 2440
rect 43717 2431 43775 2437
rect 43717 2428 43729 2431
rect 42024 2400 43729 2428
rect 42024 2388 42030 2400
rect 43717 2397 43729 2400
rect 43763 2397 43775 2431
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 43717 2391 43775 2397
rect 45526 2400 45661 2428
rect 39540 2332 41184 2360
rect 39540 2320 39546 2332
rect 43898 2320 43904 2372
rect 43956 2360 43962 2372
rect 45526 2360 45554 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 45830 2388 45836 2440
rect 45888 2428 45894 2440
rect 47581 2431 47639 2437
rect 47581 2428 47593 2431
rect 45888 2400 47593 2428
rect 45888 2388 45894 2400
rect 47581 2397 47593 2400
rect 47627 2397 47639 2431
rect 47581 2391 47639 2397
rect 48869 2431 48927 2437
rect 48869 2397 48881 2431
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 43956 2332 45554 2360
rect 43956 2320 43962 2332
rect 47210 2320 47216 2372
rect 47268 2360 47274 2372
rect 48884 2360 48912 2391
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 51445 2431 51503 2437
rect 51445 2428 51457 2431
rect 49752 2400 51457 2428
rect 49752 2388 49758 2400
rect 51445 2397 51457 2400
rect 51491 2397 51503 2431
rect 51445 2391 51503 2397
rect 51626 2388 51632 2440
rect 51684 2428 51690 2440
rect 53377 2431 53435 2437
rect 53377 2428 53389 2431
rect 51684 2400 53389 2428
rect 51684 2388 51690 2400
rect 53377 2397 53389 2400
rect 53423 2397 53435 2431
rect 53377 2391 53435 2397
rect 55953 2431 56011 2437
rect 55953 2397 55965 2431
rect 55999 2397 56011 2431
rect 55953 2391 56011 2397
rect 47268 2332 48912 2360
rect 47268 2320 47274 2332
rect 54110 2320 54116 2372
rect 54168 2360 54174 2372
rect 55968 2360 55996 2391
rect 56410 2388 56416 2440
rect 56468 2428 56474 2440
rect 59173 2431 59231 2437
rect 59173 2428 59185 2431
rect 56468 2400 59185 2428
rect 56468 2388 56474 2400
rect 59173 2397 59185 2400
rect 59219 2397 59231 2431
rect 59173 2391 59231 2397
rect 54168 2332 55996 2360
rect 54168 2320 54174 2332
rect 13780 2264 17448 2292
rect 17497 2295 17555 2301
rect 13780 2252 13786 2264
rect 17497 2261 17509 2295
rect 17543 2292 17555 2295
rect 17586 2292 17592 2304
rect 17543 2264 17592 2292
rect 17543 2261 17555 2264
rect 17497 2255 17555 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 56870 2252 56876 2304
rect 56928 2292 56934 2304
rect 60568 2292 60596 2468
rect 63678 2456 63684 2468
rect 63736 2456 63742 2508
rect 61746 2428 61752 2440
rect 61707 2400 61752 2428
rect 61746 2388 61752 2400
rect 61804 2388 61810 2440
rect 63034 2428 63040 2440
rect 62995 2400 63040 2428
rect 63034 2388 63040 2400
rect 63092 2388 63098 2440
rect 66990 2428 66996 2440
rect 66951 2400 66996 2428
rect 66990 2388 66996 2400
rect 67048 2388 67054 2440
rect 67542 2388 67548 2440
rect 67600 2428 67606 2440
rect 67637 2431 67695 2437
rect 67637 2428 67649 2431
rect 67600 2400 67649 2428
rect 67600 2388 67606 2400
rect 67637 2397 67649 2400
rect 67683 2397 67695 2431
rect 67637 2391 67695 2397
rect 56928 2264 60596 2292
rect 56928 2252 56934 2264
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
rect 6638 2048 6644 2100
rect 6696 2088 6702 2100
rect 11238 2088 11244 2100
rect 6696 2060 11244 2088
rect 6696 2048 6702 2060
rect 11238 2048 11244 2060
rect 11296 2048 11302 2100
rect 14550 2088 14556 2100
rect 12406 2060 14556 2088
rect 3878 1980 3884 2032
rect 3936 2020 3942 2032
rect 11974 2020 11980 2032
rect 3936 1992 11980 2020
rect 3936 1980 3942 1992
rect 11974 1980 11980 1992
rect 12032 2020 12038 2032
rect 12406 2020 12434 2060
rect 14550 2048 14556 2060
rect 14608 2048 14614 2100
rect 18782 2048 18788 2100
rect 18840 2088 18846 2100
rect 19794 2088 19800 2100
rect 18840 2060 19800 2088
rect 18840 2048 18846 2060
rect 19794 2048 19800 2060
rect 19852 2048 19858 2100
rect 58066 2048 58072 2100
rect 58124 2088 58130 2100
rect 61746 2088 61752 2100
rect 58124 2060 61752 2088
rect 58124 2048 58130 2060
rect 61746 2048 61752 2060
rect 61804 2048 61810 2100
rect 12032 1992 12434 2020
rect 12032 1980 12038 1992
rect 17586 1980 17592 2032
rect 17644 2020 17650 2032
rect 24670 2020 24676 2032
rect 17644 1992 24676 2020
rect 17644 1980 17650 1992
rect 24670 1980 24676 1992
rect 24728 1980 24734 2032
rect 59078 1980 59084 2032
rect 59136 2020 59142 2032
rect 63678 2020 63684 2032
rect 59136 1992 63684 2020
rect 59136 1980 59142 1992
rect 63678 1980 63684 1992
rect 63736 1980 63742 2032
rect 5074 1912 5080 1964
rect 5132 1952 5138 1964
rect 14642 1952 14648 1964
rect 5132 1924 14648 1952
rect 5132 1912 5138 1924
rect 14642 1912 14648 1924
rect 14700 1912 14706 1964
rect 58526 1912 58532 1964
rect 58584 1952 58590 1964
rect 63034 1952 63040 1964
rect 58584 1924 63040 1952
rect 58584 1912 58590 1924
rect 63034 1912 63040 1924
rect 63092 1912 63098 1964
rect 5626 1844 5632 1896
rect 5684 1884 5690 1896
rect 12710 1884 12716 1896
rect 5684 1856 12716 1884
rect 5684 1844 5690 1856
rect 12710 1844 12716 1856
rect 12768 1844 12774 1896
rect 3234 1776 3240 1828
rect 3292 1816 3298 1828
rect 12618 1816 12624 1828
rect 3292 1788 12624 1816
rect 3292 1776 3298 1788
rect 12618 1776 12624 1788
rect 12676 1776 12682 1828
rect 9674 1708 9680 1760
rect 9732 1748 9738 1760
rect 9732 1720 13032 1748
rect 9732 1708 9738 1720
rect 8110 1640 8116 1692
rect 8168 1680 8174 1692
rect 10042 1680 10048 1692
rect 8168 1652 10048 1680
rect 8168 1640 8174 1652
rect 10042 1640 10048 1652
rect 10100 1640 10106 1692
rect 9766 1572 9772 1624
rect 9824 1612 9830 1624
rect 10686 1612 10692 1624
rect 9824 1584 10692 1612
rect 9824 1572 9830 1584
rect 10686 1572 10692 1584
rect 10744 1572 10750 1624
rect 10318 1436 10324 1488
rect 10376 1476 10382 1488
rect 10376 1448 11008 1476
rect 10376 1436 10382 1448
rect 10134 1368 10140 1420
rect 10192 1408 10198 1420
rect 10870 1408 10876 1420
rect 10192 1380 10876 1408
rect 10192 1368 10198 1380
rect 10870 1368 10876 1380
rect 10928 1368 10934 1420
rect 10980 1408 11008 1448
rect 12434 1408 12440 1420
rect 10980 1380 12440 1408
rect 12434 1368 12440 1380
rect 12492 1368 12498 1420
rect 12710 1368 12716 1420
rect 12768 1408 12774 1420
rect 12768 1380 12940 1408
rect 12768 1368 12774 1380
rect 12912 1352 12940 1380
rect 13004 1352 13032 1720
rect 14274 1436 14280 1488
rect 14332 1476 14338 1488
rect 15010 1476 15016 1488
rect 14332 1448 15016 1476
rect 14332 1436 14338 1448
rect 15010 1436 15016 1448
rect 15068 1436 15074 1488
rect 13722 1408 13728 1420
rect 13096 1380 13728 1408
rect 12894 1300 12900 1352
rect 12952 1300 12958 1352
rect 12986 1300 12992 1352
rect 13044 1300 13050 1352
rect 12710 1232 12716 1284
rect 12768 1272 12774 1284
rect 13096 1272 13124 1380
rect 13722 1368 13728 1380
rect 13780 1368 13786 1420
rect 14182 1368 14188 1420
rect 14240 1408 14246 1420
rect 14826 1408 14832 1420
rect 14240 1380 14832 1408
rect 14240 1368 14246 1380
rect 14826 1368 14832 1380
rect 14884 1368 14890 1420
rect 19518 1300 19524 1352
rect 19576 1340 19582 1352
rect 20346 1340 20352 1352
rect 19576 1312 20352 1340
rect 19576 1300 19582 1312
rect 20346 1300 20352 1312
rect 20404 1300 20410 1352
rect 12768 1244 13124 1272
rect 12768 1232 12774 1244
rect 12802 1164 12808 1216
rect 12860 1204 12866 1216
rect 15654 1204 15660 1216
rect 12860 1176 15660 1204
rect 12860 1164 12866 1176
rect 15654 1164 15660 1176
rect 15712 1164 15718 1216
rect 56778 1164 56784 1216
rect 56836 1204 56842 1216
rect 57054 1204 57060 1216
rect 56836 1176 57060 1204
rect 56836 1164 56842 1176
rect 57054 1164 57060 1176
rect 57112 1164 57118 1216
rect 12342 1096 12348 1148
rect 12400 1096 12406 1148
rect 19334 1096 19340 1148
rect 19392 1136 19398 1148
rect 19702 1136 19708 1148
rect 19392 1108 19708 1136
rect 19392 1096 19398 1108
rect 19702 1096 19708 1108
rect 19760 1096 19766 1148
rect 12250 892 12256 944
rect 12308 932 12314 944
rect 12360 932 12388 1096
rect 57054 1028 57060 1080
rect 57112 1068 57118 1080
rect 59446 1068 59452 1080
rect 57112 1040 59452 1068
rect 57112 1028 57118 1040
rect 59446 1028 59452 1040
rect 59504 1028 59510 1080
rect 12308 904 12388 932
rect 12308 892 12314 904
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 5172 57400 5224 57452
rect 15200 57443 15252 57452
rect 15200 57409 15209 57443
rect 15209 57409 15243 57443
rect 15243 57409 15252 57443
rect 15200 57400 15252 57409
rect 25044 57400 25096 57452
rect 34980 57400 35032 57452
rect 44916 57400 44968 57452
rect 54852 57400 54904 57452
rect 64788 57400 64840 57452
rect 66996 57443 67048 57452
rect 66996 57409 67005 57443
rect 67005 57409 67039 57443
rect 67039 57409 67048 57443
rect 66996 57400 67048 57409
rect 67548 57400 67600 57452
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 68100 56831 68152 56840
rect 68100 56797 68109 56831
rect 68109 56797 68143 56831
rect 68143 56797 68152 56831
rect 68100 56788 68152 56797
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 67640 55131 67692 55140
rect 67640 55097 67649 55131
rect 67649 55097 67683 55131
rect 67683 55097 67692 55131
rect 67640 55088 67692 55097
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 67548 53932 67600 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 68100 52479 68152 52488
rect 68100 52445 68109 52479
rect 68109 52445 68143 52479
rect 68143 52445 68152 52479
rect 68100 52436 68152 52445
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 68100 51391 68152 51400
rect 68100 51357 68109 51391
rect 68109 51357 68143 51391
rect 68143 51357 68152 51391
rect 68100 51348 68152 51357
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 67640 49759 67692 49768
rect 67640 49725 67649 49759
rect 67649 49725 67683 49759
rect 67683 49725 67692 49759
rect 67640 49716 67692 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 67640 48535 67692 48544
rect 67640 48501 67649 48535
rect 67649 48501 67683 48535
rect 67683 48501 67692 48535
rect 67640 48492 67692 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 68100 47039 68152 47048
rect 68100 47005 68109 47039
rect 68109 47005 68143 47039
rect 68143 47005 68152 47039
rect 68100 46996 68152 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 68100 45951 68152 45960
rect 68100 45917 68109 45951
rect 68109 45917 68143 45951
rect 68143 45917 68152 45951
rect 68100 45908 68152 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 67640 44251 67692 44260
rect 67640 44217 67649 44251
rect 67649 44217 67683 44251
rect 67683 44217 67692 44251
rect 67640 44208 67692 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 67640 43095 67692 43104
rect 67640 43061 67649 43095
rect 67649 43061 67683 43095
rect 67683 43061 67692 43095
rect 67640 43052 67692 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 68100 41599 68152 41608
rect 68100 41565 68109 41599
rect 68109 41565 68143 41599
rect 68143 41565 68152 41599
rect 68100 41556 68152 41565
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 68100 40511 68152 40520
rect 68100 40477 68109 40511
rect 68109 40477 68143 40511
rect 68143 40477 68152 40511
rect 68100 40468 68152 40477
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 67640 38811 67692 38820
rect 67640 38777 67649 38811
rect 67649 38777 67683 38811
rect 67683 38777 67692 38811
rect 67640 38768 67692 38777
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 67640 37655 67692 37664
rect 67640 37621 67649 37655
rect 67649 37621 67683 37655
rect 67683 37621 67692 37655
rect 67640 37612 67692 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 68100 36159 68152 36168
rect 68100 36125 68109 36159
rect 68109 36125 68143 36159
rect 68143 36125 68152 36159
rect 68100 36116 68152 36125
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 68100 35071 68152 35080
rect 68100 35037 68109 35071
rect 68109 35037 68143 35071
rect 68143 35037 68152 35071
rect 68100 35028 68152 35037
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 67640 33371 67692 33380
rect 67640 33337 67649 33371
rect 67649 33337 67683 33371
rect 67683 33337 67692 33371
rect 67640 33328 67692 33337
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 67640 32215 67692 32224
rect 67640 32181 67649 32215
rect 67649 32181 67683 32215
rect 67683 32181 67692 32215
rect 67640 32172 67692 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 15108 31696 15160 31748
rect 20536 31696 20588 31748
rect 17408 31628 17460 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 7840 31356 7892 31408
rect 8392 31288 8444 31340
rect 12072 31331 12124 31340
rect 12072 31297 12081 31331
rect 12081 31297 12115 31331
rect 12115 31297 12124 31331
rect 12072 31288 12124 31297
rect 12624 31288 12676 31340
rect 12900 31331 12952 31340
rect 12900 31297 12909 31331
rect 12909 31297 12943 31331
rect 12943 31297 12952 31331
rect 12900 31288 12952 31297
rect 15292 31356 15344 31408
rect 13176 31331 13228 31340
rect 13176 31297 13185 31331
rect 13185 31297 13219 31331
rect 13219 31297 13228 31331
rect 13176 31288 13228 31297
rect 15200 31331 15252 31340
rect 15200 31297 15209 31331
rect 15209 31297 15243 31331
rect 15243 31297 15252 31331
rect 15200 31288 15252 31297
rect 16672 31288 16724 31340
rect 17776 31356 17828 31408
rect 22744 31356 22796 31408
rect 23020 31356 23072 31408
rect 17224 31331 17276 31340
rect 17224 31297 17233 31331
rect 17233 31297 17267 31331
rect 17267 31297 17276 31331
rect 17224 31288 17276 31297
rect 15476 31152 15528 31204
rect 16580 31152 16632 31204
rect 17408 31331 17460 31340
rect 17408 31297 17417 31331
rect 17417 31297 17451 31331
rect 17451 31297 17460 31331
rect 20536 31331 20588 31340
rect 17408 31288 17460 31297
rect 20536 31297 20545 31331
rect 20545 31297 20579 31331
rect 20579 31297 20588 31331
rect 20536 31288 20588 31297
rect 20720 31331 20772 31340
rect 20720 31297 20729 31331
rect 20729 31297 20763 31331
rect 20763 31297 20772 31331
rect 20720 31288 20772 31297
rect 20904 31331 20956 31340
rect 20904 31297 20913 31331
rect 20913 31297 20947 31331
rect 20947 31297 20956 31331
rect 23296 31331 23348 31340
rect 20904 31288 20956 31297
rect 23296 31297 23305 31331
rect 23305 31297 23339 31331
rect 23339 31297 23348 31331
rect 23296 31288 23348 31297
rect 24032 31288 24084 31340
rect 22100 31220 22152 31272
rect 23756 31220 23808 31272
rect 24492 31331 24544 31340
rect 24492 31297 24501 31331
rect 24501 31297 24535 31331
rect 24535 31297 24544 31331
rect 24492 31288 24544 31297
rect 17776 31152 17828 31204
rect 9404 31084 9456 31136
rect 13544 31127 13596 31136
rect 13544 31093 13553 31127
rect 13553 31093 13587 31127
rect 13587 31093 13596 31127
rect 13544 31084 13596 31093
rect 15384 31127 15436 31136
rect 15384 31093 15393 31127
rect 15393 31093 15427 31127
rect 15427 31093 15436 31127
rect 15384 31084 15436 31093
rect 18052 31084 18104 31136
rect 20260 31127 20312 31136
rect 20260 31093 20269 31127
rect 20269 31093 20303 31127
rect 20303 31093 20312 31127
rect 20260 31084 20312 31093
rect 26148 31084 26200 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 9312 30880 9364 30932
rect 15108 30880 15160 30932
rect 17224 30880 17276 30932
rect 20720 30880 20772 30932
rect 8392 30719 8444 30728
rect 8392 30685 8401 30719
rect 8401 30685 8435 30719
rect 8435 30685 8444 30719
rect 8392 30676 8444 30685
rect 8208 30651 8260 30660
rect 8208 30617 8217 30651
rect 8217 30617 8251 30651
rect 8251 30617 8260 30651
rect 8208 30608 8260 30617
rect 9312 30676 9364 30728
rect 9680 30744 9732 30796
rect 13268 30812 13320 30864
rect 9772 30719 9824 30728
rect 9772 30685 9781 30719
rect 9781 30685 9815 30719
rect 9815 30685 9824 30719
rect 11888 30744 11940 30796
rect 17408 30812 17460 30864
rect 9772 30676 9824 30685
rect 9680 30608 9732 30660
rect 9128 30583 9180 30592
rect 9128 30549 9137 30583
rect 9137 30549 9171 30583
rect 9171 30549 9180 30583
rect 9128 30540 9180 30549
rect 11336 30583 11388 30592
rect 11336 30549 11345 30583
rect 11345 30549 11379 30583
rect 11379 30549 11388 30583
rect 11336 30540 11388 30549
rect 11980 30719 12032 30728
rect 11980 30685 11989 30719
rect 11989 30685 12023 30719
rect 12023 30685 12032 30719
rect 11980 30676 12032 30685
rect 15108 30676 15160 30728
rect 15384 30719 15436 30728
rect 15384 30685 15393 30719
rect 15393 30685 15427 30719
rect 15427 30685 15436 30719
rect 15384 30676 15436 30685
rect 16212 30719 16264 30728
rect 16212 30685 16221 30719
rect 16221 30685 16255 30719
rect 16255 30685 16264 30719
rect 16212 30676 16264 30685
rect 16580 30744 16632 30796
rect 18420 30744 18472 30796
rect 16396 30719 16448 30728
rect 16396 30685 16405 30719
rect 16405 30685 16439 30719
rect 16439 30685 16448 30719
rect 16396 30676 16448 30685
rect 16672 30608 16724 30660
rect 14924 30583 14976 30592
rect 14924 30549 14933 30583
rect 14933 30549 14967 30583
rect 14967 30549 14976 30583
rect 14924 30540 14976 30549
rect 15292 30540 15344 30592
rect 17224 30608 17276 30660
rect 20720 30676 20772 30728
rect 68100 30719 68152 30728
rect 68100 30685 68109 30719
rect 68109 30685 68143 30719
rect 68143 30685 68152 30719
rect 68100 30676 68152 30685
rect 20628 30651 20680 30660
rect 20628 30617 20637 30651
rect 20637 30617 20671 30651
rect 20671 30617 20680 30651
rect 20628 30608 20680 30617
rect 18328 30540 18380 30592
rect 24400 30583 24452 30592
rect 24400 30549 24409 30583
rect 24409 30549 24443 30583
rect 24443 30549 24452 30583
rect 24400 30540 24452 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 7840 30336 7892 30388
rect 11888 30379 11940 30388
rect 11888 30345 11897 30379
rect 11897 30345 11931 30379
rect 11931 30345 11940 30379
rect 11888 30336 11940 30345
rect 16212 30336 16264 30388
rect 3792 30200 3844 30252
rect 9128 30268 9180 30320
rect 9680 30268 9732 30320
rect 10416 30268 10468 30320
rect 13544 30268 13596 30320
rect 6828 30175 6880 30184
rect 6828 30141 6837 30175
rect 6837 30141 6871 30175
rect 6871 30141 6880 30175
rect 6828 30132 6880 30141
rect 9404 30243 9456 30252
rect 9404 30209 9413 30243
rect 9413 30209 9447 30243
rect 9447 30209 9456 30243
rect 9404 30200 9456 30209
rect 12072 30200 12124 30252
rect 12440 30200 12492 30252
rect 17316 30268 17368 30320
rect 18052 30268 18104 30320
rect 20260 30268 20312 30320
rect 23296 30268 23348 30320
rect 24952 30268 25004 30320
rect 15292 30243 15344 30252
rect 15292 30209 15301 30243
rect 15301 30209 15335 30243
rect 15335 30209 15344 30243
rect 15292 30200 15344 30209
rect 18880 30243 18932 30252
rect 18880 30209 18889 30243
rect 18889 30209 18923 30243
rect 18923 30209 18932 30243
rect 18880 30200 18932 30209
rect 21916 30200 21968 30252
rect 24492 30200 24544 30252
rect 26148 30243 26200 30252
rect 26148 30209 26166 30243
rect 26166 30209 26200 30243
rect 26148 30200 26200 30209
rect 27620 30200 27672 30252
rect 28264 30200 28316 30252
rect 12900 30132 12952 30184
rect 14004 30175 14056 30184
rect 14004 30141 14013 30175
rect 14013 30141 14047 30175
rect 14047 30141 14056 30175
rect 14004 30132 14056 30141
rect 21824 30175 21876 30184
rect 21824 30141 21833 30175
rect 21833 30141 21867 30175
rect 21867 30141 21876 30175
rect 21824 30132 21876 30141
rect 8208 30039 8260 30048
rect 8208 30005 8217 30039
rect 8217 30005 8251 30039
rect 8251 30005 8260 30039
rect 8208 29996 8260 30005
rect 12624 30039 12676 30048
rect 12624 30005 12633 30039
rect 12633 30005 12667 30039
rect 12667 30005 12676 30039
rect 12624 29996 12676 30005
rect 17776 30064 17828 30116
rect 23020 30064 23072 30116
rect 16396 29996 16448 30048
rect 17132 29996 17184 30048
rect 20720 30039 20772 30048
rect 20720 30005 20729 30039
rect 20729 30005 20763 30039
rect 20763 30005 20772 30039
rect 20720 29996 20772 30005
rect 22468 29996 22520 30048
rect 23112 29996 23164 30048
rect 23940 29996 23992 30048
rect 29276 29996 29328 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 10140 29792 10192 29844
rect 10416 29835 10468 29844
rect 10416 29801 10425 29835
rect 10425 29801 10459 29835
rect 10459 29801 10468 29835
rect 10416 29792 10468 29801
rect 11980 29792 12032 29844
rect 16764 29792 16816 29844
rect 17316 29835 17368 29844
rect 17316 29801 17325 29835
rect 17325 29801 17359 29835
rect 17359 29801 17368 29835
rect 17316 29792 17368 29801
rect 18328 29792 18380 29844
rect 21548 29792 21600 29844
rect 21916 29792 21968 29844
rect 3792 29699 3844 29708
rect 3792 29665 3801 29699
rect 3801 29665 3835 29699
rect 3835 29665 3844 29699
rect 3792 29656 3844 29665
rect 10508 29588 10560 29640
rect 14004 29656 14056 29708
rect 3332 29520 3384 29572
rect 11336 29520 11388 29572
rect 5172 29495 5224 29504
rect 5172 29461 5181 29495
rect 5181 29461 5215 29495
rect 5215 29461 5224 29495
rect 5172 29452 5224 29461
rect 11060 29452 11112 29504
rect 12716 29631 12768 29640
rect 12716 29597 12725 29631
rect 12725 29597 12759 29631
rect 12759 29597 12768 29631
rect 12716 29588 12768 29597
rect 12900 29631 12952 29640
rect 12900 29597 12909 29631
rect 12909 29597 12943 29631
rect 12943 29597 12952 29631
rect 12900 29588 12952 29597
rect 18052 29588 18104 29640
rect 18880 29588 18932 29640
rect 20904 29588 20956 29640
rect 23756 29724 23808 29776
rect 13268 29520 13320 29572
rect 15568 29452 15620 29504
rect 16212 29520 16264 29572
rect 18420 29563 18472 29572
rect 18420 29529 18438 29563
rect 18438 29529 18472 29563
rect 21548 29631 21600 29640
rect 21548 29597 21557 29631
rect 21557 29597 21591 29631
rect 21591 29597 21600 29631
rect 22468 29631 22520 29640
rect 21548 29588 21600 29597
rect 22468 29597 22477 29631
rect 22477 29597 22511 29631
rect 22511 29597 22520 29631
rect 22468 29588 22520 29597
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 23296 29588 23348 29640
rect 18420 29520 18472 29529
rect 22100 29520 22152 29572
rect 24032 29588 24084 29640
rect 24952 29631 25004 29640
rect 24952 29597 24961 29631
rect 24961 29597 24995 29631
rect 24995 29597 25004 29631
rect 24952 29588 25004 29597
rect 27620 29588 27672 29640
rect 68100 29631 68152 29640
rect 68100 29597 68109 29631
rect 68109 29597 68143 29631
rect 68143 29597 68152 29631
rect 68100 29588 68152 29597
rect 16672 29452 16724 29504
rect 17592 29452 17644 29504
rect 23296 29452 23348 29504
rect 23940 29520 23992 29572
rect 25228 29563 25280 29572
rect 25228 29529 25262 29563
rect 25262 29529 25280 29563
rect 25228 29520 25280 29529
rect 25596 29520 25648 29572
rect 25136 29452 25188 29504
rect 25872 29452 25924 29504
rect 27804 29520 27856 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 6736 29248 6788 29300
rect 12164 29291 12216 29300
rect 6828 29180 6880 29232
rect 11796 29223 11848 29232
rect 6644 29155 6696 29164
rect 6644 29121 6678 29155
rect 6678 29121 6696 29155
rect 6644 29112 6696 29121
rect 11796 29189 11805 29223
rect 11805 29189 11839 29223
rect 11839 29189 11848 29223
rect 11796 29180 11848 29189
rect 11336 29112 11388 29164
rect 12164 29257 12173 29291
rect 12173 29257 12207 29291
rect 12207 29257 12216 29291
rect 12164 29248 12216 29257
rect 12716 29248 12768 29300
rect 12256 29180 12308 29232
rect 9588 29044 9640 29096
rect 11980 29155 12032 29164
rect 11980 29121 11994 29155
rect 11994 29121 12028 29155
rect 12028 29121 12032 29155
rect 11980 29112 12032 29121
rect 12164 29112 12216 29164
rect 15200 29248 15252 29300
rect 17592 29291 17644 29300
rect 17592 29257 17601 29291
rect 17601 29257 17635 29291
rect 17635 29257 17644 29291
rect 17592 29248 17644 29257
rect 20904 29248 20956 29300
rect 21272 29248 21324 29300
rect 24032 29248 24084 29300
rect 14004 29180 14056 29232
rect 15292 29180 15344 29232
rect 20628 29223 20680 29232
rect 20628 29189 20637 29223
rect 20637 29189 20671 29223
rect 20671 29189 20680 29223
rect 20628 29180 20680 29189
rect 14924 29112 14976 29164
rect 17316 29112 17368 29164
rect 20076 29112 20128 29164
rect 21088 29180 21140 29232
rect 21824 29180 21876 29232
rect 22652 29112 22704 29164
rect 24952 29180 25004 29232
rect 29276 29180 29328 29232
rect 23296 29112 23348 29164
rect 29092 29155 29144 29164
rect 29092 29121 29101 29155
rect 29101 29121 29135 29155
rect 29135 29121 29144 29155
rect 29092 29112 29144 29121
rect 30840 29155 30892 29164
rect 30840 29121 30858 29155
rect 30858 29121 30892 29155
rect 30840 29112 30892 29121
rect 32496 29112 32548 29164
rect 33508 29155 33560 29164
rect 33508 29121 33517 29155
rect 33517 29121 33551 29155
rect 33551 29121 33560 29155
rect 33508 29112 33560 29121
rect 10508 28976 10560 29028
rect 7288 28908 7340 28960
rect 9680 28908 9732 28960
rect 12256 28976 12308 29028
rect 20260 28976 20312 29028
rect 22192 28976 22244 29028
rect 24492 28976 24544 29028
rect 26240 28976 26292 29028
rect 29920 28976 29972 29028
rect 11888 28908 11940 28960
rect 15016 28908 15068 28960
rect 17408 28908 17460 28960
rect 20996 28951 21048 28960
rect 20996 28917 21005 28951
rect 21005 28917 21039 28951
rect 21039 28917 21048 28951
rect 20996 28908 21048 28917
rect 21548 28908 21600 28960
rect 25780 28908 25832 28960
rect 28724 28951 28776 28960
rect 28724 28917 28733 28951
rect 28733 28917 28767 28951
rect 28767 28917 28776 28951
rect 28724 28908 28776 28917
rect 32128 28951 32180 28960
rect 32128 28917 32137 28951
rect 32137 28917 32171 28951
rect 32171 28917 32180 28951
rect 32128 28908 32180 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 6644 28704 6696 28756
rect 5172 28636 5224 28688
rect 16212 28747 16264 28756
rect 8116 28636 8168 28688
rect 3424 28500 3476 28552
rect 5356 28500 5408 28552
rect 1768 28432 1820 28484
rect 2228 28364 2280 28416
rect 3240 28432 3292 28484
rect 5172 28364 5224 28416
rect 5448 28407 5500 28416
rect 5448 28373 5457 28407
rect 5457 28373 5491 28407
rect 5491 28373 5500 28407
rect 5448 28364 5500 28373
rect 7012 28543 7064 28552
rect 7012 28509 7021 28543
rect 7021 28509 7055 28543
rect 7055 28509 7064 28543
rect 7012 28500 7064 28509
rect 7288 28500 7340 28552
rect 7840 28543 7892 28552
rect 7840 28509 7849 28543
rect 7849 28509 7883 28543
rect 7883 28509 7892 28543
rect 7840 28500 7892 28509
rect 9680 28636 9732 28688
rect 16212 28713 16221 28747
rect 16221 28713 16255 28747
rect 16255 28713 16264 28747
rect 16212 28704 16264 28713
rect 22652 28704 22704 28756
rect 27620 28704 27672 28756
rect 28264 28747 28316 28756
rect 28264 28713 28273 28747
rect 28273 28713 28307 28747
rect 28307 28713 28316 28747
rect 28264 28704 28316 28713
rect 32496 28704 32548 28756
rect 12440 28636 12492 28688
rect 14648 28636 14700 28688
rect 17316 28679 17368 28688
rect 17316 28645 17325 28679
rect 17325 28645 17359 28679
rect 17359 28645 17368 28679
rect 17316 28636 17368 28645
rect 21088 28611 21140 28620
rect 12532 28543 12584 28552
rect 7380 28432 7432 28484
rect 9128 28432 9180 28484
rect 10508 28432 10560 28484
rect 11060 28432 11112 28484
rect 11796 28432 11848 28484
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 12716 28500 12768 28552
rect 15292 28500 15344 28552
rect 16580 28543 16632 28552
rect 15568 28475 15620 28484
rect 15568 28441 15577 28475
rect 15577 28441 15611 28475
rect 15611 28441 15620 28475
rect 15568 28432 15620 28441
rect 16580 28509 16589 28543
rect 16589 28509 16623 28543
rect 16623 28509 16632 28543
rect 16580 28500 16632 28509
rect 21088 28577 21097 28611
rect 21097 28577 21131 28611
rect 21131 28577 21140 28611
rect 21088 28568 21140 28577
rect 22376 28568 22428 28620
rect 22744 28611 22796 28620
rect 22744 28577 22753 28611
rect 22753 28577 22787 28611
rect 22787 28577 22796 28611
rect 22744 28568 22796 28577
rect 17960 28500 18012 28552
rect 18052 28500 18104 28552
rect 21824 28500 21876 28552
rect 8944 28407 8996 28416
rect 8944 28373 8953 28407
rect 8953 28373 8987 28407
rect 8987 28373 8996 28407
rect 8944 28364 8996 28373
rect 11336 28407 11388 28416
rect 11336 28373 11345 28407
rect 11345 28373 11379 28407
rect 11379 28373 11388 28407
rect 11336 28364 11388 28373
rect 12808 28407 12860 28416
rect 12808 28373 12817 28407
rect 12817 28373 12851 28407
rect 12851 28373 12860 28407
rect 12808 28364 12860 28373
rect 17868 28432 17920 28484
rect 20628 28432 20680 28484
rect 16672 28364 16724 28416
rect 16948 28364 17000 28416
rect 20076 28364 20128 28416
rect 23204 28407 23256 28416
rect 23204 28373 23213 28407
rect 23213 28373 23247 28407
rect 23247 28373 23256 28407
rect 23204 28364 23256 28373
rect 23848 28543 23900 28552
rect 23848 28509 23857 28543
rect 23857 28509 23891 28543
rect 23891 28509 23900 28543
rect 23848 28500 23900 28509
rect 28172 28500 28224 28552
rect 24308 28432 24360 28484
rect 24860 28432 24912 28484
rect 25872 28432 25924 28484
rect 26240 28432 26292 28484
rect 28724 28543 28776 28552
rect 28724 28509 28733 28543
rect 28733 28509 28767 28543
rect 28767 28509 28776 28543
rect 28724 28500 28776 28509
rect 28908 28543 28960 28552
rect 28908 28509 28917 28543
rect 28917 28509 28951 28543
rect 28951 28509 28960 28543
rect 28908 28500 28960 28509
rect 30380 28500 30432 28552
rect 30656 28636 30708 28688
rect 30564 28543 30616 28552
rect 30564 28509 30573 28543
rect 30573 28509 30607 28543
rect 30607 28509 30616 28543
rect 30564 28500 30616 28509
rect 30748 28500 30800 28552
rect 29000 28432 29052 28484
rect 23756 28364 23808 28416
rect 25688 28364 25740 28416
rect 27344 28364 27396 28416
rect 30472 28364 30524 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 3240 28203 3292 28212
rect 3240 28169 3249 28203
rect 3249 28169 3283 28203
rect 3283 28169 3292 28203
rect 3240 28160 3292 28169
rect 7012 28160 7064 28212
rect 8116 28160 8168 28212
rect 5448 28092 5500 28144
rect 9588 28160 9640 28212
rect 10324 28135 10376 28144
rect 1768 28067 1820 28076
rect 1768 28033 1777 28067
rect 1777 28033 1811 28067
rect 1811 28033 1820 28067
rect 1768 28024 1820 28033
rect 2320 28024 2372 28076
rect 2872 28067 2924 28076
rect 2872 28033 2881 28067
rect 2881 28033 2915 28067
rect 2915 28033 2924 28067
rect 2872 28024 2924 28033
rect 5356 28024 5408 28076
rect 5632 28067 5684 28076
rect 5632 28033 5641 28067
rect 5641 28033 5675 28067
rect 5675 28033 5684 28067
rect 5632 28024 5684 28033
rect 6736 28024 6788 28076
rect 7104 27956 7156 28008
rect 8208 28024 8260 28076
rect 9128 28067 9180 28076
rect 9128 28033 9137 28067
rect 9137 28033 9171 28067
rect 9171 28033 9180 28067
rect 10324 28101 10333 28135
rect 10333 28101 10367 28135
rect 10367 28101 10376 28135
rect 10324 28092 10376 28101
rect 9128 28024 9180 28033
rect 10140 28067 10192 28076
rect 10140 28033 10149 28067
rect 10149 28033 10183 28067
rect 10183 28033 10192 28067
rect 10140 28024 10192 28033
rect 10416 28067 10468 28076
rect 10416 28033 10425 28067
rect 10425 28033 10459 28067
rect 10459 28033 10468 28067
rect 10416 28024 10468 28033
rect 15292 28160 15344 28212
rect 17868 28203 17920 28212
rect 17868 28169 17877 28203
rect 17877 28169 17911 28203
rect 17911 28169 17920 28203
rect 17868 28160 17920 28169
rect 20628 28203 20680 28212
rect 20628 28169 20637 28203
rect 20637 28169 20671 28203
rect 20671 28169 20680 28203
rect 20628 28160 20680 28169
rect 11152 28092 11204 28144
rect 11796 28092 11848 28144
rect 12164 28092 12216 28144
rect 10232 27956 10284 28008
rect 10324 27888 10376 27940
rect 11888 27956 11940 28008
rect 12716 28024 12768 28076
rect 13268 28067 13320 28076
rect 13268 28033 13277 28067
rect 13277 28033 13311 28067
rect 13311 28033 13320 28067
rect 13268 28024 13320 28033
rect 14096 27956 14148 28008
rect 17132 28092 17184 28144
rect 14740 28024 14792 28076
rect 15936 28024 15988 28076
rect 17960 28092 18012 28144
rect 17408 28067 17460 28076
rect 17408 28033 17417 28067
rect 17417 28033 17451 28067
rect 17451 28033 17460 28067
rect 17408 28024 17460 28033
rect 6828 27820 6880 27872
rect 7932 27820 7984 27872
rect 12256 27863 12308 27872
rect 12256 27829 12265 27863
rect 12265 27829 12299 27863
rect 12299 27829 12308 27863
rect 12256 27820 12308 27829
rect 12992 27820 13044 27872
rect 16580 27956 16632 28008
rect 15476 27888 15528 27940
rect 18052 27820 18104 27872
rect 18880 28024 18932 28076
rect 20904 28067 20956 28076
rect 20904 28033 20913 28067
rect 20913 28033 20947 28067
rect 20947 28033 20956 28067
rect 20904 28024 20956 28033
rect 22100 28160 22152 28212
rect 25228 28203 25280 28212
rect 25228 28169 25237 28203
rect 25237 28169 25271 28203
rect 25271 28169 25280 28203
rect 25228 28160 25280 28169
rect 25780 28160 25832 28212
rect 27344 28160 27396 28212
rect 27804 28160 27856 28212
rect 28172 28203 28224 28212
rect 28172 28169 28181 28203
rect 28181 28169 28215 28203
rect 28215 28169 28224 28203
rect 28172 28160 28224 28169
rect 22192 28135 22244 28144
rect 22192 28101 22201 28135
rect 22201 28101 22235 28135
rect 22235 28101 22244 28135
rect 22192 28092 22244 28101
rect 22376 28135 22428 28144
rect 22376 28101 22385 28135
rect 22385 28101 22419 28135
rect 22419 28101 22428 28135
rect 22376 28092 22428 28101
rect 23204 28092 23256 28144
rect 23756 28092 23808 28144
rect 21088 28067 21140 28076
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 21272 28067 21324 28076
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 26424 28092 26476 28144
rect 21272 28024 21324 28033
rect 21548 27956 21600 28008
rect 22836 27999 22888 28008
rect 22836 27965 22845 27999
rect 22845 27965 22879 27999
rect 22879 27965 22888 27999
rect 22836 27956 22888 27965
rect 25688 28067 25740 28076
rect 25688 28033 25697 28067
rect 25697 28033 25731 28067
rect 25731 28033 25740 28067
rect 25688 28024 25740 28033
rect 19984 27820 20036 27872
rect 24400 27888 24452 27940
rect 24584 27820 24636 27872
rect 25780 27956 25832 28008
rect 26148 27956 26200 28008
rect 28080 28024 28132 28076
rect 28908 28160 28960 28212
rect 29000 28160 29052 28212
rect 30656 28160 30708 28212
rect 30380 28092 30432 28144
rect 29184 28024 29236 28076
rect 32128 28092 32180 28144
rect 30840 28067 30892 28076
rect 30840 28033 30849 28067
rect 30849 28033 30883 28067
rect 30883 28033 30892 28067
rect 30840 28024 30892 28033
rect 32496 28024 32548 28076
rect 33508 28067 33560 28076
rect 33508 28033 33517 28067
rect 33517 28033 33551 28067
rect 33551 28033 33560 28067
rect 33508 28024 33560 28033
rect 29368 27956 29420 28008
rect 30380 27956 30432 28008
rect 67640 27931 67692 27940
rect 67640 27897 67649 27931
rect 67649 27897 67683 27931
rect 67683 27897 67692 27931
rect 67640 27888 67692 27897
rect 31024 27820 31076 27872
rect 32128 27863 32180 27872
rect 32128 27829 32137 27863
rect 32137 27829 32171 27863
rect 32171 27829 32180 27863
rect 32128 27820 32180 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 5632 27616 5684 27668
rect 10784 27616 10836 27668
rect 11336 27616 11388 27668
rect 14740 27659 14792 27668
rect 2596 27548 2648 27600
rect 3332 27548 3384 27600
rect 10324 27591 10376 27600
rect 10324 27557 10333 27591
rect 10333 27557 10367 27591
rect 10367 27557 10376 27591
rect 10324 27548 10376 27557
rect 11244 27548 11296 27600
rect 14740 27625 14749 27659
rect 14749 27625 14783 27659
rect 14783 27625 14792 27659
rect 14740 27616 14792 27625
rect 17500 27616 17552 27668
rect 20444 27659 20496 27668
rect 20444 27625 20453 27659
rect 20453 27625 20487 27659
rect 20487 27625 20496 27659
rect 20444 27616 20496 27625
rect 20904 27616 20956 27668
rect 24308 27616 24360 27668
rect 18144 27548 18196 27600
rect 2228 27455 2280 27464
rect 2228 27421 2237 27455
rect 2237 27421 2271 27455
rect 2271 27421 2280 27455
rect 2228 27412 2280 27421
rect 2872 27480 2924 27532
rect 2596 27412 2648 27464
rect 7748 27455 7800 27464
rect 6552 27344 6604 27396
rect 7748 27421 7757 27455
rect 7757 27421 7791 27455
rect 7791 27421 7800 27455
rect 7748 27412 7800 27421
rect 7932 27455 7984 27464
rect 7932 27421 7941 27455
rect 7941 27421 7975 27455
rect 7975 27421 7984 27455
rect 7932 27412 7984 27421
rect 8024 27455 8076 27464
rect 8024 27421 8033 27455
rect 8033 27421 8067 27455
rect 8067 27421 8076 27455
rect 8024 27412 8076 27421
rect 10508 27412 10560 27464
rect 10876 27455 10928 27464
rect 10876 27421 10885 27455
rect 10885 27421 10919 27455
rect 10919 27421 10928 27455
rect 10876 27412 10928 27421
rect 15568 27480 15620 27532
rect 16580 27480 16632 27532
rect 17776 27480 17828 27532
rect 25136 27548 25188 27600
rect 26148 27591 26200 27600
rect 26148 27557 26157 27591
rect 26157 27557 26191 27591
rect 26191 27557 26200 27591
rect 26148 27548 26200 27557
rect 27712 27548 27764 27600
rect 32496 27548 32548 27600
rect 22100 27480 22152 27532
rect 11888 27412 11940 27464
rect 12992 27412 13044 27464
rect 14188 27412 14240 27464
rect 11152 27387 11204 27396
rect 11152 27353 11161 27387
rect 11161 27353 11195 27387
rect 11195 27353 11204 27387
rect 11152 27344 11204 27353
rect 2320 27276 2372 27328
rect 7380 27276 7432 27328
rect 8024 27276 8076 27328
rect 8208 27276 8260 27328
rect 12900 27344 12952 27396
rect 12072 27276 12124 27328
rect 14096 27276 14148 27328
rect 15200 27412 15252 27464
rect 16304 27412 16356 27464
rect 17960 27412 18012 27464
rect 18512 27455 18564 27464
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 22008 27455 22060 27464
rect 16580 27344 16632 27396
rect 17592 27344 17644 27396
rect 19432 27387 19484 27396
rect 19432 27353 19441 27387
rect 19441 27353 19475 27387
rect 19475 27353 19484 27387
rect 19432 27344 19484 27353
rect 22008 27421 22017 27455
rect 22017 27421 22051 27455
rect 22051 27421 22060 27455
rect 22008 27412 22060 27421
rect 27988 27480 28040 27532
rect 25596 27412 25648 27464
rect 28080 27455 28132 27464
rect 28080 27421 28089 27455
rect 28089 27421 28123 27455
rect 28123 27421 28132 27455
rect 28080 27412 28132 27421
rect 30288 27455 30340 27464
rect 30288 27421 30297 27455
rect 30297 27421 30331 27455
rect 30331 27421 30340 27455
rect 30288 27412 30340 27421
rect 30564 27480 30616 27532
rect 24584 27387 24636 27396
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 24860 27344 24912 27396
rect 26148 27344 26200 27396
rect 26332 27344 26384 27396
rect 30748 27412 30800 27464
rect 18236 27276 18288 27328
rect 25228 27276 25280 27328
rect 25688 27276 25740 27328
rect 26700 27319 26752 27328
rect 26700 27285 26709 27319
rect 26709 27285 26743 27319
rect 26743 27285 26752 27319
rect 26700 27276 26752 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 6552 27115 6604 27124
rect 6552 27081 6561 27115
rect 6561 27081 6595 27115
rect 6595 27081 6604 27115
rect 6552 27072 6604 27081
rect 10232 27072 10284 27124
rect 10876 27115 10928 27124
rect 10140 27004 10192 27056
rect 10876 27081 10885 27115
rect 10885 27081 10919 27115
rect 10919 27081 10928 27115
rect 10876 27072 10928 27081
rect 16580 27072 16632 27124
rect 20444 27115 20496 27124
rect 20444 27081 20453 27115
rect 20453 27081 20487 27115
rect 20487 27081 20496 27115
rect 20444 27072 20496 27081
rect 23572 27072 23624 27124
rect 29184 27072 29236 27124
rect 29368 27115 29420 27124
rect 29368 27081 29377 27115
rect 29377 27081 29411 27115
rect 29411 27081 29420 27115
rect 29368 27072 29420 27081
rect 30288 27072 30340 27124
rect 18144 27047 18196 27056
rect 2320 26979 2372 26988
rect 2320 26945 2329 26979
rect 2329 26945 2363 26979
rect 2363 26945 2372 26979
rect 2320 26936 2372 26945
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 3424 26979 3476 26988
rect 2872 26868 2924 26920
rect 3424 26945 3433 26979
rect 3433 26945 3467 26979
rect 3467 26945 3476 26979
rect 3424 26936 3476 26945
rect 7012 26979 7064 26988
rect 7012 26945 7021 26979
rect 7021 26945 7055 26979
rect 7055 26945 7064 26979
rect 7012 26936 7064 26945
rect 7288 26936 7340 26988
rect 9680 26936 9732 26988
rect 7380 26868 7432 26920
rect 7472 26868 7524 26920
rect 10692 26979 10744 26988
rect 10692 26945 10701 26979
rect 10701 26945 10735 26979
rect 10735 26945 10744 26979
rect 18144 27013 18153 27047
rect 18153 27013 18187 27047
rect 18187 27013 18196 27047
rect 18144 27004 18196 27013
rect 20996 27004 21048 27056
rect 24400 27004 24452 27056
rect 25136 27004 25188 27056
rect 10692 26936 10744 26945
rect 14004 26936 14056 26988
rect 14096 26936 14148 26988
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 20168 26936 20220 26988
rect 21180 26936 21232 26988
rect 21824 26979 21876 26988
rect 21824 26945 21833 26979
rect 21833 26945 21867 26979
rect 21867 26945 21876 26979
rect 21824 26936 21876 26945
rect 23204 26936 23256 26988
rect 13636 26868 13688 26920
rect 13912 26911 13964 26920
rect 13912 26877 13921 26911
rect 13921 26877 13955 26911
rect 13955 26877 13964 26911
rect 13912 26868 13964 26877
rect 16304 26868 16356 26920
rect 17868 26868 17920 26920
rect 24032 26936 24084 26988
rect 25228 26979 25280 26988
rect 25228 26945 25237 26979
rect 25237 26945 25271 26979
rect 25271 26945 25280 26979
rect 25228 26936 25280 26945
rect 25780 26979 25832 26988
rect 26332 27004 26384 27056
rect 25780 26945 25795 26979
rect 25795 26945 25829 26979
rect 25829 26945 25832 26979
rect 25780 26936 25832 26945
rect 27620 27004 27672 27056
rect 28172 27004 28224 27056
rect 29092 27004 29144 27056
rect 30840 27004 30892 27056
rect 24860 26868 24912 26920
rect 9128 26800 9180 26852
rect 9496 26800 9548 26852
rect 11888 26800 11940 26852
rect 29920 26936 29972 26988
rect 32128 27004 32180 27056
rect 26332 26868 26384 26920
rect 29644 26868 29696 26920
rect 26608 26800 26660 26852
rect 3700 26732 3752 26784
rect 10416 26732 10468 26784
rect 12900 26775 12952 26784
rect 12900 26741 12909 26775
rect 12909 26741 12943 26775
rect 12943 26741 12952 26775
rect 12900 26732 12952 26741
rect 15200 26732 15252 26784
rect 16028 26732 16080 26784
rect 18052 26732 18104 26784
rect 19248 26732 19300 26784
rect 22652 26732 22704 26784
rect 23388 26732 23440 26784
rect 26424 26732 26476 26784
rect 31024 26732 31076 26784
rect 67640 26775 67692 26784
rect 67640 26741 67649 26775
rect 67649 26741 67683 26775
rect 67683 26741 67692 26775
rect 67640 26732 67692 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 2504 26528 2556 26580
rect 5172 26571 5224 26580
rect 5172 26537 5181 26571
rect 5181 26537 5215 26571
rect 5215 26537 5224 26571
rect 5172 26528 5224 26537
rect 7472 26528 7524 26580
rect 8208 26571 8260 26580
rect 8208 26537 8217 26571
rect 8217 26537 8251 26571
rect 8251 26537 8260 26571
rect 8208 26528 8260 26537
rect 12164 26528 12216 26580
rect 12808 26528 12860 26580
rect 14096 26528 14148 26580
rect 3700 26460 3752 26512
rect 11888 26460 11940 26512
rect 3424 26392 3476 26444
rect 3792 26435 3844 26444
rect 3792 26401 3801 26435
rect 3801 26401 3835 26435
rect 3835 26401 3844 26435
rect 3792 26392 3844 26401
rect 12624 26460 12676 26512
rect 13084 26460 13136 26512
rect 6828 26367 6880 26376
rect 6828 26333 6837 26367
rect 6837 26333 6871 26367
rect 6871 26333 6880 26367
rect 6828 26324 6880 26333
rect 1768 26256 1820 26308
rect 3240 26256 3292 26308
rect 6920 26256 6972 26308
rect 10600 26367 10652 26376
rect 10600 26333 10609 26367
rect 10609 26333 10643 26367
rect 10643 26333 10652 26367
rect 10600 26324 10652 26333
rect 5724 26188 5776 26240
rect 10416 26299 10468 26308
rect 10416 26265 10425 26299
rect 10425 26265 10459 26299
rect 10459 26265 10468 26299
rect 10416 26256 10468 26265
rect 10692 26256 10744 26308
rect 12532 26367 12584 26376
rect 12532 26333 12541 26367
rect 12541 26333 12575 26367
rect 12575 26333 12584 26367
rect 12532 26324 12584 26333
rect 12808 26324 12860 26376
rect 12900 26324 12952 26376
rect 14004 26324 14056 26376
rect 13912 26256 13964 26308
rect 14924 26324 14976 26376
rect 15016 26367 15068 26376
rect 15016 26333 15025 26367
rect 15025 26333 15059 26367
rect 15059 26333 15068 26367
rect 15016 26324 15068 26333
rect 16488 26256 16540 26308
rect 18512 26460 18564 26512
rect 20996 26503 21048 26512
rect 16764 26324 16816 26376
rect 17868 26392 17920 26444
rect 20996 26469 21005 26503
rect 21005 26469 21039 26503
rect 21039 26469 21048 26503
rect 20996 26460 21048 26469
rect 17960 26324 18012 26376
rect 18236 26367 18288 26376
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 22836 26392 22888 26444
rect 19708 26367 19760 26376
rect 19340 26256 19392 26308
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 22744 26324 22796 26376
rect 25780 26528 25832 26580
rect 26608 26571 26660 26580
rect 26608 26537 26617 26571
rect 26617 26537 26651 26571
rect 26651 26537 26660 26571
rect 26608 26528 26660 26537
rect 27712 26571 27764 26580
rect 27712 26537 27721 26571
rect 27721 26537 27755 26571
rect 27755 26537 27764 26571
rect 27712 26528 27764 26537
rect 23388 26460 23440 26512
rect 24400 26503 24452 26512
rect 24400 26469 24409 26503
rect 24409 26469 24443 26503
rect 24443 26469 24452 26503
rect 24400 26460 24452 26469
rect 26700 26460 26752 26512
rect 23756 26392 23808 26444
rect 25780 26435 25832 26444
rect 25780 26401 25789 26435
rect 25789 26401 25823 26435
rect 25823 26401 25832 26435
rect 25780 26392 25832 26401
rect 27712 26392 27764 26444
rect 23572 26367 23624 26376
rect 23572 26333 23601 26367
rect 23601 26333 23624 26367
rect 23572 26324 23624 26333
rect 26056 26324 26108 26376
rect 30748 26392 30800 26444
rect 30656 26367 30708 26376
rect 12440 26188 12492 26240
rect 12624 26188 12676 26240
rect 16304 26188 16356 26240
rect 18788 26188 18840 26240
rect 19708 26188 19760 26240
rect 22100 26299 22152 26308
rect 22100 26265 22118 26299
rect 22118 26265 22152 26299
rect 22100 26256 22152 26265
rect 26148 26256 26200 26308
rect 26424 26299 26476 26308
rect 26424 26265 26433 26299
rect 26433 26265 26467 26299
rect 26467 26265 26476 26299
rect 26424 26256 26476 26265
rect 27068 26299 27120 26308
rect 27068 26265 27077 26299
rect 27077 26265 27111 26299
rect 27111 26265 27120 26299
rect 27068 26256 27120 26265
rect 29736 26256 29788 26308
rect 30656 26333 30665 26367
rect 30665 26333 30699 26367
rect 30699 26333 30708 26367
rect 30656 26324 30708 26333
rect 30840 26367 30892 26376
rect 30840 26333 30849 26367
rect 30849 26333 30883 26367
rect 30883 26333 30892 26367
rect 30840 26324 30892 26333
rect 31024 26367 31076 26376
rect 31024 26333 31033 26367
rect 31033 26333 31067 26367
rect 31067 26333 31076 26367
rect 33508 26392 33560 26444
rect 31024 26324 31076 26333
rect 34060 26324 34112 26376
rect 31208 26256 31260 26308
rect 24768 26188 24820 26240
rect 29552 26231 29604 26240
rect 29552 26197 29561 26231
rect 29561 26197 29595 26231
rect 29595 26197 29604 26231
rect 29552 26188 29604 26197
rect 31852 26188 31904 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 3240 26027 3292 26036
rect 3240 25993 3249 26027
rect 3249 25993 3283 26027
rect 3283 25993 3292 26027
rect 3240 25984 3292 25993
rect 6828 25984 6880 26036
rect 12440 25984 12492 26036
rect 13084 25984 13136 26036
rect 15936 25984 15988 26036
rect 22100 25984 22152 26036
rect 25780 25984 25832 26036
rect 27804 25984 27856 26036
rect 30840 25984 30892 26036
rect 33508 25984 33560 26036
rect 34428 25984 34480 26036
rect 1768 25959 1820 25968
rect 1768 25925 1777 25959
rect 1777 25925 1811 25959
rect 1811 25925 1820 25959
rect 1768 25916 1820 25925
rect 5172 25916 5224 25968
rect 2320 25848 2372 25900
rect 2872 25891 2924 25900
rect 2872 25857 2881 25891
rect 2881 25857 2915 25891
rect 2915 25857 2924 25891
rect 2872 25848 2924 25857
rect 6644 25891 6696 25900
rect 6644 25857 6653 25891
rect 6653 25857 6687 25891
rect 6687 25857 6696 25891
rect 6644 25848 6696 25857
rect 6828 25891 6880 25900
rect 6828 25857 6837 25891
rect 6837 25857 6871 25891
rect 6871 25857 6880 25891
rect 6828 25848 6880 25857
rect 7012 25891 7064 25900
rect 7012 25857 7021 25891
rect 7021 25857 7055 25891
rect 7055 25857 7064 25891
rect 7012 25848 7064 25857
rect 7748 25848 7800 25900
rect 10692 25916 10744 25968
rect 16028 25916 16080 25968
rect 16856 25916 16908 25968
rect 7380 25780 7432 25832
rect 10232 25712 10284 25764
rect 12624 25848 12676 25900
rect 14004 25848 14056 25900
rect 15016 25891 15068 25900
rect 15016 25857 15025 25891
rect 15025 25857 15059 25891
rect 15059 25857 15068 25891
rect 15016 25848 15068 25857
rect 12532 25780 12584 25832
rect 12992 25780 13044 25832
rect 14832 25823 14884 25832
rect 14832 25789 14841 25823
rect 14841 25789 14875 25823
rect 14875 25789 14884 25823
rect 14832 25780 14884 25789
rect 14004 25712 14056 25764
rect 16672 25848 16724 25900
rect 19340 25848 19392 25900
rect 22468 25891 22520 25900
rect 22468 25857 22477 25891
rect 22477 25857 22511 25891
rect 22511 25857 22520 25891
rect 22468 25848 22520 25857
rect 19248 25823 19300 25832
rect 19248 25789 19257 25823
rect 19257 25789 19291 25823
rect 19291 25789 19300 25823
rect 19248 25780 19300 25789
rect 22008 25780 22060 25832
rect 22652 25891 22704 25900
rect 22652 25857 22661 25891
rect 22661 25857 22695 25891
rect 22695 25857 22704 25891
rect 28080 25916 28132 25968
rect 29552 25959 29604 25968
rect 29552 25925 29586 25959
rect 29586 25925 29604 25959
rect 29552 25916 29604 25925
rect 22652 25848 22704 25857
rect 23756 25848 23808 25900
rect 26240 25848 26292 25900
rect 27988 25891 28040 25900
rect 23296 25823 23348 25832
rect 23296 25789 23305 25823
rect 23305 25789 23339 25823
rect 23339 25789 23348 25823
rect 23296 25780 23348 25789
rect 6920 25644 6972 25696
rect 16212 25644 16264 25696
rect 16396 25644 16448 25696
rect 19432 25644 19484 25696
rect 27988 25857 27997 25891
rect 27997 25857 28031 25891
rect 28031 25857 28040 25891
rect 27988 25848 28040 25857
rect 28172 25848 28224 25900
rect 30656 25848 30708 25900
rect 30932 25848 30984 25900
rect 31852 25848 31904 25900
rect 32496 25891 32548 25900
rect 32496 25857 32505 25891
rect 32505 25857 32539 25891
rect 32539 25857 32548 25891
rect 32496 25848 32548 25857
rect 32680 25891 32732 25900
rect 32680 25857 32689 25891
rect 32689 25857 32723 25891
rect 32723 25857 32732 25891
rect 32680 25848 32732 25857
rect 32864 25891 32916 25900
rect 32864 25857 32873 25891
rect 32873 25857 32907 25891
rect 32907 25857 32916 25891
rect 32864 25848 32916 25857
rect 32956 25780 33008 25832
rect 34704 25848 34756 25900
rect 31576 25644 31628 25696
rect 33140 25687 33192 25696
rect 33140 25653 33149 25687
rect 33149 25653 33183 25687
rect 33183 25653 33192 25687
rect 33140 25644 33192 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 5724 25483 5776 25492
rect 5724 25449 5733 25483
rect 5733 25449 5767 25483
rect 5767 25449 5776 25483
rect 5724 25440 5776 25449
rect 6828 25440 6880 25492
rect 16672 25483 16724 25492
rect 16672 25449 16681 25483
rect 16681 25449 16715 25483
rect 16715 25449 16724 25483
rect 16672 25440 16724 25449
rect 12256 25372 12308 25424
rect 18604 25372 18656 25424
rect 18788 25372 18840 25424
rect 19064 25372 19116 25424
rect 3792 25304 3844 25356
rect 10508 25347 10560 25356
rect 10508 25313 10517 25347
rect 10517 25313 10551 25347
rect 10551 25313 10560 25347
rect 10508 25304 10560 25313
rect 11704 25304 11756 25356
rect 23204 25440 23256 25492
rect 31208 25440 31260 25492
rect 32680 25440 32732 25492
rect 20904 25372 20956 25424
rect 26240 25415 26292 25424
rect 26240 25381 26249 25415
rect 26249 25381 26283 25415
rect 26283 25381 26292 25415
rect 26240 25372 26292 25381
rect 2320 25236 2372 25288
rect 2872 25279 2924 25288
rect 2872 25245 2881 25279
rect 2881 25245 2915 25279
rect 2915 25245 2924 25279
rect 2872 25236 2924 25245
rect 5632 25236 5684 25288
rect 8208 25236 8260 25288
rect 14464 25236 14516 25288
rect 16212 25279 16264 25288
rect 7104 25211 7156 25220
rect 7104 25177 7113 25211
rect 7113 25177 7147 25211
rect 7147 25177 7156 25211
rect 7104 25168 7156 25177
rect 12348 25168 12400 25220
rect 12624 25168 12676 25220
rect 2872 25100 2924 25152
rect 12440 25100 12492 25152
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 13820 25100 13872 25152
rect 14832 25168 14884 25220
rect 16212 25245 16221 25279
rect 16221 25245 16255 25279
rect 16255 25245 16264 25279
rect 16212 25236 16264 25245
rect 16304 25279 16356 25288
rect 16304 25245 16313 25279
rect 16313 25245 16347 25279
rect 16347 25245 16356 25279
rect 16304 25236 16356 25245
rect 16856 25236 16908 25288
rect 17592 25279 17644 25288
rect 17592 25245 17601 25279
rect 17601 25245 17635 25279
rect 17635 25245 17644 25279
rect 17592 25236 17644 25245
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 21916 25236 21968 25288
rect 23664 25304 23716 25356
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 22652 25279 22704 25288
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 26056 25304 26108 25356
rect 16764 25168 16816 25220
rect 19340 25168 19392 25220
rect 20536 25168 20588 25220
rect 25228 25236 25280 25288
rect 25688 25236 25740 25288
rect 28172 25347 28224 25356
rect 28172 25313 28181 25347
rect 28181 25313 28215 25347
rect 28215 25313 28224 25347
rect 28172 25304 28224 25313
rect 30748 25304 30800 25356
rect 34428 25304 34480 25356
rect 29552 25279 29604 25288
rect 23480 25211 23532 25220
rect 23480 25177 23489 25211
rect 23489 25177 23523 25211
rect 23523 25177 23532 25211
rect 23480 25168 23532 25177
rect 24032 25168 24084 25220
rect 29552 25245 29561 25279
rect 29561 25245 29595 25279
rect 29595 25245 29604 25279
rect 29552 25236 29604 25245
rect 33140 25236 33192 25288
rect 68100 25279 68152 25288
rect 68100 25245 68109 25279
rect 68109 25245 68143 25279
rect 68143 25245 68152 25279
rect 68100 25236 68152 25245
rect 26332 25168 26384 25220
rect 31576 25168 31628 25220
rect 31760 25168 31812 25220
rect 32680 25168 32732 25220
rect 14372 25100 14424 25152
rect 18144 25100 18196 25152
rect 23572 25100 23624 25152
rect 25504 25100 25556 25152
rect 34704 25100 34756 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 2872 24939 2924 24948
rect 2872 24905 2881 24939
rect 2881 24905 2915 24939
rect 2915 24905 2924 24939
rect 2872 24896 2924 24905
rect 1768 24828 1820 24880
rect 4712 24760 4764 24812
rect 5724 24692 5776 24744
rect 6736 24760 6788 24812
rect 13452 24828 13504 24880
rect 13912 24896 13964 24948
rect 22560 24896 22612 24948
rect 24768 24939 24820 24948
rect 24768 24905 24777 24939
rect 24777 24905 24811 24939
rect 24811 24905 24820 24939
rect 24768 24896 24820 24905
rect 25136 24896 25188 24948
rect 25780 24896 25832 24948
rect 7564 24692 7616 24744
rect 4804 24624 4856 24676
rect 4712 24556 4764 24608
rect 7104 24624 7156 24676
rect 7380 24624 7432 24676
rect 7748 24692 7800 24744
rect 11980 24803 12032 24812
rect 11980 24769 11989 24803
rect 11989 24769 12023 24803
rect 12023 24769 12032 24803
rect 12164 24803 12216 24812
rect 11980 24760 12032 24769
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 16948 24828 17000 24880
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 12348 24692 12400 24744
rect 13360 24692 13412 24744
rect 14832 24760 14884 24812
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 19432 24803 19484 24812
rect 14188 24692 14240 24744
rect 14924 24692 14976 24744
rect 16120 24735 16172 24744
rect 16120 24701 16129 24735
rect 16129 24701 16163 24735
rect 16163 24701 16172 24735
rect 16120 24692 16172 24701
rect 17500 24692 17552 24744
rect 17868 24692 17920 24744
rect 6644 24556 6696 24608
rect 9588 24556 9640 24608
rect 14464 24556 14516 24608
rect 18144 24624 18196 24676
rect 19432 24769 19441 24803
rect 19441 24769 19475 24803
rect 19475 24769 19484 24803
rect 19432 24760 19484 24769
rect 19984 24803 20036 24812
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 20352 24760 20404 24812
rect 21088 24803 21140 24812
rect 21088 24769 21097 24803
rect 21097 24769 21131 24803
rect 21131 24769 21140 24803
rect 21088 24760 21140 24769
rect 22008 24803 22060 24812
rect 19340 24692 19392 24744
rect 22008 24769 22017 24803
rect 22017 24769 22051 24803
rect 22051 24769 22060 24803
rect 22008 24760 22060 24769
rect 19524 24624 19576 24676
rect 20904 24624 20956 24676
rect 23480 24760 23532 24812
rect 23572 24760 23624 24812
rect 24216 24803 24268 24812
rect 24216 24769 24225 24803
rect 24225 24769 24259 24803
rect 24259 24769 24268 24803
rect 24216 24760 24268 24769
rect 25228 24760 25280 24812
rect 25504 24803 25556 24812
rect 25504 24769 25513 24803
rect 25513 24769 25547 24803
rect 25547 24769 25556 24803
rect 25504 24760 25556 24769
rect 26240 24828 26292 24880
rect 27160 24803 27212 24812
rect 24216 24624 24268 24676
rect 25504 24624 25556 24676
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 25780 24692 25832 24744
rect 26332 24692 26384 24744
rect 27344 24803 27396 24812
rect 27344 24769 27353 24803
rect 27353 24769 27387 24803
rect 27387 24769 27396 24803
rect 27344 24760 27396 24769
rect 27712 24760 27764 24812
rect 28356 24760 28408 24812
rect 30932 24896 30984 24948
rect 30288 24803 30340 24812
rect 30288 24769 30297 24803
rect 30297 24769 30331 24803
rect 30331 24769 30340 24803
rect 30288 24760 30340 24769
rect 32864 24896 32916 24948
rect 32496 24760 32548 24812
rect 33140 24760 33192 24812
rect 32864 24692 32916 24744
rect 33416 24803 33468 24812
rect 33416 24769 33425 24803
rect 33425 24769 33459 24803
rect 33459 24769 33468 24803
rect 33416 24760 33468 24769
rect 34428 24760 34480 24812
rect 31760 24624 31812 24676
rect 22008 24556 22060 24608
rect 27528 24556 27580 24608
rect 32956 24556 33008 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 1768 24395 1820 24404
rect 1768 24361 1777 24395
rect 1777 24361 1811 24395
rect 1811 24361 1820 24395
rect 1768 24352 1820 24361
rect 2964 24352 3016 24404
rect 11980 24352 12032 24404
rect 13728 24352 13780 24404
rect 14832 24395 14884 24404
rect 14832 24361 14841 24395
rect 14841 24361 14875 24395
rect 14875 24361 14884 24395
rect 14832 24352 14884 24361
rect 14924 24352 14976 24404
rect 6644 24284 6696 24336
rect 14556 24284 14608 24336
rect 16488 24284 16540 24336
rect 23296 24352 23348 24404
rect 27160 24352 27212 24404
rect 5172 24216 5224 24268
rect 2504 24080 2556 24132
rect 2872 24080 2924 24132
rect 3332 24148 3384 24200
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 2688 24012 2740 24064
rect 7840 24148 7892 24200
rect 9588 24191 9640 24200
rect 9588 24157 9597 24191
rect 9597 24157 9631 24191
rect 9631 24157 9640 24191
rect 9588 24148 9640 24157
rect 10232 24191 10284 24200
rect 10232 24157 10241 24191
rect 10241 24157 10275 24191
rect 10275 24157 10284 24191
rect 10232 24148 10284 24157
rect 6644 24080 6696 24132
rect 4436 24055 4488 24064
rect 4436 24021 4445 24055
rect 4445 24021 4479 24055
rect 4479 24021 4488 24055
rect 4436 24012 4488 24021
rect 6736 24012 6788 24064
rect 10140 24080 10192 24132
rect 17500 24216 17552 24268
rect 10600 24191 10652 24200
rect 10600 24157 10609 24191
rect 10609 24157 10643 24191
rect 10643 24157 10652 24191
rect 10600 24148 10652 24157
rect 12440 24148 12492 24200
rect 13360 24148 13412 24200
rect 14372 24191 14424 24200
rect 14372 24157 14381 24191
rect 14381 24157 14415 24191
rect 14415 24157 14424 24191
rect 14372 24148 14424 24157
rect 12624 24080 12676 24132
rect 13176 24080 13228 24132
rect 13912 24080 13964 24132
rect 15200 24148 15252 24200
rect 17592 24148 17644 24200
rect 17960 24148 18012 24200
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 16856 24080 16908 24132
rect 18236 24080 18288 24132
rect 19156 24080 19208 24132
rect 22284 24284 22336 24336
rect 23848 24284 23900 24336
rect 25688 24284 25740 24336
rect 21824 24216 21876 24268
rect 20904 24148 20956 24200
rect 22652 24148 22704 24200
rect 24216 24216 24268 24268
rect 27804 24259 27856 24268
rect 27804 24225 27813 24259
rect 27813 24225 27847 24259
rect 27847 24225 27856 24259
rect 27804 24216 27856 24225
rect 23204 24148 23256 24200
rect 23572 24148 23624 24200
rect 24860 24148 24912 24200
rect 27528 24191 27580 24200
rect 27528 24157 27546 24191
rect 27546 24157 27580 24191
rect 28356 24191 28408 24200
rect 27528 24148 27580 24157
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 33140 24395 33192 24404
rect 33140 24361 33149 24395
rect 33149 24361 33183 24395
rect 33183 24361 33192 24395
rect 33140 24352 33192 24361
rect 30564 24284 30616 24336
rect 33416 24284 33468 24336
rect 28908 24216 28960 24268
rect 29460 24216 29512 24268
rect 23756 24080 23808 24132
rect 11152 24012 11204 24064
rect 11520 24012 11572 24064
rect 17592 24012 17644 24064
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 19340 24012 19392 24064
rect 19984 24012 20036 24064
rect 20352 24055 20404 24064
rect 20352 24021 20361 24055
rect 20361 24021 20395 24055
rect 20395 24021 20404 24055
rect 20352 24012 20404 24021
rect 24308 24012 24360 24064
rect 28172 24080 28224 24132
rect 31944 24148 31996 24200
rect 34428 24148 34480 24200
rect 68100 24191 68152 24200
rect 68100 24157 68109 24191
rect 68109 24157 68143 24191
rect 68143 24157 68152 24191
rect 68100 24148 68152 24157
rect 30288 24080 30340 24132
rect 27344 24012 27396 24064
rect 30564 24012 30616 24064
rect 31300 24012 31352 24064
rect 31668 24080 31720 24132
rect 32220 24055 32272 24064
rect 32220 24021 32229 24055
rect 32229 24021 32263 24055
rect 32263 24021 32272 24055
rect 32220 24012 32272 24021
rect 32772 24123 32824 24132
rect 32772 24089 32781 24123
rect 32781 24089 32815 24123
rect 32815 24089 32824 24123
rect 32956 24123 33008 24132
rect 32772 24080 32824 24089
rect 32956 24089 32965 24123
rect 32965 24089 32999 24123
rect 32999 24089 33008 24123
rect 32956 24080 33008 24089
rect 36728 24012 36780 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 5632 23808 5684 23860
rect 4436 23740 4488 23792
rect 7104 23808 7156 23860
rect 2320 23715 2372 23724
rect 2320 23681 2329 23715
rect 2329 23681 2363 23715
rect 2363 23681 2372 23715
rect 2320 23672 2372 23681
rect 3792 23715 3844 23724
rect 3792 23681 3801 23715
rect 3801 23681 3835 23715
rect 3835 23681 3844 23715
rect 3792 23672 3844 23681
rect 6828 23672 6880 23724
rect 7472 23672 7524 23724
rect 9588 23672 9640 23724
rect 10140 23715 10192 23724
rect 10140 23681 10149 23715
rect 10149 23681 10183 23715
rect 10183 23681 10192 23715
rect 10140 23672 10192 23681
rect 5172 23579 5224 23588
rect 5172 23545 5181 23579
rect 5181 23545 5215 23579
rect 5215 23545 5224 23579
rect 5172 23536 5224 23545
rect 5632 23536 5684 23588
rect 3148 23511 3200 23520
rect 3148 23477 3157 23511
rect 3157 23477 3191 23511
rect 3191 23477 3200 23511
rect 3148 23468 3200 23477
rect 6920 23511 6972 23520
rect 6920 23477 6929 23511
rect 6929 23477 6963 23511
rect 6963 23477 6972 23511
rect 6920 23468 6972 23477
rect 10600 23672 10652 23724
rect 11612 23468 11664 23520
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 14648 23808 14700 23860
rect 15200 23808 15252 23860
rect 16028 23808 16080 23860
rect 12164 23536 12216 23588
rect 12348 23715 12400 23724
rect 12348 23681 12362 23715
rect 12362 23681 12396 23715
rect 12396 23681 12400 23715
rect 13360 23715 13412 23724
rect 12348 23672 12400 23681
rect 13360 23681 13369 23715
rect 13369 23681 13403 23715
rect 13403 23681 13412 23715
rect 13360 23672 13412 23681
rect 13544 23715 13596 23724
rect 13544 23681 13553 23715
rect 13553 23681 13587 23715
rect 13587 23681 13596 23715
rect 13544 23672 13596 23681
rect 13912 23740 13964 23792
rect 19432 23808 19484 23860
rect 15476 23672 15528 23724
rect 16764 23672 16816 23724
rect 17408 23715 17460 23724
rect 17408 23681 17417 23715
rect 17417 23681 17451 23715
rect 17451 23681 17460 23715
rect 17408 23672 17460 23681
rect 16120 23647 16172 23656
rect 16120 23613 16129 23647
rect 16129 23613 16163 23647
rect 16163 23613 16172 23647
rect 16120 23604 16172 23613
rect 17592 23715 17644 23724
rect 17592 23681 17601 23715
rect 17601 23681 17635 23715
rect 17635 23681 17644 23715
rect 22284 23851 22336 23860
rect 22284 23817 22293 23851
rect 22293 23817 22327 23851
rect 22327 23817 22336 23851
rect 22284 23808 22336 23817
rect 19984 23740 20036 23792
rect 20352 23740 20404 23792
rect 20996 23740 21048 23792
rect 23480 23808 23532 23860
rect 24860 23808 24912 23860
rect 28172 23851 28224 23860
rect 28172 23817 28181 23851
rect 28181 23817 28215 23851
rect 28215 23817 28224 23851
rect 28172 23808 28224 23817
rect 17592 23672 17644 23681
rect 18236 23715 18288 23724
rect 18236 23681 18245 23715
rect 18245 23681 18279 23715
rect 18279 23681 18288 23715
rect 18236 23672 18288 23681
rect 21180 23672 21232 23724
rect 19248 23604 19300 23656
rect 17500 23536 17552 23588
rect 12532 23511 12584 23520
rect 12532 23477 12541 23511
rect 12541 23477 12575 23511
rect 12575 23477 12584 23511
rect 12532 23468 12584 23477
rect 15200 23468 15252 23520
rect 16120 23468 16172 23520
rect 21732 23604 21784 23656
rect 23664 23672 23716 23724
rect 24308 23672 24360 23724
rect 26976 23740 27028 23792
rect 27804 23740 27856 23792
rect 31760 23808 31812 23860
rect 32496 23808 32548 23860
rect 25228 23715 25280 23724
rect 25228 23681 25237 23715
rect 25237 23681 25271 23715
rect 25271 23681 25280 23715
rect 25228 23672 25280 23681
rect 24216 23604 24268 23656
rect 25044 23604 25096 23656
rect 25503 23715 25555 23724
rect 25503 23681 25534 23715
rect 25534 23681 25555 23715
rect 25503 23672 25555 23681
rect 29552 23715 29604 23724
rect 29552 23681 29561 23715
rect 29561 23681 29595 23715
rect 29595 23681 29604 23715
rect 29552 23672 29604 23681
rect 29736 23672 29788 23724
rect 25780 23604 25832 23656
rect 27160 23604 27212 23656
rect 31484 23672 31536 23724
rect 31668 23672 31720 23724
rect 32404 23715 32456 23724
rect 32404 23681 32413 23715
rect 32413 23681 32447 23715
rect 32447 23681 32456 23715
rect 32404 23672 32456 23681
rect 33692 23808 33744 23860
rect 33784 23808 33836 23860
rect 36728 23851 36780 23860
rect 32864 23740 32916 23792
rect 34428 23740 34480 23792
rect 36728 23817 36737 23851
rect 36737 23817 36771 23851
rect 36771 23817 36780 23851
rect 36728 23808 36780 23817
rect 32128 23604 32180 23656
rect 30472 23536 30524 23588
rect 21180 23511 21232 23520
rect 21180 23477 21189 23511
rect 21189 23477 21223 23511
rect 21223 23477 21232 23511
rect 21180 23468 21232 23477
rect 25688 23468 25740 23520
rect 27068 23468 27120 23520
rect 27160 23468 27212 23520
rect 27804 23468 27856 23520
rect 32220 23536 32272 23588
rect 32404 23468 32456 23520
rect 32588 23468 32640 23520
rect 32772 23468 32824 23520
rect 33416 23468 33468 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 5632 23307 5684 23316
rect 5632 23273 5641 23307
rect 5641 23273 5675 23307
rect 5675 23273 5684 23307
rect 5632 23264 5684 23273
rect 7472 23264 7524 23316
rect 12072 23264 12124 23316
rect 14556 23264 14608 23316
rect 16672 23264 16724 23316
rect 16856 23264 16908 23316
rect 17776 23264 17828 23316
rect 19156 23264 19208 23316
rect 19340 23307 19392 23316
rect 19340 23273 19349 23307
rect 19349 23273 19383 23307
rect 19383 23273 19392 23307
rect 21088 23307 21140 23316
rect 19340 23264 19392 23273
rect 21088 23273 21097 23307
rect 21097 23273 21131 23307
rect 21131 23273 21140 23307
rect 21088 23264 21140 23273
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 22928 23264 22980 23316
rect 25044 23264 25096 23316
rect 28908 23307 28960 23316
rect 6828 23196 6880 23248
rect 1584 23060 1636 23112
rect 3332 23128 3384 23180
rect 3792 23128 3844 23180
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 2964 23060 3016 23112
rect 5540 23060 5592 23112
rect 5724 23060 5776 23112
rect 7380 23128 7432 23180
rect 6920 23060 6972 23112
rect 7012 23103 7064 23112
rect 7012 23069 7021 23103
rect 7021 23069 7055 23103
rect 7055 23069 7064 23103
rect 7472 23103 7524 23112
rect 7012 23060 7064 23069
rect 7472 23069 7481 23103
rect 7481 23069 7515 23103
rect 7515 23069 7524 23103
rect 7472 23060 7524 23069
rect 7748 23196 7800 23248
rect 10140 23128 10192 23180
rect 2688 22992 2740 23044
rect 4620 22992 4672 23044
rect 2504 22924 2556 22976
rect 5448 22924 5500 22976
rect 7104 22992 7156 23044
rect 7840 23103 7892 23112
rect 7840 23069 7849 23103
rect 7849 23069 7883 23103
rect 7883 23069 7892 23103
rect 7840 23060 7892 23069
rect 8024 23060 8076 23112
rect 8852 23060 8904 23112
rect 9496 23060 9548 23112
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 10600 23060 10652 23069
rect 14464 23196 14516 23248
rect 12992 23171 13044 23180
rect 12992 23137 13001 23171
rect 13001 23137 13035 23171
rect 13035 23137 13044 23171
rect 12992 23128 13044 23137
rect 16120 23128 16172 23180
rect 15200 23103 15252 23112
rect 15200 23069 15218 23103
rect 15218 23069 15252 23103
rect 15200 23060 15252 23069
rect 16764 23060 16816 23112
rect 11520 22992 11572 23044
rect 8208 22924 8260 22976
rect 13268 22924 13320 22976
rect 13360 22924 13412 22976
rect 21180 23196 21232 23248
rect 23204 23196 23256 23248
rect 28908 23273 28917 23307
rect 28917 23273 28951 23307
rect 28951 23273 28960 23307
rect 28908 23264 28960 23273
rect 30288 23264 30340 23316
rect 33692 23307 33744 23316
rect 33692 23273 33701 23307
rect 33701 23273 33735 23307
rect 33735 23273 33744 23307
rect 33692 23264 33744 23273
rect 17500 23128 17552 23180
rect 17592 23060 17644 23112
rect 18236 23060 18288 23112
rect 20628 23060 20680 23112
rect 20904 23103 20956 23112
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 21272 23060 21324 23112
rect 25504 23128 25556 23180
rect 25780 23128 25832 23180
rect 26976 23171 27028 23180
rect 26976 23137 26985 23171
rect 26985 23137 27019 23171
rect 27019 23137 27028 23171
rect 26976 23128 27028 23137
rect 22100 23060 22152 23112
rect 23020 23060 23072 23112
rect 23296 23060 23348 23112
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 27068 23060 27120 23112
rect 33784 23196 33836 23248
rect 29552 23103 29604 23112
rect 29552 23069 29561 23103
rect 29561 23069 29595 23103
rect 29595 23069 29604 23103
rect 29552 23060 29604 23069
rect 31944 23128 31996 23180
rect 29920 23060 29972 23112
rect 32220 23103 32272 23112
rect 32220 23069 32229 23103
rect 32229 23069 32263 23103
rect 32263 23069 32272 23103
rect 32220 23060 32272 23069
rect 32404 23103 32456 23112
rect 32404 23069 32408 23103
rect 32408 23069 32442 23103
rect 32442 23069 32456 23103
rect 32404 23060 32456 23069
rect 32588 23103 32640 23112
rect 32588 23069 32597 23103
rect 32597 23069 32631 23103
rect 32631 23069 32640 23103
rect 32588 23060 32640 23069
rect 32772 23060 32824 23112
rect 18328 23035 18380 23044
rect 18328 23001 18337 23035
rect 18337 23001 18371 23035
rect 18371 23001 18380 23035
rect 18328 22992 18380 23001
rect 21180 22992 21232 23044
rect 21364 22992 21416 23044
rect 22008 22992 22060 23044
rect 23480 23035 23532 23044
rect 23480 23001 23489 23035
rect 23489 23001 23523 23035
rect 23523 23001 23532 23035
rect 23480 22992 23532 23001
rect 17684 22967 17736 22976
rect 17684 22933 17693 22967
rect 17693 22933 17727 22967
rect 17727 22933 17736 22967
rect 17684 22924 17736 22933
rect 22744 22967 22796 22976
rect 22744 22933 22753 22967
rect 22753 22933 22787 22967
rect 22787 22933 22796 22967
rect 22744 22924 22796 22933
rect 23664 22924 23716 22976
rect 24768 22924 24820 22976
rect 30656 22992 30708 23044
rect 32128 22992 32180 23044
rect 33416 22992 33468 23044
rect 30104 22924 30156 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 3976 22720 4028 22772
rect 4620 22720 4672 22772
rect 5448 22763 5500 22772
rect 5448 22729 5457 22763
rect 5457 22729 5491 22763
rect 5491 22729 5500 22763
rect 5448 22720 5500 22729
rect 13544 22763 13596 22772
rect 2136 22627 2188 22636
rect 2136 22593 2145 22627
rect 2145 22593 2179 22627
rect 2179 22593 2188 22627
rect 2136 22584 2188 22593
rect 3792 22652 3844 22704
rect 3240 22584 3292 22636
rect 6736 22584 6788 22636
rect 8208 22627 8260 22636
rect 8208 22593 8242 22627
rect 8242 22593 8260 22627
rect 8208 22584 8260 22593
rect 10600 22584 10652 22636
rect 11152 22584 11204 22636
rect 12164 22695 12216 22704
rect 12164 22661 12173 22695
rect 12173 22661 12207 22695
rect 12207 22661 12216 22695
rect 12164 22652 12216 22661
rect 13544 22729 13553 22763
rect 13553 22729 13587 22763
rect 13587 22729 13596 22763
rect 13544 22720 13596 22729
rect 17592 22720 17644 22772
rect 18144 22763 18196 22772
rect 18144 22729 18153 22763
rect 18153 22729 18187 22763
rect 18187 22729 18196 22763
rect 18144 22720 18196 22729
rect 18328 22720 18380 22772
rect 21272 22720 21324 22772
rect 29552 22720 29604 22772
rect 30472 22720 30524 22772
rect 32588 22720 32640 22772
rect 13176 22695 13228 22704
rect 5908 22516 5960 22568
rect 7104 22516 7156 22568
rect 7564 22516 7616 22568
rect 7748 22516 7800 22568
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 7932 22448 7984 22500
rect 9312 22491 9364 22500
rect 9312 22457 9321 22491
rect 9321 22457 9355 22491
rect 9355 22457 9364 22491
rect 12348 22627 12400 22636
rect 12348 22593 12362 22627
rect 12362 22593 12396 22627
rect 12396 22593 12400 22627
rect 12348 22584 12400 22593
rect 13176 22661 13185 22695
rect 13185 22661 13219 22695
rect 13219 22661 13228 22695
rect 13176 22652 13228 22661
rect 13360 22695 13412 22704
rect 13360 22661 13369 22695
rect 13369 22661 13403 22695
rect 13403 22661 13412 22695
rect 13360 22652 13412 22661
rect 13452 22652 13504 22704
rect 17684 22652 17736 22704
rect 22008 22695 22060 22704
rect 22008 22661 22017 22695
rect 22017 22661 22051 22695
rect 22051 22661 22060 22695
rect 22008 22652 22060 22661
rect 30104 22652 30156 22704
rect 15476 22584 15528 22636
rect 17408 22584 17460 22636
rect 20444 22584 20496 22636
rect 20812 22584 20864 22636
rect 24400 22627 24452 22636
rect 24400 22593 24410 22627
rect 24410 22593 24444 22627
rect 24444 22593 24452 22627
rect 24400 22584 24452 22593
rect 16304 22516 16356 22568
rect 22008 22516 22060 22568
rect 23204 22516 23256 22568
rect 9312 22448 9364 22457
rect 16396 22448 16448 22500
rect 22100 22448 22152 22500
rect 5172 22380 5224 22432
rect 8116 22380 8168 22432
rect 13268 22380 13320 22432
rect 15936 22380 15988 22432
rect 20628 22423 20680 22432
rect 20628 22389 20637 22423
rect 20637 22389 20671 22423
rect 20671 22389 20680 22423
rect 20628 22380 20680 22389
rect 23572 22448 23624 22500
rect 24952 22584 25004 22636
rect 31668 22584 31720 22636
rect 33508 22584 33560 22636
rect 37372 22584 37424 22636
rect 37556 22627 37608 22636
rect 37556 22593 37590 22627
rect 37590 22593 37608 22627
rect 37556 22584 37608 22593
rect 24676 22448 24728 22500
rect 67640 22491 67692 22500
rect 67640 22457 67649 22491
rect 67649 22457 67683 22491
rect 67683 22457 67692 22491
rect 67640 22448 67692 22457
rect 23480 22380 23532 22432
rect 24860 22380 24912 22432
rect 31116 22380 31168 22432
rect 32036 22380 32088 22432
rect 32956 22423 33008 22432
rect 32956 22389 32965 22423
rect 32965 22389 32999 22423
rect 32999 22389 33008 22423
rect 32956 22380 33008 22389
rect 38660 22423 38712 22432
rect 38660 22389 38669 22423
rect 38669 22389 38703 22423
rect 38703 22389 38712 22423
rect 38660 22380 38712 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 2320 22176 2372 22228
rect 3792 22108 3844 22160
rect 6736 22176 6788 22228
rect 9496 22151 9548 22160
rect 4620 22040 4672 22092
rect 9496 22117 9505 22151
rect 9505 22117 9539 22151
rect 9539 22117 9548 22151
rect 9496 22108 9548 22117
rect 10968 22108 11020 22160
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 2136 21972 2188 22024
rect 1768 21947 1820 21956
rect 1768 21913 1777 21947
rect 1777 21913 1811 21947
rect 1811 21913 1820 21947
rect 1768 21904 1820 21913
rect 5632 21972 5684 22024
rect 9312 22040 9364 22092
rect 12072 22108 12124 22160
rect 12256 22151 12308 22160
rect 12256 22117 12265 22151
rect 12265 22117 12299 22151
rect 12299 22117 12308 22151
rect 12256 22108 12308 22117
rect 17592 22176 17644 22228
rect 12532 22108 12584 22160
rect 14188 22108 14240 22160
rect 19432 22176 19484 22228
rect 20628 22176 20680 22228
rect 23572 22176 23624 22228
rect 27344 22176 27396 22228
rect 27620 22219 27672 22228
rect 27620 22185 27629 22219
rect 27629 22185 27663 22219
rect 27663 22185 27672 22219
rect 27620 22176 27672 22185
rect 1676 21836 1728 21888
rect 2780 21836 2832 21888
rect 3056 21879 3108 21888
rect 3056 21845 3065 21879
rect 3065 21845 3099 21879
rect 3099 21845 3108 21879
rect 3056 21836 3108 21845
rect 4620 21904 4672 21956
rect 7196 21947 7248 21956
rect 3332 21836 3384 21888
rect 6552 21836 6604 21888
rect 7196 21913 7205 21947
rect 7205 21913 7239 21947
rect 7239 21913 7248 21947
rect 7196 21904 7248 21913
rect 7932 21972 7984 22024
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 11704 22015 11756 22024
rect 11704 21981 11714 22015
rect 11714 21981 11748 22015
rect 11748 21981 11756 22015
rect 15476 22040 15528 22092
rect 11704 21972 11756 21981
rect 12348 21972 12400 22024
rect 13452 21972 13504 22024
rect 14648 22015 14700 22024
rect 8852 21904 8904 21956
rect 11980 21947 12032 21956
rect 11980 21913 11989 21947
rect 11989 21913 12023 21947
rect 12023 21913 12032 21947
rect 14648 21981 14657 22015
rect 14657 21981 14691 22015
rect 14691 21981 14700 22015
rect 14648 21972 14700 21981
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 16028 22015 16080 22024
rect 16028 21981 16038 22015
rect 16038 21981 16072 22015
rect 16072 21981 16080 22015
rect 20536 22108 20588 22160
rect 20996 22108 21048 22160
rect 20720 22040 20772 22092
rect 22008 22040 22060 22092
rect 22192 22040 22244 22092
rect 16028 21972 16080 21981
rect 11980 21904 12032 21913
rect 14372 21904 14424 21956
rect 15016 21904 15068 21956
rect 15476 21904 15528 21956
rect 13452 21836 13504 21888
rect 15752 21836 15804 21888
rect 18788 21904 18840 21956
rect 18512 21836 18564 21888
rect 19432 21904 19484 21956
rect 20536 21947 20588 21956
rect 20536 21913 20545 21947
rect 20545 21913 20579 21947
rect 20579 21913 20588 21947
rect 20536 21904 20588 21913
rect 20904 21972 20956 22024
rect 21824 21972 21876 22024
rect 22100 22015 22152 22024
rect 22100 21981 22109 22015
rect 22109 21981 22143 22015
rect 22143 21981 22152 22015
rect 22100 21972 22152 21981
rect 22284 22015 22336 22024
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 23388 22108 23440 22160
rect 22468 22015 22520 22024
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 22468 21972 22520 21981
rect 22652 21972 22704 22024
rect 22836 22040 22888 22092
rect 23388 22015 23440 22024
rect 23388 21981 23397 22015
rect 23397 21981 23431 22015
rect 23431 21981 23440 22015
rect 23388 21972 23440 21981
rect 24584 22015 24636 22024
rect 24584 21981 24591 22015
rect 24591 21981 24636 22015
rect 20720 21836 20772 21888
rect 21272 21836 21324 21888
rect 22192 21904 22244 21956
rect 22560 21904 22612 21956
rect 24584 21972 24636 21981
rect 24676 21947 24728 21956
rect 24676 21913 24685 21947
rect 24685 21913 24719 21947
rect 24719 21913 24728 21947
rect 24676 21904 24728 21913
rect 24952 21972 25004 22024
rect 25688 21972 25740 22024
rect 28172 22015 28224 22024
rect 28172 21981 28181 22015
rect 28181 21981 28215 22015
rect 28215 21981 28224 22015
rect 28172 21972 28224 21981
rect 28264 21972 28316 22024
rect 28448 22015 28500 22024
rect 28448 21981 28457 22015
rect 28457 21981 28491 22015
rect 28491 21981 28500 22015
rect 28448 21972 28500 21981
rect 31392 22040 31444 22092
rect 27620 21904 27672 21956
rect 30104 21972 30156 22024
rect 31760 21972 31812 22024
rect 32404 22040 32456 22092
rect 32036 22015 32088 22024
rect 32036 21981 32045 22015
rect 32045 21981 32079 22015
rect 32079 21981 32088 22015
rect 32036 21972 32088 21981
rect 31208 21904 31260 21956
rect 32220 22015 32272 22024
rect 32220 21981 32229 22015
rect 32229 21981 32263 22015
rect 32263 21981 32272 22015
rect 32220 21972 32272 21981
rect 33140 22015 33192 22024
rect 33140 21981 33149 22015
rect 33149 21981 33183 22015
rect 33183 21981 33192 22015
rect 33140 21972 33192 21981
rect 33324 22015 33376 22024
rect 33324 21981 33333 22015
rect 33333 21981 33367 22015
rect 33367 21981 33376 22015
rect 33324 21972 33376 21981
rect 34336 21972 34388 22024
rect 34520 21972 34572 22024
rect 37464 21972 37516 22024
rect 23388 21836 23440 21888
rect 25228 21836 25280 21888
rect 26976 21879 27028 21888
rect 26976 21845 26985 21879
rect 26985 21845 27019 21879
rect 27019 21845 27028 21879
rect 26976 21836 27028 21845
rect 27436 21836 27488 21888
rect 31392 21836 31444 21888
rect 32404 21836 32456 21888
rect 33968 21836 34020 21888
rect 34888 21879 34940 21888
rect 34888 21845 34897 21879
rect 34897 21845 34931 21879
rect 34931 21845 34940 21879
rect 34888 21836 34940 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 3240 21632 3292 21684
rect 1584 21539 1636 21548
rect 1584 21505 1593 21539
rect 1593 21505 1627 21539
rect 1627 21505 1636 21539
rect 1584 21496 1636 21505
rect 1676 21496 1728 21548
rect 5448 21564 5500 21616
rect 9404 21632 9456 21684
rect 10232 21632 10284 21684
rect 10600 21675 10652 21684
rect 10600 21641 10609 21675
rect 10609 21641 10643 21675
rect 10643 21641 10652 21675
rect 10600 21632 10652 21641
rect 15200 21632 15252 21684
rect 9496 21607 9548 21616
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 7840 21496 7892 21548
rect 9496 21573 9530 21607
rect 9530 21573 9548 21607
rect 9496 21564 9548 21573
rect 9588 21564 9640 21616
rect 11520 21496 11572 21548
rect 2780 21428 2832 21480
rect 2320 21360 2372 21412
rect 9220 21471 9272 21480
rect 9220 21437 9229 21471
rect 9229 21437 9263 21471
rect 9263 21437 9272 21471
rect 9220 21428 9272 21437
rect 4804 21360 4856 21412
rect 13084 21564 13136 21616
rect 15476 21607 15528 21616
rect 15476 21573 15485 21607
rect 15485 21573 15519 21607
rect 15519 21573 15528 21607
rect 15476 21564 15528 21573
rect 16580 21564 16632 21616
rect 28264 21675 28316 21684
rect 22284 21564 22336 21616
rect 24676 21564 24728 21616
rect 13268 21496 13320 21548
rect 13544 21539 13596 21548
rect 13544 21505 13553 21539
rect 13553 21505 13587 21539
rect 13587 21505 13596 21539
rect 13544 21496 13596 21505
rect 15200 21539 15252 21548
rect 15200 21505 15209 21539
rect 15209 21505 15243 21539
rect 15243 21505 15252 21539
rect 15200 21496 15252 21505
rect 15384 21539 15436 21548
rect 15384 21505 15391 21539
rect 15391 21505 15436 21539
rect 15384 21496 15436 21505
rect 2688 21292 2740 21344
rect 5908 21292 5960 21344
rect 9220 21292 9272 21344
rect 9588 21292 9640 21344
rect 12532 21292 12584 21344
rect 13268 21292 13320 21344
rect 13452 21360 13504 21412
rect 14464 21428 14516 21480
rect 15752 21496 15804 21548
rect 15844 21496 15896 21548
rect 18880 21496 18932 21548
rect 19432 21496 19484 21548
rect 20076 21496 20128 21548
rect 20536 21539 20588 21548
rect 18052 21471 18104 21480
rect 13728 21292 13780 21344
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 20536 21505 20545 21539
rect 20545 21505 20579 21539
rect 20579 21505 20588 21539
rect 20536 21496 20588 21505
rect 20904 21496 20956 21548
rect 22928 21539 22980 21548
rect 22928 21505 22937 21539
rect 22937 21505 22971 21539
rect 22971 21505 22980 21539
rect 22928 21496 22980 21505
rect 23848 21496 23900 21548
rect 24952 21496 25004 21548
rect 22468 21360 22520 21412
rect 22652 21471 22704 21480
rect 22652 21437 22661 21471
rect 22661 21437 22695 21471
rect 22695 21437 22704 21471
rect 25412 21539 25464 21548
rect 25412 21505 25421 21539
rect 25421 21505 25455 21539
rect 25455 21505 25464 21539
rect 25596 21539 25648 21548
rect 25412 21496 25464 21505
rect 25596 21505 25604 21539
rect 25604 21505 25638 21539
rect 25638 21505 25648 21539
rect 25596 21496 25648 21505
rect 28264 21641 28273 21675
rect 28273 21641 28307 21675
rect 28307 21641 28316 21675
rect 28264 21632 28316 21641
rect 30656 21675 30708 21684
rect 30656 21641 30665 21675
rect 30665 21641 30699 21675
rect 30699 21641 30708 21675
rect 30656 21632 30708 21641
rect 27436 21564 27488 21616
rect 27988 21496 28040 21548
rect 29276 21496 29328 21548
rect 32588 21632 32640 21684
rect 33140 21632 33192 21684
rect 33508 21675 33560 21684
rect 33508 21641 33517 21675
rect 33517 21641 33551 21675
rect 33551 21641 33560 21675
rect 33508 21632 33560 21641
rect 31208 21564 31260 21616
rect 31668 21564 31720 21616
rect 34888 21632 34940 21684
rect 37556 21632 37608 21684
rect 31116 21539 31168 21548
rect 31116 21505 31125 21539
rect 31125 21505 31159 21539
rect 31159 21505 31168 21539
rect 31116 21496 31168 21505
rect 31392 21496 31444 21548
rect 33968 21564 34020 21616
rect 34336 21496 34388 21548
rect 35992 21539 36044 21548
rect 35992 21505 36001 21539
rect 36001 21505 36035 21539
rect 36035 21505 36044 21539
rect 35992 21496 36044 21505
rect 36176 21539 36228 21548
rect 36176 21505 36185 21539
rect 36185 21505 36219 21539
rect 36219 21505 36228 21539
rect 36176 21496 36228 21505
rect 36268 21539 36320 21548
rect 36268 21505 36280 21539
rect 36280 21505 36314 21539
rect 36314 21505 36320 21539
rect 36268 21496 36320 21505
rect 39304 21564 39356 21616
rect 37464 21539 37516 21548
rect 37464 21505 37473 21539
rect 37473 21505 37507 21539
rect 37507 21505 37516 21539
rect 37464 21496 37516 21505
rect 37740 21539 37792 21548
rect 37740 21505 37774 21539
rect 37774 21505 37792 21539
rect 37740 21496 37792 21505
rect 22652 21428 22704 21437
rect 23112 21360 23164 21412
rect 25504 21360 25556 21412
rect 15384 21292 15436 21344
rect 16580 21292 16632 21344
rect 20812 21292 20864 21344
rect 25044 21335 25096 21344
rect 25044 21301 25053 21335
rect 25053 21301 25087 21335
rect 25087 21301 25096 21335
rect 25044 21292 25096 21301
rect 32956 21360 33008 21412
rect 34520 21292 34572 21344
rect 38844 21335 38896 21344
rect 38844 21301 38853 21335
rect 38853 21301 38887 21335
rect 38887 21301 38896 21335
rect 38844 21292 38896 21301
rect 67640 21335 67692 21344
rect 67640 21301 67649 21335
rect 67649 21301 67683 21335
rect 67683 21301 67692 21335
rect 67640 21292 67692 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 13452 21088 13504 21140
rect 14464 21088 14516 21140
rect 15568 21088 15620 21140
rect 15844 21131 15896 21140
rect 15844 21097 15853 21131
rect 15853 21097 15887 21131
rect 15887 21097 15896 21131
rect 15844 21088 15896 21097
rect 16212 21088 16264 21140
rect 18512 21088 18564 21140
rect 19432 21088 19484 21140
rect 20904 21088 20956 21140
rect 22468 21088 22520 21140
rect 34060 21131 34112 21140
rect 34060 21097 34069 21131
rect 34069 21097 34103 21131
rect 34103 21097 34112 21131
rect 34060 21088 34112 21097
rect 36176 21088 36228 21140
rect 37740 21088 37792 21140
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 2504 20884 2556 20936
rect 3884 20884 3936 20936
rect 9312 20927 9364 20936
rect 1768 20816 1820 20868
rect 2228 20791 2280 20800
rect 2228 20757 2237 20791
rect 2237 20757 2271 20791
rect 2271 20757 2280 20791
rect 2228 20748 2280 20757
rect 3424 20816 3476 20868
rect 7748 20816 7800 20868
rect 7840 20816 7892 20868
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 3056 20748 3108 20800
rect 5724 20748 5776 20800
rect 8208 20748 8260 20800
rect 9680 20816 9732 20868
rect 14188 21020 14240 21072
rect 15292 21020 15344 21072
rect 10692 20952 10744 21004
rect 10508 20884 10560 20936
rect 12900 20952 12952 21004
rect 11520 20884 11572 20936
rect 12164 20927 12216 20936
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 12992 20927 13044 20936
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 13452 20884 13504 20936
rect 15200 20927 15252 20936
rect 15200 20893 15209 20927
rect 15209 20893 15243 20927
rect 15243 20893 15252 20927
rect 15200 20884 15252 20893
rect 15384 20927 15436 20936
rect 15384 20893 15393 20927
rect 15393 20893 15427 20927
rect 15427 20893 15436 20927
rect 15384 20884 15436 20893
rect 20536 21020 20588 21072
rect 25136 21020 25188 21072
rect 26332 21063 26384 21072
rect 26332 21029 26341 21063
rect 26341 21029 26375 21063
rect 26375 21029 26384 21063
rect 26332 21020 26384 21029
rect 30656 21020 30708 21072
rect 31208 21020 31260 21072
rect 13176 20859 13228 20868
rect 13176 20825 13185 20859
rect 13185 20825 13219 20859
rect 13219 20825 13228 20859
rect 13176 20816 13228 20825
rect 13820 20816 13872 20868
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 18236 20884 18288 20936
rect 18880 20884 18932 20936
rect 16856 20816 16908 20868
rect 17960 20816 18012 20868
rect 20168 20884 20220 20936
rect 23664 20884 23716 20936
rect 25412 20927 25464 20936
rect 25412 20893 25421 20927
rect 25421 20893 25455 20927
rect 25455 20893 25464 20927
rect 25412 20884 25464 20893
rect 30288 20952 30340 21004
rect 31392 20952 31444 21004
rect 11704 20791 11756 20800
rect 11704 20757 11713 20791
rect 11713 20757 11747 20791
rect 11747 20757 11756 20791
rect 11704 20748 11756 20757
rect 13912 20748 13964 20800
rect 18512 20748 18564 20800
rect 19984 20816 20036 20868
rect 20720 20748 20772 20800
rect 21824 20791 21876 20800
rect 21824 20757 21833 20791
rect 21833 20757 21867 20791
rect 21867 20757 21876 20791
rect 21824 20748 21876 20757
rect 22192 20816 22244 20868
rect 23388 20816 23440 20868
rect 27620 20884 27672 20936
rect 31116 20884 31168 20936
rect 31668 20884 31720 20936
rect 34428 20952 34480 21004
rect 28448 20816 28500 20868
rect 31944 20859 31996 20868
rect 22376 20748 22428 20800
rect 29276 20748 29328 20800
rect 30288 20748 30340 20800
rect 31944 20825 31953 20859
rect 31953 20825 31987 20859
rect 31987 20825 31996 20859
rect 31944 20816 31996 20825
rect 32956 20927 33008 20936
rect 32956 20893 32965 20927
rect 32965 20893 32999 20927
rect 32999 20893 33008 20927
rect 32956 20884 33008 20893
rect 34612 20884 34664 20936
rect 35992 20884 36044 20936
rect 37188 20927 37240 20936
rect 37188 20893 37197 20927
rect 37197 20893 37231 20927
rect 37231 20893 37240 20927
rect 37188 20884 37240 20893
rect 37372 20927 37424 20936
rect 37372 20893 37381 20927
rect 37381 20893 37415 20927
rect 37415 20893 37424 20927
rect 37372 20884 37424 20893
rect 32220 20748 32272 20800
rect 33232 20791 33284 20800
rect 33232 20757 33241 20791
rect 33241 20757 33275 20791
rect 33275 20757 33284 20791
rect 33232 20748 33284 20757
rect 36084 20748 36136 20800
rect 36268 20816 36320 20868
rect 37556 20927 37608 20936
rect 37556 20893 37565 20927
rect 37565 20893 37599 20927
rect 37599 20893 37608 20927
rect 37556 20884 37608 20893
rect 37648 20816 37700 20868
rect 38660 20748 38712 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 3424 20544 3476 20596
rect 4620 20544 4672 20596
rect 7748 20587 7800 20596
rect 7748 20553 7757 20587
rect 7757 20553 7791 20587
rect 7791 20553 7800 20587
rect 7748 20544 7800 20553
rect 7932 20544 7984 20596
rect 8944 20544 8996 20596
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 16856 20544 16908 20596
rect 19984 20587 20036 20596
rect 19984 20553 19993 20587
rect 19993 20553 20027 20587
rect 20027 20553 20036 20587
rect 19984 20544 20036 20553
rect 20444 20544 20496 20596
rect 22008 20544 22060 20596
rect 24308 20544 24360 20596
rect 25412 20544 25464 20596
rect 1584 20408 1636 20460
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 2320 20451 2372 20460
rect 2320 20417 2329 20451
rect 2329 20417 2363 20451
rect 2363 20417 2372 20451
rect 2320 20408 2372 20417
rect 2136 20340 2188 20392
rect 4804 20476 4856 20528
rect 7196 20519 7248 20528
rect 7196 20485 7205 20519
rect 7205 20485 7239 20519
rect 7239 20485 7248 20519
rect 7196 20476 7248 20485
rect 9220 20476 9272 20528
rect 9404 20476 9456 20528
rect 11704 20476 11756 20528
rect 3424 20451 3476 20460
rect 3424 20417 3433 20451
rect 3433 20417 3467 20451
rect 3467 20417 3476 20451
rect 3424 20408 3476 20417
rect 6552 20408 6604 20460
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 5816 20272 5868 20324
rect 7932 20408 7984 20460
rect 8116 20451 8168 20460
rect 8116 20417 8125 20451
rect 8125 20417 8159 20451
rect 8159 20417 8168 20451
rect 8116 20408 8168 20417
rect 8208 20451 8260 20460
rect 8208 20417 8217 20451
rect 8217 20417 8251 20451
rect 8251 20417 8260 20451
rect 8208 20408 8260 20417
rect 15568 20408 15620 20460
rect 18052 20476 18104 20528
rect 20720 20476 20772 20528
rect 22744 20519 22796 20528
rect 22744 20485 22778 20519
rect 22778 20485 22796 20519
rect 22744 20476 22796 20485
rect 31944 20544 31996 20596
rect 17960 20451 18012 20460
rect 17960 20417 17994 20451
rect 17994 20417 18012 20451
rect 10508 20340 10560 20392
rect 11980 20272 12032 20324
rect 5080 20204 5132 20256
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 5724 20204 5776 20213
rect 6460 20204 6512 20256
rect 6736 20204 6788 20256
rect 9496 20247 9548 20256
rect 9496 20213 9505 20247
rect 9505 20213 9539 20247
rect 9539 20213 9548 20247
rect 9496 20204 9548 20213
rect 11520 20247 11572 20256
rect 11520 20213 11529 20247
rect 11529 20213 11563 20247
rect 11563 20213 11572 20247
rect 11520 20204 11572 20213
rect 13176 20204 13228 20256
rect 15752 20204 15804 20256
rect 17960 20408 18012 20417
rect 20812 20408 20864 20460
rect 21824 20408 21876 20460
rect 24952 20408 25004 20460
rect 25320 20451 25372 20460
rect 25320 20417 25329 20451
rect 25329 20417 25363 20451
rect 25363 20417 25372 20451
rect 25320 20408 25372 20417
rect 21088 20340 21140 20392
rect 22468 20272 22520 20324
rect 25596 20451 25648 20460
rect 25596 20417 25605 20451
rect 25605 20417 25639 20451
rect 25639 20417 25648 20451
rect 25596 20408 25648 20417
rect 31392 20476 31444 20528
rect 26516 20408 26568 20460
rect 27988 20451 28040 20460
rect 27988 20417 27997 20451
rect 27997 20417 28031 20451
rect 28031 20417 28040 20451
rect 27988 20408 28040 20417
rect 26332 20340 26384 20392
rect 26424 20272 26476 20324
rect 29000 20408 29052 20460
rect 31760 20408 31812 20460
rect 32404 20408 32456 20460
rect 33232 20408 33284 20460
rect 34520 20451 34572 20460
rect 34520 20417 34529 20451
rect 34529 20417 34563 20451
rect 34563 20417 34572 20451
rect 34520 20408 34572 20417
rect 34704 20408 34756 20460
rect 23388 20204 23440 20256
rect 23848 20247 23900 20256
rect 23848 20213 23857 20247
rect 23857 20213 23891 20247
rect 23891 20213 23900 20247
rect 23848 20204 23900 20213
rect 26056 20204 26108 20256
rect 28540 20204 28592 20256
rect 31944 20204 31996 20256
rect 32956 20204 33008 20256
rect 37556 20204 37608 20256
rect 40408 20204 40460 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 9404 20000 9456 20052
rect 9588 20000 9640 20052
rect 2320 19932 2372 19984
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 2044 19796 2096 19848
rect 2504 19839 2556 19848
rect 2504 19805 2513 19839
rect 2513 19805 2547 19839
rect 2547 19805 2556 19839
rect 2504 19796 2556 19805
rect 2412 19728 2464 19780
rect 5448 19796 5500 19848
rect 6460 19839 6512 19848
rect 6460 19805 6469 19839
rect 6469 19805 6503 19839
rect 6503 19805 6512 19839
rect 6460 19796 6512 19805
rect 7104 19932 7156 19984
rect 10048 19932 10100 19984
rect 10692 19932 10744 19984
rect 6736 19796 6788 19848
rect 7472 19864 7524 19916
rect 8116 19864 8168 19916
rect 12716 20000 12768 20052
rect 13728 20000 13780 20052
rect 21088 20000 21140 20052
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 24124 20000 24176 20052
rect 13820 19932 13872 19984
rect 5264 19728 5316 19780
rect 9128 19796 9180 19848
rect 7472 19728 7524 19780
rect 2688 19660 2740 19712
rect 2964 19703 3016 19712
rect 2964 19669 2973 19703
rect 2973 19669 3007 19703
rect 3007 19669 3016 19703
rect 2964 19660 3016 19669
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 6184 19703 6236 19712
rect 6184 19669 6193 19703
rect 6193 19669 6227 19703
rect 6227 19669 6236 19703
rect 6184 19660 6236 19669
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 10508 19839 10560 19848
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 10692 19839 10744 19848
rect 10692 19805 10701 19839
rect 10701 19805 10735 19839
rect 10735 19805 10744 19839
rect 10692 19796 10744 19805
rect 10968 19796 11020 19848
rect 14740 19796 14792 19848
rect 17776 19932 17828 19984
rect 15752 19907 15804 19916
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 20720 19864 20772 19916
rect 13728 19728 13780 19780
rect 15016 19839 15068 19848
rect 15016 19805 15025 19839
rect 15025 19805 15059 19839
rect 15059 19805 15068 19839
rect 15016 19796 15068 19805
rect 17316 19796 17368 19848
rect 22468 19932 22520 19984
rect 22100 19839 22152 19848
rect 13820 19660 13872 19712
rect 15200 19728 15252 19780
rect 16856 19728 16908 19780
rect 15016 19660 15068 19712
rect 15476 19660 15528 19712
rect 22100 19805 22109 19839
rect 22109 19805 22143 19839
rect 22143 19805 22152 19839
rect 22100 19796 22152 19805
rect 23296 19839 23348 19848
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 23296 19796 23348 19805
rect 24124 19796 24176 19848
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 25596 20000 25648 20052
rect 27804 20043 27856 20052
rect 27804 20009 27813 20043
rect 27813 20009 27847 20043
rect 27847 20009 27856 20043
rect 27804 20000 27856 20009
rect 29000 20043 29052 20052
rect 29000 20009 29009 20043
rect 29009 20009 29043 20043
rect 29043 20009 29052 20043
rect 29000 20000 29052 20009
rect 32220 20000 32272 20052
rect 25688 19864 25740 19916
rect 20628 19728 20680 19780
rect 23940 19728 23992 19780
rect 20260 19660 20312 19712
rect 20996 19660 21048 19712
rect 22192 19660 22244 19712
rect 25964 19839 26016 19848
rect 25964 19805 25974 19839
rect 25974 19805 26008 19839
rect 26008 19805 26016 19839
rect 28448 19864 28500 19916
rect 25964 19796 26016 19805
rect 28172 19796 28224 19848
rect 28540 19839 28592 19848
rect 28540 19805 28549 19839
rect 28549 19805 28583 19839
rect 28583 19805 28592 19839
rect 28540 19796 28592 19805
rect 34704 20000 34756 20052
rect 37372 20000 37424 20052
rect 35532 19975 35584 19984
rect 35532 19941 35541 19975
rect 35541 19941 35575 19975
rect 35575 19941 35584 19975
rect 35532 19932 35584 19941
rect 37464 19864 37516 19916
rect 26148 19771 26200 19780
rect 26148 19737 26157 19771
rect 26157 19737 26191 19771
rect 26191 19737 26200 19771
rect 26148 19728 26200 19737
rect 32404 19796 32456 19848
rect 36084 19839 36136 19848
rect 36084 19805 36093 19839
rect 36093 19805 36127 19839
rect 36127 19805 36136 19839
rect 36084 19796 36136 19805
rect 37096 19796 37148 19848
rect 37372 19796 37424 19848
rect 68100 19839 68152 19848
rect 31116 19728 31168 19780
rect 31208 19728 31260 19780
rect 36176 19728 36228 19780
rect 38108 19728 38160 19780
rect 26516 19703 26568 19712
rect 26516 19669 26525 19703
rect 26525 19669 26559 19703
rect 26559 19669 26568 19703
rect 26516 19660 26568 19669
rect 30748 19660 30800 19712
rect 36544 19660 36596 19712
rect 37188 19660 37240 19712
rect 38844 19660 38896 19712
rect 68100 19805 68109 19839
rect 68109 19805 68143 19839
rect 68143 19805 68152 19839
rect 68100 19796 68152 19805
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 2504 19456 2556 19508
rect 2596 19499 2648 19508
rect 2596 19465 2605 19499
rect 2605 19465 2639 19499
rect 2639 19465 2648 19499
rect 5816 19499 5868 19508
rect 2596 19456 2648 19465
rect 5816 19465 5825 19499
rect 5825 19465 5859 19499
rect 5859 19465 5868 19499
rect 5816 19456 5868 19465
rect 1768 19431 1820 19440
rect 1768 19397 1777 19431
rect 1777 19397 1811 19431
rect 1811 19397 1820 19431
rect 1768 19388 1820 19397
rect 2964 19388 3016 19440
rect 6184 19388 6236 19440
rect 6644 19388 6696 19440
rect 3884 19320 3936 19372
rect 5080 19320 5132 19372
rect 11060 19456 11112 19508
rect 11520 19456 11572 19508
rect 11796 19456 11848 19508
rect 9588 19388 9640 19440
rect 10140 19388 10192 19440
rect 6920 19252 6972 19304
rect 10416 19320 10468 19372
rect 12716 19456 12768 19508
rect 13452 19456 13504 19508
rect 15384 19456 15436 19508
rect 15936 19456 15988 19508
rect 14740 19388 14792 19440
rect 15292 19388 15344 19440
rect 15568 19431 15620 19440
rect 15568 19397 15577 19431
rect 15577 19397 15611 19431
rect 15611 19397 15620 19431
rect 15568 19388 15620 19397
rect 13452 19320 13504 19372
rect 13912 19363 13964 19372
rect 13912 19329 13921 19363
rect 13921 19329 13955 19363
rect 13955 19329 13964 19363
rect 13912 19320 13964 19329
rect 14004 19363 14056 19372
rect 14004 19329 14014 19363
rect 14014 19329 14048 19363
rect 14048 19329 14056 19363
rect 14004 19320 14056 19329
rect 10692 19252 10744 19304
rect 14372 19363 14424 19372
rect 14372 19329 14386 19363
rect 14386 19329 14420 19363
rect 14420 19329 14424 19363
rect 14372 19320 14424 19329
rect 15476 19320 15528 19372
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 17408 19320 17460 19372
rect 20260 19320 20312 19372
rect 20904 19363 20956 19372
rect 20904 19329 20913 19363
rect 20913 19329 20947 19363
rect 20947 19329 20956 19363
rect 20904 19320 20956 19329
rect 14648 19252 14700 19304
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 16856 19295 16908 19304
rect 16856 19261 16865 19295
rect 16865 19261 16899 19295
rect 16899 19261 16908 19295
rect 16856 19252 16908 19261
rect 20996 19329 21002 19346
rect 21002 19329 21036 19346
rect 21036 19329 21048 19346
rect 20996 19294 21048 19329
rect 12808 19227 12860 19236
rect 5356 19116 5408 19168
rect 6460 19116 6512 19168
rect 10140 19116 10192 19168
rect 12808 19193 12817 19227
rect 12817 19193 12851 19227
rect 12851 19193 12860 19227
rect 12808 19184 12860 19193
rect 14004 19184 14056 19236
rect 14188 19184 14240 19236
rect 20628 19227 20680 19236
rect 20628 19193 20637 19227
rect 20637 19193 20671 19227
rect 20671 19193 20680 19227
rect 20628 19184 20680 19193
rect 14464 19116 14516 19168
rect 16672 19116 16724 19168
rect 20076 19116 20128 19168
rect 22008 19320 22060 19372
rect 22189 19363 22241 19372
rect 22189 19329 22198 19363
rect 22198 19329 22232 19363
rect 22232 19329 22241 19363
rect 22189 19320 22241 19329
rect 23940 19388 23992 19440
rect 25596 19456 25648 19508
rect 31208 19499 31260 19508
rect 31208 19465 31217 19499
rect 31217 19465 31251 19499
rect 31251 19465 31260 19499
rect 31208 19456 31260 19465
rect 37280 19456 37332 19508
rect 38108 19499 38160 19508
rect 38108 19465 38117 19499
rect 38117 19465 38151 19499
rect 38151 19465 38160 19499
rect 38108 19456 38160 19465
rect 22560 19294 22612 19346
rect 22928 19252 22980 19304
rect 21456 19116 21508 19168
rect 22652 19184 22704 19236
rect 24032 19363 24084 19372
rect 24032 19329 24041 19363
rect 24041 19329 24075 19363
rect 24075 19329 24084 19363
rect 24032 19320 24084 19329
rect 24124 19320 24176 19372
rect 25688 19320 25740 19372
rect 26148 19363 26200 19372
rect 26148 19329 26157 19363
rect 26157 19329 26191 19363
rect 26191 19329 26200 19363
rect 26332 19363 26384 19372
rect 26148 19320 26200 19329
rect 26332 19329 26340 19363
rect 26340 19329 26374 19363
rect 26374 19329 26384 19363
rect 26332 19320 26384 19329
rect 30656 19388 30708 19440
rect 26700 19320 26752 19372
rect 28816 19320 28868 19372
rect 29828 19320 29880 19372
rect 30104 19320 30156 19372
rect 30748 19363 30800 19372
rect 30748 19329 30757 19363
rect 30757 19329 30791 19363
rect 30791 19329 30800 19363
rect 30748 19320 30800 19329
rect 34520 19388 34572 19440
rect 26884 19252 26936 19304
rect 34888 19320 34940 19372
rect 35532 19388 35584 19440
rect 22100 19116 22152 19168
rect 22560 19116 22612 19168
rect 24860 19116 24912 19168
rect 26608 19116 26660 19168
rect 36544 19363 36596 19372
rect 36544 19329 36553 19363
rect 36553 19329 36587 19363
rect 36587 19329 36596 19363
rect 36544 19320 36596 19329
rect 37096 19320 37148 19372
rect 37372 19320 37424 19372
rect 37556 19320 37608 19372
rect 38476 19363 38528 19372
rect 38476 19329 38485 19363
rect 38485 19329 38519 19363
rect 38519 19329 38528 19363
rect 38476 19320 38528 19329
rect 38844 19320 38896 19372
rect 30288 19116 30340 19168
rect 33968 19116 34020 19168
rect 36268 19184 36320 19236
rect 36452 19184 36504 19236
rect 37556 19116 37608 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 6920 18912 6972 18964
rect 8944 18955 8996 18964
rect 8944 18921 8953 18955
rect 8953 18921 8987 18955
rect 8987 18921 8996 18955
rect 8944 18912 8996 18921
rect 11336 18912 11388 18964
rect 17316 18912 17368 18964
rect 18696 18955 18748 18964
rect 18696 18921 18705 18955
rect 18705 18921 18739 18955
rect 18739 18921 18748 18955
rect 18696 18912 18748 18921
rect 20536 18912 20588 18964
rect 2044 18776 2096 18828
rect 3148 18776 3200 18828
rect 7564 18844 7616 18896
rect 10508 18844 10560 18896
rect 11704 18844 11756 18896
rect 15844 18844 15896 18896
rect 24860 18912 24912 18964
rect 6552 18640 6604 18692
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 13912 18776 13964 18828
rect 15568 18776 15620 18828
rect 20720 18776 20772 18828
rect 9680 18640 9732 18692
rect 10048 18640 10100 18692
rect 3148 18615 3200 18624
rect 3148 18581 3157 18615
rect 3157 18581 3191 18615
rect 3191 18581 3200 18615
rect 3148 18572 3200 18581
rect 3792 18572 3844 18624
rect 4896 18572 4948 18624
rect 5264 18572 5316 18624
rect 12440 18708 12492 18760
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 12624 18708 12676 18717
rect 13360 18708 13412 18760
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 18512 18708 18564 18760
rect 18696 18708 18748 18760
rect 20076 18708 20128 18760
rect 21456 18708 21508 18760
rect 21732 18708 21784 18760
rect 21916 18708 21968 18760
rect 22560 18708 22612 18760
rect 23940 18708 23992 18760
rect 29828 18912 29880 18964
rect 34796 18912 34848 18964
rect 35072 18912 35124 18964
rect 36268 18912 36320 18964
rect 37648 18912 37700 18964
rect 38476 18912 38528 18964
rect 27436 18776 27488 18828
rect 30656 18844 30708 18896
rect 31116 18844 31168 18896
rect 30380 18776 30432 18828
rect 31944 18776 31996 18828
rect 13084 18640 13136 18692
rect 15016 18640 15068 18692
rect 19984 18640 20036 18692
rect 10876 18572 10928 18624
rect 13728 18572 13780 18624
rect 15568 18572 15620 18624
rect 18144 18572 18196 18624
rect 18696 18572 18748 18624
rect 22284 18615 22336 18624
rect 22284 18581 22293 18615
rect 22293 18581 22327 18615
rect 22327 18581 22336 18615
rect 22284 18572 22336 18581
rect 22928 18572 22980 18624
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 26700 18751 26752 18760
rect 25412 18708 25464 18717
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 27620 18708 27672 18760
rect 28540 18708 28592 18760
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 30840 18708 30892 18717
rect 32220 18708 32272 18760
rect 32404 18708 32456 18760
rect 34244 18708 34296 18760
rect 35069 18751 35121 18760
rect 35069 18717 35078 18751
rect 35078 18717 35112 18751
rect 35112 18717 35121 18751
rect 35069 18708 35121 18717
rect 25136 18683 25188 18692
rect 25136 18649 25145 18683
rect 25145 18649 25179 18683
rect 25179 18649 25188 18683
rect 25136 18640 25188 18649
rect 26148 18640 26200 18692
rect 26884 18683 26936 18692
rect 26884 18649 26893 18683
rect 26893 18649 26927 18683
rect 26927 18649 26936 18683
rect 26884 18640 26936 18649
rect 25688 18572 25740 18624
rect 27344 18572 27396 18624
rect 27804 18683 27856 18692
rect 27804 18649 27838 18683
rect 27838 18649 27856 18683
rect 27804 18640 27856 18649
rect 30748 18640 30800 18692
rect 33968 18683 34020 18692
rect 33968 18649 33977 18683
rect 33977 18649 34011 18683
rect 34011 18649 34020 18683
rect 33968 18640 34020 18649
rect 36084 18776 36136 18828
rect 34060 18572 34112 18624
rect 37280 18751 37332 18760
rect 37280 18717 37298 18751
rect 37298 18717 37332 18751
rect 37280 18708 37332 18717
rect 37464 18708 37516 18760
rect 68100 18751 68152 18760
rect 68100 18717 68109 18751
rect 68109 18717 68143 18751
rect 68143 18717 68152 18751
rect 68100 18708 68152 18717
rect 36268 18572 36320 18624
rect 37280 18572 37332 18624
rect 37556 18572 37608 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 6920 18368 6972 18420
rect 10140 18368 10192 18420
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 7656 18343 7708 18352
rect 7656 18309 7665 18343
rect 7665 18309 7699 18343
rect 7699 18309 7708 18343
rect 7656 18300 7708 18309
rect 8852 18300 8904 18352
rect 11980 18300 12032 18352
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 2320 18275 2372 18284
rect 2320 18241 2329 18275
rect 2329 18241 2363 18275
rect 2363 18241 2372 18275
rect 2320 18232 2372 18241
rect 2228 18164 2280 18216
rect 3240 18232 3292 18284
rect 7564 18232 7616 18284
rect 13820 18368 13872 18420
rect 15016 18411 15068 18420
rect 15016 18377 15025 18411
rect 15025 18377 15059 18411
rect 15059 18377 15068 18411
rect 15016 18368 15068 18377
rect 17408 18368 17460 18420
rect 8116 18275 8168 18284
rect 8116 18241 8125 18275
rect 8125 18241 8159 18275
rect 8159 18241 8168 18275
rect 8116 18232 8168 18241
rect 3608 18207 3660 18216
rect 3608 18173 3617 18207
rect 3617 18173 3651 18207
rect 3651 18173 3660 18207
rect 3608 18164 3660 18173
rect 5816 18164 5868 18216
rect 7288 18164 7340 18216
rect 5356 18096 5408 18148
rect 9588 18232 9640 18284
rect 10232 18232 10284 18284
rect 12072 18232 12124 18284
rect 12716 18232 12768 18284
rect 5448 18028 5500 18080
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 15568 18300 15620 18352
rect 17684 18300 17736 18352
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14096 18232 14148 18241
rect 14372 18232 14424 18284
rect 15108 18232 15160 18284
rect 15292 18232 15344 18284
rect 15660 18275 15712 18284
rect 14740 18164 14792 18216
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 15568 18164 15620 18216
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 16856 18232 16908 18284
rect 17316 18232 17368 18284
rect 20720 18300 20772 18352
rect 25412 18368 25464 18420
rect 27804 18411 27856 18420
rect 27804 18377 27813 18411
rect 27813 18377 27847 18411
rect 27847 18377 27856 18411
rect 27804 18368 27856 18377
rect 30748 18411 30800 18420
rect 30748 18377 30757 18411
rect 30757 18377 30791 18411
rect 30791 18377 30800 18411
rect 30748 18368 30800 18377
rect 32588 18368 32640 18420
rect 34244 18411 34296 18420
rect 34244 18377 34253 18411
rect 34253 18377 34287 18411
rect 34287 18377 34296 18411
rect 34244 18368 34296 18377
rect 36452 18411 36504 18420
rect 36452 18377 36461 18411
rect 36461 18377 36495 18411
rect 36495 18377 36504 18411
rect 36452 18368 36504 18377
rect 24216 18300 24268 18352
rect 20628 18232 20680 18284
rect 23020 18232 23072 18284
rect 23756 18275 23808 18284
rect 23756 18241 23765 18275
rect 23765 18241 23799 18275
rect 23799 18241 23808 18275
rect 23756 18232 23808 18241
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 24124 18275 24176 18284
rect 24124 18241 24133 18275
rect 24133 18241 24167 18275
rect 24167 18241 24176 18275
rect 24768 18275 24820 18284
rect 24124 18232 24176 18241
rect 24768 18241 24777 18275
rect 24777 18241 24811 18275
rect 24811 18241 24820 18275
rect 24768 18232 24820 18241
rect 16028 18164 16080 18216
rect 9680 18096 9732 18148
rect 12808 18096 12860 18148
rect 22100 18164 22152 18216
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 10048 18028 10100 18080
rect 11980 18028 12032 18080
rect 14096 18028 14148 18080
rect 17132 18028 17184 18080
rect 17224 18028 17276 18080
rect 17592 18028 17644 18080
rect 24124 18096 24176 18148
rect 26976 18232 27028 18284
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 25780 18207 25832 18216
rect 25780 18173 25789 18207
rect 25789 18173 25823 18207
rect 25823 18173 25832 18207
rect 25780 18164 25832 18173
rect 27988 18232 28040 18284
rect 28540 18275 28592 18284
rect 28540 18241 28549 18275
rect 28549 18241 28583 18275
rect 28583 18241 28592 18275
rect 28540 18232 28592 18241
rect 34428 18300 34480 18352
rect 36084 18343 36136 18352
rect 36084 18309 36093 18343
rect 36093 18309 36127 18343
rect 36127 18309 36136 18343
rect 36084 18300 36136 18309
rect 30104 18275 30156 18284
rect 30104 18241 30119 18275
rect 30119 18241 30153 18275
rect 30153 18241 30156 18275
rect 30288 18275 30340 18284
rect 30104 18232 30156 18241
rect 30288 18241 30297 18275
rect 30297 18241 30331 18275
rect 30331 18241 30340 18275
rect 30288 18232 30340 18241
rect 35072 18275 35124 18284
rect 27712 18164 27764 18216
rect 26148 18096 26200 18148
rect 19524 18028 19576 18080
rect 20996 18028 21048 18080
rect 22560 18028 22612 18080
rect 22744 18028 22796 18080
rect 25136 18028 25188 18080
rect 25872 18028 25924 18080
rect 30380 18096 30432 18148
rect 30288 18028 30340 18080
rect 35072 18241 35081 18275
rect 35081 18241 35115 18275
rect 35115 18241 35124 18275
rect 35072 18232 35124 18241
rect 36268 18275 36320 18284
rect 36268 18241 36277 18275
rect 36277 18241 36311 18275
rect 36311 18241 36320 18275
rect 36268 18232 36320 18241
rect 37464 18232 37516 18284
rect 38016 18275 38068 18284
rect 38016 18241 38050 18275
rect 38050 18241 38068 18275
rect 38016 18232 38068 18241
rect 34796 18207 34848 18216
rect 34796 18173 34805 18207
rect 34805 18173 34839 18207
rect 34839 18173 34848 18207
rect 34796 18164 34848 18173
rect 34060 18096 34112 18148
rect 38752 18028 38804 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 2228 17756 2280 17808
rect 2044 17620 2096 17672
rect 8116 17824 8168 17876
rect 7748 17756 7800 17808
rect 8024 17756 8076 17808
rect 11704 17824 11756 17876
rect 11980 17867 12032 17876
rect 11980 17833 11989 17867
rect 11989 17833 12023 17867
rect 12023 17833 12032 17867
rect 11980 17824 12032 17833
rect 12164 17824 12216 17876
rect 14832 17824 14884 17876
rect 15476 17824 15528 17876
rect 15752 17867 15804 17876
rect 15752 17833 15761 17867
rect 15761 17833 15795 17867
rect 15795 17833 15804 17867
rect 15752 17824 15804 17833
rect 17684 17867 17736 17876
rect 17684 17833 17693 17867
rect 17693 17833 17727 17867
rect 17727 17833 17736 17867
rect 17684 17824 17736 17833
rect 20904 17824 20956 17876
rect 21456 17867 21508 17876
rect 21456 17833 21465 17867
rect 21465 17833 21499 17867
rect 21499 17833 21508 17867
rect 21456 17824 21508 17833
rect 21640 17824 21692 17876
rect 23572 17824 23624 17876
rect 28816 17867 28868 17876
rect 3608 17688 3660 17740
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 7104 17688 7156 17740
rect 9220 17688 9272 17740
rect 2688 17620 2740 17672
rect 6828 17620 6880 17672
rect 2780 17552 2832 17604
rect 2964 17552 3016 17604
rect 2596 17527 2648 17536
rect 2596 17493 2605 17527
rect 2605 17493 2639 17527
rect 2639 17493 2648 17527
rect 2596 17484 2648 17493
rect 2688 17484 2740 17536
rect 5448 17484 5500 17536
rect 6736 17527 6788 17536
rect 6736 17493 6745 17527
rect 6745 17493 6779 17527
rect 6779 17493 6788 17527
rect 6736 17484 6788 17493
rect 7288 17620 7340 17672
rect 9588 17688 9640 17740
rect 9864 17620 9916 17672
rect 10048 17620 10100 17672
rect 10876 17663 10928 17672
rect 10876 17629 10910 17663
rect 10910 17629 10928 17663
rect 10876 17620 10928 17629
rect 14372 17756 14424 17808
rect 16672 17756 16724 17808
rect 16028 17688 16080 17740
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 12992 17663 13044 17672
rect 12992 17629 13001 17663
rect 13001 17629 13035 17663
rect 13035 17629 13044 17663
rect 12992 17620 13044 17629
rect 14740 17663 14792 17672
rect 13452 17552 13504 17604
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 16948 17620 17000 17672
rect 17224 17663 17276 17672
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 16856 17552 16908 17604
rect 17592 17620 17644 17672
rect 20168 17620 20220 17672
rect 20352 17620 20404 17672
rect 20812 17756 20864 17808
rect 22468 17756 22520 17808
rect 28816 17833 28825 17867
rect 28825 17833 28859 17867
rect 28859 17833 28868 17867
rect 28816 17824 28868 17833
rect 29828 17824 29880 17876
rect 33968 17824 34020 17876
rect 26240 17756 26292 17808
rect 29460 17756 29512 17808
rect 32312 17756 32364 17808
rect 34612 17824 34664 17876
rect 36084 17824 36136 17876
rect 38016 17824 38068 17876
rect 34428 17756 34480 17808
rect 24124 17688 24176 17740
rect 25136 17688 25188 17740
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 22008 17663 22060 17672
rect 20812 17620 20864 17629
rect 22008 17629 22017 17663
rect 22017 17629 22051 17663
rect 22051 17629 22060 17663
rect 22008 17620 22060 17629
rect 17776 17552 17828 17604
rect 19432 17552 19484 17604
rect 20536 17552 20588 17604
rect 7564 17484 7616 17536
rect 9772 17527 9824 17536
rect 9772 17493 9781 17527
rect 9781 17493 9815 17527
rect 9815 17493 9824 17527
rect 9772 17484 9824 17493
rect 9864 17484 9916 17536
rect 15200 17484 15252 17536
rect 23020 17552 23072 17604
rect 25688 17620 25740 17672
rect 25964 17688 26016 17740
rect 26056 17663 26108 17672
rect 26056 17629 26064 17663
rect 26064 17629 26098 17663
rect 26098 17629 26108 17663
rect 26056 17620 26108 17629
rect 26148 17663 26200 17672
rect 26148 17629 26157 17663
rect 26157 17629 26191 17663
rect 26191 17629 26200 17663
rect 26148 17620 26200 17629
rect 26700 17620 26752 17672
rect 26792 17663 26844 17672
rect 26792 17629 26801 17663
rect 26801 17629 26835 17663
rect 26835 17629 26844 17663
rect 29368 17688 29420 17740
rect 32220 17731 32272 17740
rect 26792 17620 26844 17629
rect 29092 17620 29144 17672
rect 29736 17663 29788 17672
rect 29736 17629 29745 17663
rect 29745 17629 29779 17663
rect 29779 17629 29788 17663
rect 29736 17620 29788 17629
rect 29828 17663 29880 17672
rect 29828 17629 29837 17663
rect 29837 17629 29871 17663
rect 29871 17629 29880 17663
rect 32220 17697 32229 17731
rect 32229 17697 32263 17731
rect 32263 17697 32272 17731
rect 32220 17688 32272 17697
rect 29828 17620 29880 17629
rect 33324 17620 33376 17672
rect 24584 17552 24636 17604
rect 25780 17595 25832 17604
rect 24124 17484 24176 17536
rect 25136 17484 25188 17536
rect 25504 17527 25556 17536
rect 25504 17493 25513 17527
rect 25513 17493 25547 17527
rect 25547 17493 25556 17527
rect 25504 17484 25556 17493
rect 25780 17561 25789 17595
rect 25789 17561 25823 17595
rect 25823 17561 25832 17595
rect 25780 17552 25832 17561
rect 29276 17552 29328 17604
rect 29920 17595 29972 17604
rect 29920 17561 29929 17595
rect 29929 17561 29963 17595
rect 29963 17561 29972 17595
rect 29920 17552 29972 17561
rect 27160 17484 27212 17536
rect 27988 17527 28040 17536
rect 27988 17493 27997 17527
rect 27997 17493 28031 17527
rect 28031 17493 28040 17527
rect 27988 17484 28040 17493
rect 29552 17527 29604 17536
rect 29552 17493 29561 17527
rect 29561 17493 29595 17527
rect 29595 17493 29604 17527
rect 29552 17484 29604 17493
rect 30840 17527 30892 17536
rect 30840 17493 30849 17527
rect 30849 17493 30883 17527
rect 30883 17493 30892 17527
rect 30840 17484 30892 17493
rect 32404 17484 32456 17536
rect 33876 17663 33928 17672
rect 33876 17629 33885 17663
rect 33885 17629 33919 17663
rect 33919 17629 33928 17663
rect 33876 17620 33928 17629
rect 34336 17620 34388 17672
rect 35992 17552 36044 17604
rect 36728 17552 36780 17604
rect 34796 17484 34848 17536
rect 35808 17484 35860 17536
rect 37740 17552 37792 17604
rect 38660 17663 38712 17672
rect 38660 17629 38669 17663
rect 38669 17629 38703 17663
rect 38703 17629 38712 17663
rect 38660 17620 38712 17629
rect 38844 17663 38896 17672
rect 38844 17629 38853 17663
rect 38853 17629 38887 17663
rect 38887 17629 38896 17663
rect 38844 17620 38896 17629
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 2780 17323 2832 17332
rect 2780 17289 2789 17323
rect 2789 17289 2823 17323
rect 2823 17289 2832 17323
rect 6828 17323 6880 17332
rect 2780 17280 2832 17289
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 7840 17280 7892 17332
rect 2596 17212 2648 17264
rect 8116 17212 8168 17264
rect 12900 17212 12952 17264
rect 15200 17255 15252 17264
rect 15200 17221 15209 17255
rect 15209 17221 15243 17255
rect 15243 17221 15252 17255
rect 15200 17212 15252 17221
rect 15476 17212 15528 17264
rect 16856 17255 16908 17264
rect 16856 17221 16865 17255
rect 16865 17221 16899 17255
rect 16899 17221 16908 17255
rect 16856 17212 16908 17221
rect 24216 17280 24268 17332
rect 1584 17144 1636 17196
rect 2688 17144 2740 17196
rect 3056 17144 3108 17196
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 4620 17144 4672 17196
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 7564 17187 7616 17196
rect 7564 17153 7573 17187
rect 7573 17153 7607 17187
rect 7607 17153 7616 17187
rect 7564 17144 7616 17153
rect 7840 17144 7892 17196
rect 9588 17144 9640 17196
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 13268 17144 13320 17196
rect 17316 17144 17368 17196
rect 3516 17076 3568 17128
rect 14372 17076 14424 17128
rect 20076 17212 20128 17264
rect 20352 17212 20404 17264
rect 20812 17212 20864 17264
rect 21180 17212 21232 17264
rect 25872 17280 25924 17332
rect 25964 17280 26016 17332
rect 24676 17212 24728 17264
rect 27620 17212 27672 17264
rect 32312 17280 32364 17332
rect 32404 17323 32456 17332
rect 32404 17289 32413 17323
rect 32413 17289 32447 17323
rect 32447 17289 32456 17323
rect 32404 17280 32456 17289
rect 33876 17280 33928 17332
rect 38660 17280 38712 17332
rect 18052 17187 18104 17196
rect 18052 17153 18086 17187
rect 18086 17153 18104 17187
rect 19984 17187 20036 17196
rect 18052 17144 18104 17153
rect 19984 17153 19993 17187
rect 19993 17153 20027 17187
rect 20027 17153 20036 17187
rect 19984 17144 20036 17153
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 22008 17144 22060 17196
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 21548 17076 21600 17128
rect 24952 17119 25004 17128
rect 24952 17085 24961 17119
rect 24961 17085 24995 17119
rect 24995 17085 25004 17119
rect 24952 17076 25004 17085
rect 25136 17076 25188 17128
rect 27804 17144 27856 17196
rect 30840 17212 30892 17264
rect 29828 17187 29880 17196
rect 29828 17153 29837 17187
rect 29837 17153 29871 17187
rect 29871 17153 29880 17187
rect 29828 17144 29880 17153
rect 30196 17187 30248 17196
rect 26240 17076 26292 17128
rect 29920 17076 29972 17128
rect 30196 17153 30205 17187
rect 30205 17153 30239 17187
rect 30239 17153 30248 17187
rect 30196 17144 30248 17153
rect 15752 17008 15804 17060
rect 3056 16940 3108 16992
rect 7840 16940 7892 16992
rect 8024 16940 8076 16992
rect 8300 16940 8352 16992
rect 9404 16940 9456 16992
rect 11888 16940 11940 16992
rect 14648 16940 14700 16992
rect 17500 16940 17552 16992
rect 21640 17008 21692 17060
rect 25780 17008 25832 17060
rect 26792 17008 26844 17060
rect 32036 17144 32088 17196
rect 32220 17187 32272 17196
rect 32220 17153 32229 17187
rect 32229 17153 32263 17187
rect 32263 17153 32272 17187
rect 32220 17144 32272 17153
rect 32864 17187 32916 17196
rect 32864 17153 32873 17187
rect 32873 17153 32907 17187
rect 32907 17153 32916 17187
rect 34336 17187 34388 17196
rect 32864 17144 32916 17153
rect 34336 17153 34345 17187
rect 34345 17153 34379 17187
rect 34379 17153 34388 17187
rect 34336 17144 34388 17153
rect 34796 17187 34848 17196
rect 34796 17153 34805 17187
rect 34805 17153 34839 17187
rect 34839 17153 34848 17187
rect 34796 17144 34848 17153
rect 35716 17212 35768 17264
rect 37740 17212 37792 17264
rect 21180 16940 21232 16992
rect 22376 16940 22428 16992
rect 23388 16940 23440 16992
rect 27344 16940 27396 16992
rect 29184 16983 29236 16992
rect 29184 16949 29193 16983
rect 29193 16949 29227 16983
rect 29227 16949 29236 16983
rect 29184 16940 29236 16949
rect 29552 16940 29604 16992
rect 32312 17076 32364 17128
rect 32036 17008 32088 17060
rect 36544 17187 36596 17196
rect 36544 17153 36553 17187
rect 36553 17153 36587 17187
rect 36587 17153 36596 17187
rect 36544 17144 36596 17153
rect 36728 17187 36780 17196
rect 36728 17153 36737 17187
rect 36737 17153 36771 17187
rect 36771 17153 36780 17187
rect 38476 17187 38528 17196
rect 36728 17144 36780 17153
rect 38476 17153 38485 17187
rect 38485 17153 38519 17187
rect 38519 17153 38528 17187
rect 38476 17144 38528 17153
rect 38660 17187 38712 17196
rect 38660 17153 38669 17187
rect 38669 17153 38703 17187
rect 38703 17153 38712 17187
rect 38660 17144 38712 17153
rect 67640 17051 67692 17060
rect 67640 17017 67649 17051
rect 67649 17017 67683 17051
rect 67683 17017 67692 17051
rect 67640 17008 67692 17017
rect 34152 16983 34204 16992
rect 34152 16949 34161 16983
rect 34161 16949 34195 16983
rect 34195 16949 34204 16983
rect 34152 16940 34204 16949
rect 36176 16940 36228 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 2044 16600 2096 16652
rect 3332 16736 3384 16788
rect 8116 16736 8168 16788
rect 10048 16736 10100 16788
rect 11704 16736 11756 16788
rect 13268 16736 13320 16788
rect 14832 16736 14884 16788
rect 2872 16668 2924 16720
rect 3148 16668 3200 16720
rect 3240 16668 3292 16720
rect 5356 16668 5408 16720
rect 9128 16668 9180 16720
rect 3516 16532 3568 16584
rect 9404 16600 9456 16652
rect 10324 16668 10376 16720
rect 13452 16668 13504 16720
rect 15568 16736 15620 16788
rect 18052 16736 18104 16788
rect 18144 16736 18196 16788
rect 17684 16668 17736 16720
rect 19432 16668 19484 16720
rect 9680 16600 9732 16652
rect 12716 16600 12768 16652
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 10600 16532 10652 16584
rect 12808 16532 12860 16584
rect 7380 16464 7432 16516
rect 10968 16464 11020 16516
rect 13544 16532 13596 16584
rect 16764 16600 16816 16652
rect 20536 16600 20588 16652
rect 21548 16600 21600 16652
rect 23020 16668 23072 16720
rect 16948 16532 17000 16584
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 14648 16464 14700 16516
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 19064 16532 19116 16584
rect 17776 16464 17828 16516
rect 20720 16532 20772 16584
rect 23388 16736 23440 16788
rect 27620 16736 27672 16788
rect 27988 16736 28040 16788
rect 30380 16668 30432 16720
rect 32864 16736 32916 16788
rect 36544 16736 36596 16788
rect 35808 16668 35860 16720
rect 24584 16600 24636 16652
rect 27528 16600 27580 16652
rect 22284 16575 22336 16584
rect 22284 16541 22292 16575
rect 22292 16541 22326 16575
rect 22326 16541 22336 16575
rect 22284 16532 22336 16541
rect 22376 16575 22428 16584
rect 22376 16541 22385 16575
rect 22385 16541 22419 16575
rect 22419 16541 22428 16575
rect 22836 16575 22888 16584
rect 22376 16532 22428 16541
rect 22836 16541 22845 16575
rect 22845 16541 22879 16575
rect 22879 16541 22888 16575
rect 22836 16532 22888 16541
rect 24952 16532 25004 16584
rect 26424 16575 26476 16584
rect 26424 16541 26433 16575
rect 26433 16541 26467 16575
rect 26467 16541 26476 16575
rect 26424 16532 26476 16541
rect 29552 16532 29604 16584
rect 29828 16600 29880 16652
rect 32220 16600 32272 16652
rect 35900 16643 35952 16652
rect 29920 16575 29972 16584
rect 29920 16541 29929 16575
rect 29929 16541 29963 16575
rect 29963 16541 29972 16575
rect 29920 16532 29972 16541
rect 30012 16532 30064 16584
rect 30932 16532 30984 16584
rect 32312 16575 32364 16584
rect 32312 16541 32321 16575
rect 32321 16541 32355 16575
rect 32355 16541 32364 16575
rect 32312 16532 32364 16541
rect 35900 16609 35909 16643
rect 35909 16609 35943 16643
rect 35943 16609 35952 16643
rect 35900 16600 35952 16609
rect 34152 16532 34204 16584
rect 36176 16575 36228 16584
rect 21640 16464 21692 16516
rect 2780 16396 2832 16448
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 11612 16396 11664 16448
rect 18972 16396 19024 16448
rect 20720 16396 20772 16448
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 20996 16396 21048 16405
rect 22744 16464 22796 16516
rect 28080 16464 28132 16516
rect 29184 16464 29236 16516
rect 29828 16507 29880 16516
rect 24216 16396 24268 16448
rect 24400 16439 24452 16448
rect 24400 16405 24409 16439
rect 24409 16405 24443 16439
rect 24443 16405 24452 16439
rect 24400 16396 24452 16405
rect 28448 16396 28500 16448
rect 28540 16396 28592 16448
rect 29828 16473 29837 16507
rect 29837 16473 29871 16507
rect 29871 16473 29880 16507
rect 29828 16464 29880 16473
rect 33232 16464 33284 16516
rect 36176 16541 36210 16575
rect 36210 16541 36228 16575
rect 36176 16532 36228 16541
rect 37648 16532 37700 16584
rect 39120 16575 39172 16584
rect 39120 16541 39129 16575
rect 39129 16541 39163 16575
rect 39163 16541 39172 16575
rect 39120 16532 39172 16541
rect 30196 16396 30248 16448
rect 33968 16439 34020 16448
rect 33968 16405 33977 16439
rect 33977 16405 34011 16439
rect 34011 16405 34020 16439
rect 33968 16396 34020 16405
rect 36544 16464 36596 16516
rect 37464 16396 37516 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 3332 16192 3384 16244
rect 5172 16192 5224 16244
rect 7932 16192 7984 16244
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 10968 16235 11020 16244
rect 9772 16192 9824 16201
rect 3792 16167 3844 16176
rect 2044 16056 2096 16108
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 3792 16133 3801 16167
rect 3801 16133 3835 16167
rect 3835 16133 3844 16167
rect 3792 16124 3844 16133
rect 2228 15988 2280 16040
rect 3700 16056 3752 16108
rect 4528 16099 4580 16108
rect 4528 16065 4537 16099
rect 4537 16065 4571 16099
rect 4571 16065 4580 16099
rect 4528 16056 4580 16065
rect 4807 16099 4859 16108
rect 4807 16065 4816 16099
rect 4816 16065 4850 16099
rect 4850 16065 4859 16099
rect 4807 16056 4859 16065
rect 5356 16056 5408 16108
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 9680 16124 9732 16176
rect 8024 16099 8076 16108
rect 8024 16065 8058 16099
rect 8058 16065 8076 16099
rect 8024 16056 8076 16065
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 10416 16056 10468 16108
rect 10968 16201 10977 16235
rect 10977 16201 11011 16235
rect 11011 16201 11020 16235
rect 10968 16192 11020 16201
rect 11336 16192 11388 16244
rect 19248 16192 19300 16244
rect 19432 16192 19484 16244
rect 12072 16124 12124 16176
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 16672 16124 16724 16176
rect 16856 16124 16908 16176
rect 20904 16192 20956 16244
rect 21824 16192 21876 16244
rect 2596 15920 2648 15972
rect 10508 15920 10560 15972
rect 12992 15988 13044 16040
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 14648 16099 14700 16108
rect 13912 16056 13964 16065
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 16120 16056 16172 16108
rect 21732 16124 21784 16176
rect 14832 15988 14884 16040
rect 16764 15988 16816 16040
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 20904 16056 20956 16108
rect 22836 16192 22888 16244
rect 25136 16192 25188 16244
rect 27804 16192 27856 16244
rect 28080 16235 28132 16244
rect 28080 16201 28089 16235
rect 28089 16201 28123 16235
rect 28123 16201 28132 16235
rect 28080 16192 28132 16201
rect 28172 16192 28224 16244
rect 33968 16192 34020 16244
rect 36544 16235 36596 16244
rect 24400 16124 24452 16176
rect 22192 16099 22244 16108
rect 20444 15988 20496 16040
rect 21088 15988 21140 16040
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 23020 16099 23072 16108
rect 22468 16056 22520 16065
rect 23020 16065 23029 16099
rect 23029 16065 23063 16099
rect 23063 16065 23072 16099
rect 23020 16056 23072 16065
rect 23480 16056 23532 16108
rect 25872 16056 25924 16108
rect 26976 16099 27028 16108
rect 26976 16065 26985 16099
rect 26985 16065 27019 16099
rect 27019 16065 27028 16099
rect 26976 16056 27028 16065
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27712 16124 27764 16176
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 28632 16124 28684 16176
rect 30840 16124 30892 16176
rect 27344 16056 27396 16065
rect 28724 16099 28776 16108
rect 23848 15988 23900 16040
rect 13728 15920 13780 15972
rect 15016 15920 15068 15972
rect 19616 15920 19668 15972
rect 22468 15920 22520 15972
rect 23020 15920 23072 15972
rect 5264 15852 5316 15904
rect 5448 15852 5500 15904
rect 7380 15852 7432 15904
rect 8944 15852 8996 15904
rect 12440 15852 12492 15904
rect 14924 15852 14976 15904
rect 16212 15852 16264 15904
rect 16764 15852 16816 15904
rect 17592 15852 17644 15904
rect 18972 15895 19024 15904
rect 18972 15861 18981 15895
rect 18981 15861 19015 15895
rect 19015 15861 19024 15895
rect 18972 15852 19024 15861
rect 20352 15852 20404 15904
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 23572 15852 23624 15904
rect 26424 15852 26476 15904
rect 28448 15920 28500 15972
rect 28724 16065 28733 16099
rect 28733 16065 28767 16099
rect 28767 16065 28776 16099
rect 28724 16056 28776 16065
rect 29920 16099 29972 16108
rect 29920 16065 29929 16099
rect 29929 16065 29963 16099
rect 29963 16065 29972 16099
rect 29920 16056 29972 16065
rect 30932 16099 30984 16108
rect 30932 16065 30941 16099
rect 30941 16065 30975 16099
rect 30975 16065 30984 16099
rect 30932 16056 30984 16065
rect 31300 16099 31352 16108
rect 31300 16065 31309 16099
rect 31309 16065 31343 16099
rect 31343 16065 31352 16099
rect 31300 16056 31352 16065
rect 32680 16056 32732 16108
rect 36544 16201 36553 16235
rect 36553 16201 36587 16235
rect 36587 16201 36596 16235
rect 36544 16192 36596 16201
rect 31208 15988 31260 16040
rect 34612 16099 34664 16108
rect 34612 16065 34621 16099
rect 34621 16065 34655 16099
rect 34655 16065 34664 16099
rect 34612 16056 34664 16065
rect 35992 16056 36044 16108
rect 37648 16167 37700 16176
rect 37648 16133 37657 16167
rect 37657 16133 37691 16167
rect 37691 16133 37700 16167
rect 37648 16124 37700 16133
rect 38476 16124 38528 16176
rect 37464 16099 37516 16108
rect 35716 15988 35768 16040
rect 29092 15920 29144 15972
rect 30288 15920 30340 15972
rect 37464 16065 37473 16099
rect 37473 16065 37507 16099
rect 37507 16065 37516 16099
rect 37464 16056 37516 16065
rect 30748 15895 30800 15904
rect 30748 15861 30757 15895
rect 30757 15861 30791 15895
rect 30791 15861 30800 15895
rect 30748 15852 30800 15861
rect 32312 15895 32364 15904
rect 32312 15861 32321 15895
rect 32321 15861 32355 15895
rect 32355 15861 32364 15895
rect 32312 15852 32364 15861
rect 67640 15895 67692 15904
rect 67640 15861 67649 15895
rect 67649 15861 67683 15895
rect 67683 15861 67692 15895
rect 67640 15852 67692 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 2964 15691 3016 15700
rect 2964 15657 2973 15691
rect 2973 15657 3007 15691
rect 3007 15657 3016 15691
rect 2964 15648 3016 15657
rect 5172 15648 5224 15700
rect 6644 15648 6696 15700
rect 7656 15691 7708 15700
rect 7656 15657 7665 15691
rect 7665 15657 7699 15691
rect 7699 15657 7708 15691
rect 7656 15648 7708 15657
rect 7932 15648 7984 15700
rect 9404 15648 9456 15700
rect 11336 15648 11388 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 15384 15691 15436 15700
rect 15384 15657 15393 15691
rect 15393 15657 15427 15691
rect 15427 15657 15436 15691
rect 15384 15648 15436 15657
rect 2044 15444 2096 15496
rect 1584 15376 1636 15428
rect 1676 15419 1728 15428
rect 1676 15385 1685 15419
rect 1685 15385 1719 15419
rect 1719 15385 1728 15419
rect 1676 15376 1728 15385
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4068 15444 4120 15496
rect 5264 15487 5316 15496
rect 5264 15453 5298 15487
rect 5298 15453 5316 15487
rect 5264 15444 5316 15453
rect 9496 15623 9548 15632
rect 7012 15512 7064 15564
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 7840 15512 7892 15564
rect 8024 15444 8076 15496
rect 8944 15487 8996 15496
rect 8944 15453 8953 15487
rect 8953 15453 8987 15487
rect 8987 15453 8996 15487
rect 8944 15444 8996 15453
rect 9496 15589 9505 15623
rect 9505 15589 9539 15623
rect 9539 15589 9548 15623
rect 9496 15580 9548 15589
rect 17040 15512 17092 15564
rect 17776 15580 17828 15632
rect 19708 15648 19760 15700
rect 20168 15648 20220 15700
rect 20260 15648 20312 15700
rect 21456 15691 21508 15700
rect 21456 15657 21465 15691
rect 21465 15657 21499 15691
rect 21499 15657 21508 15691
rect 21456 15648 21508 15657
rect 22376 15691 22428 15700
rect 22376 15657 22385 15691
rect 22385 15657 22419 15691
rect 22419 15657 22428 15691
rect 22376 15648 22428 15657
rect 22836 15648 22888 15700
rect 27344 15648 27396 15700
rect 34612 15648 34664 15700
rect 19984 15580 20036 15632
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 11796 15444 11848 15496
rect 7012 15376 7064 15428
rect 7288 15419 7340 15428
rect 7288 15385 7297 15419
rect 7297 15385 7331 15419
rect 7331 15385 7340 15419
rect 7288 15376 7340 15385
rect 7840 15376 7892 15428
rect 8208 15419 8260 15428
rect 8208 15385 8217 15419
rect 8217 15385 8251 15419
rect 8251 15385 8260 15419
rect 8208 15376 8260 15385
rect 9128 15419 9180 15428
rect 9128 15385 9137 15419
rect 9137 15385 9171 15419
rect 9171 15385 9180 15419
rect 9128 15376 9180 15385
rect 13452 15419 13504 15428
rect 13452 15385 13461 15419
rect 13461 15385 13495 15419
rect 13495 15385 13504 15419
rect 13452 15376 13504 15385
rect 16764 15444 16816 15496
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 17592 15512 17644 15564
rect 19616 15512 19668 15564
rect 15476 15376 15528 15428
rect 17868 15444 17920 15496
rect 19064 15444 19116 15496
rect 19156 15444 19208 15496
rect 19340 15444 19392 15496
rect 19708 15444 19760 15496
rect 20168 15444 20220 15496
rect 20444 15512 20496 15564
rect 21456 15512 21508 15564
rect 22008 15512 22060 15564
rect 24216 15512 24268 15564
rect 29552 15580 29604 15632
rect 38660 15648 38712 15700
rect 20352 15487 20404 15496
rect 20352 15453 20361 15487
rect 20361 15453 20395 15487
rect 20395 15453 20404 15487
rect 20352 15444 20404 15453
rect 21732 15444 21784 15496
rect 22928 15444 22980 15496
rect 23112 15487 23164 15496
rect 23112 15453 23121 15487
rect 23121 15453 23155 15487
rect 23155 15453 23164 15487
rect 23112 15444 23164 15453
rect 26332 15444 26384 15496
rect 26700 15444 26752 15496
rect 27068 15444 27120 15496
rect 17684 15376 17736 15428
rect 3148 15308 3200 15360
rect 3976 15308 4028 15360
rect 8944 15308 8996 15360
rect 12624 15308 12676 15360
rect 14556 15308 14608 15360
rect 15200 15351 15252 15360
rect 15200 15317 15209 15351
rect 15209 15317 15243 15351
rect 15243 15317 15252 15351
rect 15200 15308 15252 15317
rect 17960 15308 18012 15360
rect 19340 15308 19392 15360
rect 20536 15376 20588 15428
rect 20260 15308 20312 15360
rect 21088 15308 21140 15360
rect 22100 15419 22152 15428
rect 22100 15385 22109 15419
rect 22109 15385 22143 15419
rect 22143 15385 22152 15419
rect 22100 15376 22152 15385
rect 22744 15376 22796 15428
rect 23480 15376 23532 15428
rect 27712 15376 27764 15428
rect 28172 15444 28224 15496
rect 29828 15444 29880 15496
rect 30196 15512 30248 15564
rect 34704 15512 34756 15564
rect 30472 15444 30524 15496
rect 32312 15444 32364 15496
rect 34152 15487 34204 15496
rect 34152 15453 34161 15487
rect 34161 15453 34195 15487
rect 34195 15453 34204 15487
rect 34152 15444 34204 15453
rect 35992 15580 36044 15632
rect 22192 15308 22244 15360
rect 22376 15308 22428 15360
rect 28264 15351 28316 15360
rect 28264 15317 28273 15351
rect 28273 15317 28307 15351
rect 28307 15317 28316 15351
rect 28264 15308 28316 15317
rect 28632 15308 28684 15360
rect 29920 15308 29972 15360
rect 32772 15376 32824 15428
rect 39120 15512 39172 15564
rect 30472 15308 30524 15360
rect 34612 15308 34664 15360
rect 35716 15376 35768 15428
rect 36176 15308 36228 15360
rect 37556 15351 37608 15360
rect 37556 15317 37565 15351
rect 37565 15317 37599 15351
rect 37599 15317 37608 15351
rect 37556 15308 37608 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 7472 15104 7524 15156
rect 10416 15104 10468 15156
rect 10508 15104 10560 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 2780 14968 2832 15020
rect 3148 14968 3200 15020
rect 3700 15011 3752 15020
rect 3700 14977 3709 15011
rect 3709 14977 3743 15011
rect 3743 14977 3752 15011
rect 3700 14968 3752 14977
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 4804 15036 4856 15088
rect 5172 15036 5224 15088
rect 7288 15036 7340 15088
rect 8024 15079 8076 15088
rect 8024 15045 8033 15079
rect 8033 15045 8067 15079
rect 8067 15045 8076 15079
rect 8024 15036 8076 15045
rect 6184 14968 6236 15020
rect 6736 14968 6788 15020
rect 7012 15011 7064 15020
rect 7012 14977 7021 15011
rect 7021 14977 7055 15011
rect 7055 14977 7064 15011
rect 7012 14968 7064 14977
rect 2228 14900 2280 14952
rect 2596 14900 2648 14952
rect 2964 14900 3016 14952
rect 1676 14832 1728 14884
rect 6828 14900 6880 14952
rect 8300 14968 8352 15020
rect 8208 14832 8260 14884
rect 4620 14764 4672 14816
rect 9772 14968 9824 15020
rect 10324 15011 10376 15020
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 12440 15036 12492 15088
rect 10692 15011 10744 15020
rect 10692 14977 10721 15011
rect 10721 14977 10744 15011
rect 10692 14968 10744 14977
rect 10968 14968 11020 15020
rect 15016 15104 15068 15156
rect 18972 15104 19024 15156
rect 12900 15036 12952 15088
rect 15384 15036 15436 15088
rect 11612 14900 11664 14952
rect 11704 14900 11756 14952
rect 14372 14900 14424 14952
rect 12532 14832 12584 14884
rect 11520 14764 11572 14816
rect 14832 14968 14884 15020
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 17960 15036 18012 15088
rect 20352 15104 20404 15156
rect 20720 15104 20772 15156
rect 20812 15036 20864 15088
rect 22652 15104 22704 15156
rect 28540 15104 28592 15156
rect 29552 15147 29604 15156
rect 29552 15113 29561 15147
rect 29561 15113 29595 15147
rect 29595 15113 29604 15147
rect 29552 15104 29604 15113
rect 30380 15147 30432 15156
rect 30380 15113 30389 15147
rect 30389 15113 30423 15147
rect 30423 15113 30432 15147
rect 30380 15104 30432 15113
rect 36176 15147 36228 15156
rect 36176 15113 36185 15147
rect 36185 15113 36219 15147
rect 36219 15113 36228 15147
rect 36176 15104 36228 15113
rect 39304 15104 39356 15156
rect 40224 15104 40276 15156
rect 21364 15036 21416 15088
rect 20628 14968 20680 15020
rect 24308 15036 24360 15088
rect 22836 14968 22888 15020
rect 23020 15011 23072 15020
rect 23020 14977 23054 15011
rect 23054 14977 23072 15011
rect 23020 14968 23072 14977
rect 26700 14968 26752 15020
rect 28264 15036 28316 15088
rect 32312 15036 32364 15088
rect 34704 15036 34756 15088
rect 35348 15036 35400 15088
rect 21916 14943 21968 14952
rect 16120 14875 16172 14884
rect 16120 14841 16129 14875
rect 16129 14841 16163 14875
rect 16163 14841 16172 14875
rect 16120 14832 16172 14841
rect 17868 14832 17920 14884
rect 21916 14909 21925 14943
rect 21925 14909 21959 14943
rect 21959 14909 21968 14943
rect 21916 14900 21968 14909
rect 22008 14900 22060 14952
rect 26792 14900 26844 14952
rect 16672 14764 16724 14816
rect 18144 14764 18196 14816
rect 18604 14764 18656 14816
rect 21180 14764 21232 14816
rect 22652 14832 22704 14884
rect 24768 14875 24820 14884
rect 24768 14841 24777 14875
rect 24777 14841 24811 14875
rect 24811 14841 24820 14875
rect 24768 14832 24820 14841
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 22284 14807 22336 14816
rect 22284 14773 22293 14807
rect 22293 14773 22327 14807
rect 22327 14773 22336 14807
rect 22284 14764 22336 14773
rect 23940 14764 23992 14816
rect 26424 14764 26476 14816
rect 28724 14968 28776 15020
rect 30748 14968 30800 15020
rect 30932 14968 30984 15020
rect 31208 15011 31260 15020
rect 31208 14977 31217 15011
rect 31217 14977 31251 15011
rect 31251 14977 31260 15011
rect 31208 14968 31260 14977
rect 31484 14968 31536 15020
rect 32956 14968 33008 15020
rect 37556 15036 37608 15088
rect 37648 14968 37700 15020
rect 27528 14900 27580 14952
rect 27712 14832 27764 14884
rect 30932 14832 30984 14884
rect 34612 14832 34664 14884
rect 30840 14807 30892 14816
rect 30840 14773 30849 14807
rect 30849 14773 30883 14807
rect 30883 14773 30892 14807
rect 30840 14764 30892 14773
rect 32680 14764 32732 14816
rect 35900 14764 35952 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 3884 14560 3936 14612
rect 8116 14560 8168 14612
rect 8944 14560 8996 14612
rect 6184 14492 6236 14544
rect 3792 14424 3844 14476
rect 7564 14492 7616 14544
rect 10508 14492 10560 14544
rect 4068 14356 4120 14408
rect 4620 14356 4672 14408
rect 4804 14356 4856 14408
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 6828 14356 6880 14408
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 7288 14399 7340 14408
rect 7288 14365 7317 14399
rect 7317 14365 7340 14399
rect 10784 14424 10836 14476
rect 8944 14399 8996 14408
rect 7288 14356 7340 14365
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 9312 14356 9364 14408
rect 14280 14603 14332 14612
rect 11520 14535 11572 14544
rect 11520 14501 11529 14535
rect 11529 14501 11563 14535
rect 11563 14501 11572 14535
rect 11520 14492 11572 14501
rect 11796 14492 11848 14544
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 12992 14492 13044 14544
rect 14924 14560 14976 14612
rect 16580 14603 16632 14612
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 17132 14560 17184 14612
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 20536 14560 20588 14612
rect 22376 14560 22428 14612
rect 24676 14603 24728 14612
rect 24676 14569 24685 14603
rect 24685 14569 24719 14603
rect 24719 14569 24728 14603
rect 24676 14560 24728 14569
rect 26700 14603 26752 14612
rect 26700 14569 26709 14603
rect 26709 14569 26743 14603
rect 26743 14569 26752 14603
rect 26700 14560 26752 14569
rect 26792 14560 26844 14612
rect 27436 14560 27488 14612
rect 28172 14560 28224 14612
rect 28724 14560 28776 14612
rect 33048 14560 33100 14612
rect 12900 14467 12952 14476
rect 12900 14433 12909 14467
rect 12909 14433 12943 14467
rect 12943 14433 12952 14467
rect 12900 14424 12952 14433
rect 12072 14356 12124 14408
rect 16304 14492 16356 14544
rect 6460 14288 6512 14340
rect 8300 14288 8352 14340
rect 9680 14288 9732 14340
rect 14924 14399 14976 14408
rect 12532 14288 12584 14340
rect 14924 14365 14933 14399
rect 14933 14365 14967 14399
rect 14967 14365 14976 14399
rect 14924 14356 14976 14365
rect 28908 14492 28960 14544
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 19984 14424 20036 14476
rect 20904 14467 20956 14476
rect 20904 14433 20913 14467
rect 20913 14433 20947 14467
rect 20947 14433 20956 14467
rect 20904 14424 20956 14433
rect 21640 14424 21692 14476
rect 24492 14467 24544 14476
rect 22744 14356 22796 14408
rect 19340 14288 19392 14340
rect 1584 14220 1636 14272
rect 2320 14263 2372 14272
rect 2320 14229 2329 14263
rect 2329 14229 2363 14263
rect 2363 14229 2372 14263
rect 2320 14220 2372 14229
rect 7104 14220 7156 14272
rect 7656 14220 7708 14272
rect 11704 14220 11756 14272
rect 12716 14220 12768 14272
rect 14464 14220 14516 14272
rect 15844 14263 15896 14272
rect 15844 14229 15853 14263
rect 15853 14229 15887 14263
rect 15887 14229 15896 14263
rect 15844 14220 15896 14229
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 19432 14220 19484 14272
rect 20720 14288 20772 14340
rect 20996 14288 21048 14340
rect 24124 14288 24176 14340
rect 24492 14433 24501 14467
rect 24501 14433 24535 14467
rect 24535 14433 24544 14467
rect 24492 14424 24544 14433
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 28448 14424 28500 14476
rect 30472 14424 30524 14476
rect 26332 14331 26384 14340
rect 26332 14297 26341 14331
rect 26341 14297 26375 14331
rect 26375 14297 26384 14331
rect 26332 14288 26384 14297
rect 28080 14399 28132 14408
rect 28080 14365 28089 14399
rect 28089 14365 28123 14399
rect 28123 14365 28132 14399
rect 28080 14356 28132 14365
rect 28264 14356 28316 14408
rect 31208 14356 31260 14408
rect 31392 14356 31444 14408
rect 31852 14399 31904 14408
rect 31852 14365 31861 14399
rect 31861 14365 31895 14399
rect 31895 14365 31904 14399
rect 31852 14356 31904 14365
rect 20076 14220 20128 14272
rect 22192 14220 22244 14272
rect 23388 14220 23440 14272
rect 24768 14220 24820 14272
rect 27988 14220 28040 14272
rect 30564 14220 30616 14272
rect 33140 14492 33192 14544
rect 33140 14399 33192 14408
rect 33140 14365 33149 14399
rect 33149 14365 33183 14399
rect 33183 14365 33192 14399
rect 33140 14356 33192 14365
rect 39948 14560 40000 14612
rect 35808 14356 35860 14408
rect 37096 14399 37148 14408
rect 37096 14365 37105 14399
rect 37105 14365 37139 14399
rect 37139 14365 37148 14399
rect 37096 14356 37148 14365
rect 38844 14399 38896 14408
rect 38844 14365 38873 14399
rect 38873 14365 38896 14399
rect 38844 14356 38896 14365
rect 39028 14356 39080 14408
rect 39396 14356 39448 14408
rect 33324 14331 33376 14340
rect 33324 14297 33333 14331
rect 33333 14297 33367 14331
rect 33367 14297 33376 14331
rect 33324 14288 33376 14297
rect 34612 14288 34664 14340
rect 33416 14220 33468 14272
rect 34796 14220 34848 14272
rect 35164 14288 35216 14340
rect 35440 14288 35492 14340
rect 39764 14288 39816 14340
rect 40224 14399 40276 14408
rect 40224 14365 40253 14399
rect 40253 14365 40276 14399
rect 68100 14399 68152 14408
rect 40224 14356 40276 14365
rect 68100 14365 68109 14399
rect 68109 14365 68143 14399
rect 68143 14365 68152 14399
rect 68100 14356 68152 14365
rect 40500 14331 40552 14340
rect 36452 14220 36504 14272
rect 40500 14297 40509 14331
rect 40509 14297 40543 14331
rect 40543 14297 40552 14331
rect 40500 14288 40552 14297
rect 40316 14220 40368 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 5540 14016 5592 14068
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 6460 14016 6512 14068
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 7748 14016 7800 14068
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 2780 13948 2832 14000
rect 2228 13812 2280 13864
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 7196 13948 7248 14000
rect 2964 13812 3016 13864
rect 2780 13744 2832 13796
rect 4620 13812 4672 13864
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 8300 13948 8352 14000
rect 11520 13948 11572 14000
rect 11888 13991 11940 14000
rect 11888 13957 11897 13991
rect 11897 13957 11931 13991
rect 11931 13957 11940 13991
rect 11888 13948 11940 13957
rect 6552 13812 6604 13864
rect 9128 13880 9180 13932
rect 9864 13880 9916 13932
rect 10600 13923 10652 13932
rect 10600 13889 10609 13923
rect 10609 13889 10643 13923
rect 10643 13889 10652 13923
rect 10600 13880 10652 13889
rect 10784 13880 10836 13932
rect 11612 13923 11664 13932
rect 11612 13889 11621 13923
rect 11621 13889 11655 13923
rect 11655 13889 11664 13923
rect 11612 13880 11664 13889
rect 11704 13880 11756 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 14464 13948 14516 14000
rect 14648 13991 14700 14000
rect 14648 13957 14657 13991
rect 14657 13957 14691 13991
rect 14691 13957 14700 13991
rect 14648 13948 14700 13957
rect 15476 14016 15528 14068
rect 15844 14016 15896 14068
rect 19892 14016 19944 14068
rect 20996 14016 21048 14068
rect 21916 14016 21968 14068
rect 22836 14016 22888 14068
rect 33048 14016 33100 14068
rect 17408 13948 17460 14000
rect 23940 13948 23992 14000
rect 25412 13948 25464 14000
rect 26424 13991 26476 14000
rect 26424 13957 26433 13991
rect 26433 13957 26467 13991
rect 26467 13957 26476 13991
rect 26424 13948 26476 13957
rect 32956 13948 33008 14000
rect 34612 13948 34664 14000
rect 35440 14016 35492 14068
rect 39304 14059 39356 14068
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 14188 13880 14240 13932
rect 15292 13880 15344 13932
rect 15844 13880 15896 13932
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 14740 13812 14792 13864
rect 15476 13812 15528 13864
rect 20536 13880 20588 13932
rect 20904 13923 20956 13932
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 19616 13812 19668 13864
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 21272 13880 21324 13932
rect 21548 13880 21600 13932
rect 14096 13787 14148 13796
rect 14096 13753 14105 13787
rect 14105 13753 14139 13787
rect 14139 13753 14148 13787
rect 14096 13744 14148 13753
rect 14280 13744 14332 13796
rect 17960 13744 18012 13796
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 23848 13880 23900 13932
rect 24124 13880 24176 13932
rect 28632 13880 28684 13932
rect 28448 13855 28500 13864
rect 28448 13821 28457 13855
rect 28457 13821 28491 13855
rect 28491 13821 28500 13855
rect 28448 13812 28500 13821
rect 30288 13855 30340 13864
rect 30288 13821 30297 13855
rect 30297 13821 30331 13855
rect 30331 13821 30340 13855
rect 30288 13812 30340 13821
rect 30748 13880 30800 13932
rect 31392 13923 31444 13932
rect 31392 13889 31401 13923
rect 31401 13889 31435 13923
rect 31435 13889 31444 13923
rect 31392 13880 31444 13889
rect 31576 13923 31628 13932
rect 31576 13889 31585 13923
rect 31585 13889 31619 13923
rect 31619 13889 31628 13923
rect 31576 13880 31628 13889
rect 33048 13923 33100 13932
rect 33048 13889 33057 13923
rect 33057 13889 33091 13923
rect 33091 13889 33100 13923
rect 33048 13880 33100 13889
rect 33324 13880 33376 13932
rect 33600 13880 33652 13932
rect 36452 13948 36504 14000
rect 23388 13744 23440 13796
rect 24308 13744 24360 13796
rect 32864 13744 32916 13796
rect 3884 13676 3936 13728
rect 8760 13676 8812 13728
rect 10876 13676 10928 13728
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 14556 13676 14608 13728
rect 21640 13676 21692 13728
rect 23664 13676 23716 13728
rect 27160 13676 27212 13728
rect 27896 13719 27948 13728
rect 27896 13685 27905 13719
rect 27905 13685 27939 13719
rect 27939 13685 27948 13719
rect 27896 13676 27948 13685
rect 28080 13676 28132 13728
rect 31024 13719 31076 13728
rect 31024 13685 31033 13719
rect 31033 13685 31067 13719
rect 31067 13685 31076 13719
rect 31024 13676 31076 13685
rect 34796 13880 34848 13932
rect 35072 13923 35124 13932
rect 35072 13889 35081 13923
rect 35081 13889 35115 13923
rect 35115 13889 35124 13923
rect 35072 13880 35124 13889
rect 35532 13880 35584 13932
rect 36176 13923 36228 13932
rect 36176 13889 36185 13923
rect 36185 13889 36219 13923
rect 36219 13889 36228 13923
rect 36176 13880 36228 13889
rect 35900 13855 35952 13864
rect 35900 13821 35909 13855
rect 35909 13821 35943 13855
rect 35943 13821 35952 13855
rect 35900 13812 35952 13821
rect 36360 13923 36412 13932
rect 36360 13889 36369 13923
rect 36369 13889 36403 13923
rect 36403 13889 36412 13923
rect 39304 14025 39313 14059
rect 39313 14025 39347 14059
rect 39347 14025 39356 14059
rect 39304 14016 39356 14025
rect 39764 14016 39816 14068
rect 39948 13991 40000 14000
rect 39948 13957 39957 13991
rect 39957 13957 39991 13991
rect 39991 13957 40000 13991
rect 39948 13948 40000 13957
rect 36360 13880 36412 13889
rect 39396 13880 39448 13932
rect 39764 13923 39816 13932
rect 39764 13889 39773 13923
rect 39773 13889 39807 13923
rect 39807 13889 39816 13923
rect 39764 13880 39816 13889
rect 34244 13676 34296 13728
rect 35164 13676 35216 13728
rect 35532 13676 35584 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 11428 13472 11480 13524
rect 2688 13404 2740 13456
rect 4068 13336 4120 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 2596 13268 2648 13320
rect 4620 13268 4672 13320
rect 12072 13404 12124 13456
rect 14280 13447 14332 13456
rect 14280 13413 14289 13447
rect 14289 13413 14323 13447
rect 14323 13413 14332 13447
rect 14280 13404 14332 13413
rect 17408 13472 17460 13524
rect 21088 13472 21140 13524
rect 21180 13472 21232 13524
rect 21640 13472 21692 13524
rect 8300 13336 8352 13388
rect 11520 13336 11572 13388
rect 13084 13336 13136 13388
rect 14004 13336 14056 13388
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 15384 13379 15436 13388
rect 15384 13345 15393 13379
rect 15393 13345 15427 13379
rect 15427 13345 15436 13379
rect 15384 13336 15436 13345
rect 21456 13404 21508 13456
rect 18880 13336 18932 13388
rect 20536 13336 20588 13388
rect 7932 13268 7984 13320
rect 10140 13268 10192 13320
rect 10968 13268 11020 13320
rect 11704 13268 11756 13320
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 19340 13268 19392 13320
rect 21272 13336 21324 13388
rect 21916 13336 21968 13388
rect 8024 13200 8076 13252
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 8300 13200 8352 13252
rect 8392 13243 8444 13252
rect 8392 13209 8401 13243
rect 8401 13209 8435 13243
rect 8435 13209 8444 13243
rect 8392 13200 8444 13209
rect 11060 13200 11112 13252
rect 17592 13200 17644 13252
rect 9864 13132 9916 13184
rect 21732 13268 21784 13320
rect 22560 13472 22612 13524
rect 23020 13472 23072 13524
rect 28632 13472 28684 13524
rect 32864 13515 32916 13524
rect 32864 13481 32873 13515
rect 32873 13481 32907 13515
rect 32907 13481 32916 13515
rect 32864 13472 32916 13481
rect 35808 13472 35860 13524
rect 22744 13404 22796 13456
rect 25504 13404 25556 13456
rect 29828 13404 29880 13456
rect 30288 13404 30340 13456
rect 23388 13336 23440 13388
rect 26792 13379 26844 13388
rect 26792 13345 26801 13379
rect 26801 13345 26835 13379
rect 26835 13345 26844 13379
rect 26792 13336 26844 13345
rect 29644 13336 29696 13388
rect 31852 13404 31904 13456
rect 32312 13404 32364 13456
rect 32588 13404 32640 13456
rect 33416 13404 33468 13456
rect 34796 13404 34848 13456
rect 34888 13404 34940 13456
rect 36176 13447 36228 13456
rect 36176 13413 36185 13447
rect 36185 13413 36219 13447
rect 36219 13413 36228 13447
rect 36176 13404 36228 13413
rect 40132 13404 40184 13456
rect 23664 13311 23716 13320
rect 23664 13277 23673 13311
rect 23673 13277 23707 13311
rect 23707 13277 23716 13311
rect 23664 13268 23716 13277
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 25044 13268 25096 13320
rect 29828 13268 29880 13320
rect 30472 13268 30524 13320
rect 30748 13311 30800 13320
rect 30748 13277 30757 13311
rect 30757 13277 30791 13311
rect 30791 13277 30800 13311
rect 30748 13268 30800 13277
rect 33048 13311 33100 13320
rect 33048 13277 33057 13311
rect 33057 13277 33091 13311
rect 33091 13277 33100 13311
rect 33048 13268 33100 13277
rect 36360 13336 36412 13388
rect 39120 13336 39172 13388
rect 20996 13243 21048 13252
rect 20996 13209 21005 13243
rect 21005 13209 21039 13243
rect 21039 13209 21048 13243
rect 20996 13200 21048 13209
rect 23940 13200 23992 13252
rect 24124 13200 24176 13252
rect 24676 13200 24728 13252
rect 18052 13132 18104 13184
rect 24032 13132 24084 13184
rect 24952 13175 25004 13184
rect 24952 13141 24961 13175
rect 24961 13141 24995 13175
rect 24995 13141 25004 13175
rect 24952 13132 25004 13141
rect 25688 13200 25740 13252
rect 27620 13200 27672 13252
rect 30012 13243 30064 13252
rect 30012 13209 30021 13243
rect 30021 13209 30055 13243
rect 30055 13209 30064 13243
rect 30012 13200 30064 13209
rect 30380 13200 30432 13252
rect 33324 13200 33376 13252
rect 29828 13132 29880 13184
rect 33048 13132 33100 13184
rect 35716 13268 35768 13320
rect 39304 13268 39356 13320
rect 40500 13311 40552 13320
rect 40500 13277 40509 13311
rect 40509 13277 40543 13311
rect 40543 13277 40552 13311
rect 40500 13268 40552 13277
rect 34704 13200 34756 13252
rect 35532 13200 35584 13252
rect 39948 13200 40000 13252
rect 68100 13311 68152 13320
rect 68100 13277 68109 13311
rect 68109 13277 68143 13311
rect 68143 13277 68152 13311
rect 68100 13268 68152 13277
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 4068 12928 4120 12980
rect 5356 12928 5408 12980
rect 8024 12971 8076 12980
rect 2320 12792 2372 12844
rect 3792 12835 3844 12844
rect 1400 12588 1452 12640
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 3884 12792 3936 12844
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 12164 12928 12216 12980
rect 8300 12860 8352 12912
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7196 12792 7248 12844
rect 8116 12792 8168 12844
rect 8392 12792 8444 12844
rect 9680 12860 9732 12912
rect 11060 12860 11112 12912
rect 11704 12860 11756 12912
rect 12072 12903 12124 12912
rect 12072 12869 12081 12903
rect 12081 12869 12115 12903
rect 12115 12869 12124 12903
rect 12072 12860 12124 12869
rect 8760 12835 8812 12844
rect 8760 12801 8794 12835
rect 8794 12801 8812 12835
rect 11796 12835 11848 12844
rect 8760 12792 8812 12801
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 11888 12724 11940 12776
rect 13360 12928 13412 12980
rect 15108 12971 15160 12980
rect 15108 12937 15117 12971
rect 15117 12937 15151 12971
rect 15151 12937 15160 12971
rect 15108 12928 15160 12937
rect 17132 12971 17184 12980
rect 17132 12937 17141 12971
rect 17141 12937 17175 12971
rect 17175 12937 17184 12971
rect 17132 12928 17184 12937
rect 17592 12971 17644 12980
rect 17592 12937 17601 12971
rect 17601 12937 17635 12971
rect 17635 12937 17644 12971
rect 17592 12928 17644 12937
rect 18972 12971 19024 12980
rect 18972 12937 18981 12971
rect 18981 12937 19015 12971
rect 19015 12937 19024 12971
rect 18972 12928 19024 12937
rect 21180 12928 21232 12980
rect 21640 12928 21692 12980
rect 24492 12928 24544 12980
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 25780 12928 25832 12980
rect 27620 12971 27672 12980
rect 15660 12860 15712 12912
rect 17684 12860 17736 12912
rect 18604 12860 18656 12912
rect 20904 12860 20956 12912
rect 22008 12860 22060 12912
rect 24032 12903 24084 12912
rect 24032 12869 24041 12903
rect 24041 12869 24075 12903
rect 24075 12869 24084 12903
rect 24032 12860 24084 12869
rect 24952 12860 25004 12912
rect 13268 12835 13320 12844
rect 13268 12801 13277 12835
rect 13277 12801 13311 12835
rect 13311 12801 13320 12835
rect 13268 12792 13320 12801
rect 14648 12792 14700 12844
rect 14464 12767 14516 12776
rect 12348 12699 12400 12708
rect 6644 12588 6696 12640
rect 12348 12665 12357 12699
rect 12357 12665 12391 12699
rect 12391 12665 12400 12699
rect 12348 12656 12400 12665
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 14556 12656 14608 12708
rect 10600 12588 10652 12640
rect 11244 12588 11296 12640
rect 12992 12588 13044 12640
rect 14280 12588 14332 12640
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 15476 12792 15528 12844
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 18236 12835 18288 12844
rect 18236 12801 18245 12835
rect 18245 12801 18279 12835
rect 18279 12801 18288 12835
rect 18236 12792 18288 12801
rect 18420 12792 18472 12844
rect 18972 12792 19024 12844
rect 20536 12792 20588 12844
rect 22284 12792 22336 12844
rect 18328 12724 18380 12776
rect 15292 12656 15344 12708
rect 14372 12588 14424 12597
rect 15384 12588 15436 12640
rect 22192 12724 22244 12776
rect 22744 12724 22796 12776
rect 22652 12631 22704 12640
rect 22652 12597 22661 12631
rect 22661 12597 22695 12631
rect 22695 12597 22704 12631
rect 22652 12588 22704 12597
rect 23112 12588 23164 12640
rect 25044 12835 25096 12844
rect 24032 12724 24084 12776
rect 23940 12656 23992 12708
rect 25044 12801 25053 12835
rect 25053 12801 25087 12835
rect 25087 12801 25096 12835
rect 25044 12792 25096 12801
rect 24952 12724 25004 12776
rect 25432 12835 25484 12844
rect 25432 12801 25467 12835
rect 25467 12801 25484 12835
rect 25432 12792 25484 12801
rect 27620 12937 27629 12971
rect 27629 12937 27663 12971
rect 27663 12937 27672 12971
rect 27620 12928 27672 12937
rect 31852 12928 31904 12980
rect 37464 12928 37516 12980
rect 30380 12860 30432 12912
rect 26976 12835 27028 12844
rect 26976 12801 26985 12835
rect 26985 12801 27019 12835
rect 27019 12801 27028 12835
rect 26976 12792 27028 12801
rect 27160 12835 27212 12844
rect 27160 12801 27164 12835
rect 27164 12801 27198 12835
rect 27198 12801 27212 12835
rect 27160 12792 27212 12801
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 28632 12792 28684 12844
rect 30288 12792 30340 12844
rect 32312 12835 32364 12844
rect 27528 12724 27580 12776
rect 29644 12767 29696 12776
rect 29644 12733 29653 12767
rect 29653 12733 29687 12767
rect 29687 12733 29696 12767
rect 29644 12724 29696 12733
rect 24676 12656 24728 12708
rect 26148 12656 26200 12708
rect 31760 12656 31812 12708
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 31944 12724 31996 12776
rect 32772 12656 32824 12708
rect 29092 12631 29144 12640
rect 29092 12597 29101 12631
rect 29101 12597 29135 12631
rect 29135 12597 29144 12631
rect 29092 12588 29144 12597
rect 30380 12588 30432 12640
rect 31392 12588 31444 12640
rect 34244 12860 34296 12912
rect 34336 12792 34388 12844
rect 35440 12792 35492 12844
rect 37096 12792 37148 12844
rect 40500 12792 40552 12844
rect 34244 12767 34296 12776
rect 34244 12733 34253 12767
rect 34253 12733 34287 12767
rect 34287 12733 34296 12767
rect 34244 12724 34296 12733
rect 33048 12656 33100 12708
rect 37372 12656 37424 12708
rect 38844 12699 38896 12708
rect 38844 12665 38853 12699
rect 38853 12665 38887 12699
rect 38887 12665 38896 12699
rect 38844 12656 38896 12665
rect 37464 12631 37516 12640
rect 37464 12597 37473 12631
rect 37473 12597 37507 12631
rect 37507 12597 37516 12631
rect 37464 12588 37516 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 1400 12180 1452 12232
rect 2780 12316 2832 12368
rect 3792 12248 3844 12300
rect 3976 12291 4028 12300
rect 3976 12257 3985 12291
rect 3985 12257 4019 12291
rect 4019 12257 4028 12291
rect 3976 12248 4028 12257
rect 2412 12112 2464 12164
rect 3240 12180 3292 12232
rect 2228 12044 2280 12096
rect 2596 12044 2648 12096
rect 3056 12112 3108 12164
rect 4712 12044 4764 12096
rect 8208 12384 8260 12436
rect 7932 12359 7984 12368
rect 7932 12325 7941 12359
rect 7941 12325 7975 12359
rect 7975 12325 7984 12359
rect 7932 12316 7984 12325
rect 9588 12316 9640 12368
rect 11520 12384 11572 12436
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 13544 12384 13596 12436
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 6644 12180 6696 12232
rect 7840 12112 7892 12164
rect 7472 12044 7524 12096
rect 9864 12112 9916 12164
rect 14096 12316 14148 12368
rect 15660 12384 15712 12436
rect 13084 12291 13136 12300
rect 13084 12257 13093 12291
rect 13093 12257 13127 12291
rect 13127 12257 13136 12291
rect 13084 12248 13136 12257
rect 14188 12248 14240 12300
rect 10784 12180 10836 12232
rect 10968 12180 11020 12232
rect 11888 12180 11940 12232
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 17868 12316 17920 12368
rect 19248 12316 19300 12368
rect 20260 12316 20312 12368
rect 11612 12112 11664 12164
rect 17408 12180 17460 12232
rect 17500 12180 17552 12232
rect 18236 12248 18288 12300
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 12440 12044 12492 12096
rect 12900 12044 12952 12096
rect 15476 12044 15528 12096
rect 16028 12112 16080 12164
rect 19248 12180 19300 12232
rect 18972 12112 19024 12164
rect 20079 12223 20131 12232
rect 20079 12189 20104 12223
rect 20104 12189 20131 12223
rect 20079 12180 20131 12189
rect 24676 12384 24728 12436
rect 26608 12384 26660 12436
rect 27528 12384 27580 12436
rect 28448 12384 28500 12436
rect 28908 12384 28960 12436
rect 29828 12427 29880 12436
rect 29828 12393 29837 12427
rect 29837 12393 29871 12427
rect 29871 12393 29880 12427
rect 29828 12384 29880 12393
rect 30288 12427 30340 12436
rect 30288 12393 30297 12427
rect 30297 12393 30331 12427
rect 30331 12393 30340 12427
rect 30288 12384 30340 12393
rect 33600 12384 33652 12436
rect 24032 12316 24084 12368
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 22652 12248 22704 12300
rect 25044 12248 25096 12300
rect 26976 12248 27028 12300
rect 17868 12044 17920 12096
rect 18052 12044 18104 12096
rect 19064 12044 19116 12096
rect 19432 12044 19484 12096
rect 22192 12180 22244 12232
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 24584 12180 24636 12232
rect 24768 12180 24820 12232
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 24032 12112 24084 12164
rect 28632 12223 28684 12232
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 28908 12248 28960 12300
rect 32404 12316 32456 12368
rect 32956 12359 33008 12368
rect 32956 12325 32965 12359
rect 32965 12325 32999 12359
rect 32999 12325 33008 12359
rect 32956 12316 33008 12325
rect 33140 12316 33192 12368
rect 32680 12248 32732 12300
rect 34520 12316 34572 12368
rect 28816 12223 28868 12232
rect 28816 12189 28825 12223
rect 28825 12189 28859 12223
rect 28859 12189 28868 12223
rect 28816 12180 28868 12189
rect 29644 12180 29696 12232
rect 31116 12180 31168 12232
rect 33416 12180 33468 12232
rect 28540 12112 28592 12164
rect 34244 12180 34296 12232
rect 35348 12384 35400 12436
rect 37464 12384 37516 12436
rect 39120 12384 39172 12436
rect 35716 12359 35768 12368
rect 35716 12325 35725 12359
rect 35725 12325 35759 12359
rect 35759 12325 35768 12359
rect 35716 12316 35768 12325
rect 34336 12112 34388 12164
rect 35900 12180 35952 12232
rect 37096 12223 37148 12232
rect 37096 12189 37105 12223
rect 37105 12189 37139 12223
rect 37139 12189 37148 12223
rect 37096 12180 37148 12189
rect 37464 12180 37516 12232
rect 39028 12180 39080 12232
rect 40408 12223 40460 12232
rect 40408 12189 40417 12223
rect 40417 12189 40451 12223
rect 40451 12189 40460 12223
rect 40408 12180 40460 12189
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 23112 12044 23164 12096
rect 23756 12044 23808 12096
rect 26516 12087 26568 12096
rect 26516 12053 26525 12087
rect 26525 12053 26559 12087
rect 26559 12053 26568 12087
rect 26516 12044 26568 12053
rect 26608 12044 26660 12096
rect 31024 12044 31076 12096
rect 32956 12044 33008 12096
rect 40684 12155 40736 12164
rect 40684 12121 40693 12155
rect 40693 12121 40727 12155
rect 40727 12121 40736 12155
rect 40684 12112 40736 12121
rect 34612 12044 34664 12096
rect 40224 12044 40276 12096
rect 40316 12044 40368 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2412 11840 2464 11892
rect 3240 11840 3292 11892
rect 5356 11840 5408 11892
rect 7196 11840 7248 11892
rect 7472 11840 7524 11892
rect 1768 11704 1820 11756
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 2596 11772 2648 11824
rect 2688 11704 2740 11756
rect 9312 11815 9364 11824
rect 9312 11781 9321 11815
rect 9321 11781 9355 11815
rect 9355 11781 9364 11815
rect 9312 11772 9364 11781
rect 9588 11772 9640 11824
rect 5816 11704 5868 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 9128 11704 9180 11756
rect 9680 11704 9732 11756
rect 2872 11636 2924 11688
rect 3148 11636 3200 11688
rect 9312 11636 9364 11688
rect 11520 11772 11572 11824
rect 11704 11772 11756 11824
rect 13636 11840 13688 11892
rect 14556 11840 14608 11892
rect 18144 11840 18196 11892
rect 18972 11840 19024 11892
rect 23388 11840 23440 11892
rect 24584 11883 24636 11892
rect 15752 11772 15804 11824
rect 17592 11772 17644 11824
rect 19708 11772 19760 11824
rect 23572 11772 23624 11824
rect 24584 11849 24593 11883
rect 24593 11849 24627 11883
rect 24627 11849 24636 11883
rect 24584 11840 24636 11849
rect 25504 11883 25556 11892
rect 25504 11849 25513 11883
rect 25513 11849 25547 11883
rect 25547 11849 25556 11883
rect 25504 11840 25556 11849
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 3056 11568 3108 11620
rect 9220 11568 9272 11620
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 6920 11500 6972 11509
rect 7932 11500 7984 11552
rect 9128 11500 9180 11552
rect 9680 11568 9732 11620
rect 10968 11704 11020 11756
rect 11336 11704 11388 11756
rect 11888 11636 11940 11688
rect 13360 11704 13412 11756
rect 14188 11704 14240 11756
rect 14556 11704 14608 11756
rect 17868 11747 17920 11756
rect 17868 11713 17877 11747
rect 17877 11713 17911 11747
rect 17911 11713 17920 11747
rect 17868 11704 17920 11713
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 19248 11704 19300 11756
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 20076 11747 20128 11756
rect 20076 11713 20085 11747
rect 20085 11713 20119 11747
rect 20119 11713 20128 11747
rect 20076 11704 20128 11713
rect 20260 11704 20312 11756
rect 20628 11704 20680 11756
rect 21088 11747 21140 11756
rect 21088 11713 21097 11747
rect 21097 11713 21131 11747
rect 21131 11713 21140 11747
rect 21088 11704 21140 11713
rect 24952 11772 25004 11824
rect 27252 11840 27304 11892
rect 27436 11840 27488 11892
rect 30656 11883 30708 11892
rect 30656 11849 30665 11883
rect 30665 11849 30699 11883
rect 30699 11849 30708 11883
rect 30656 11840 30708 11849
rect 26516 11772 26568 11824
rect 12440 11636 12492 11688
rect 17500 11636 17552 11688
rect 19524 11636 19576 11688
rect 21916 11636 21968 11688
rect 23940 11747 23992 11756
rect 23940 11713 23949 11747
rect 23949 11713 23983 11747
rect 23983 11713 23992 11747
rect 23940 11704 23992 11713
rect 24676 11704 24728 11756
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 25964 11747 26016 11756
rect 25964 11713 25973 11747
rect 25973 11713 26007 11747
rect 26007 11713 26016 11747
rect 25964 11704 26016 11713
rect 26976 11747 27028 11756
rect 26976 11713 26985 11747
rect 26985 11713 27019 11747
rect 27019 11713 27028 11747
rect 26976 11704 27028 11713
rect 28540 11772 28592 11824
rect 27528 11704 27580 11756
rect 28448 11747 28500 11756
rect 28448 11713 28457 11747
rect 28457 11713 28491 11747
rect 28491 11713 28500 11747
rect 28448 11704 28500 11713
rect 28632 11747 28684 11756
rect 28632 11713 28641 11747
rect 28641 11713 28675 11747
rect 28675 11713 28684 11747
rect 28632 11704 28684 11713
rect 28816 11747 28868 11756
rect 28816 11713 28825 11747
rect 28825 11713 28859 11747
rect 28859 11713 28868 11747
rect 28816 11704 28868 11713
rect 23020 11679 23072 11688
rect 23020 11645 23029 11679
rect 23029 11645 23063 11679
rect 23063 11645 23072 11679
rect 24860 11679 24912 11688
rect 23020 11636 23072 11645
rect 24860 11645 24869 11679
rect 24869 11645 24903 11679
rect 24903 11645 24912 11679
rect 24860 11636 24912 11645
rect 25780 11679 25832 11688
rect 25780 11645 25789 11679
rect 25789 11645 25823 11679
rect 25823 11645 25832 11679
rect 25780 11636 25832 11645
rect 9588 11543 9640 11552
rect 9588 11509 9597 11543
rect 9597 11509 9631 11543
rect 9631 11509 9640 11543
rect 9588 11500 9640 11509
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 19800 11568 19852 11620
rect 18328 11500 18380 11552
rect 20076 11500 20128 11552
rect 20444 11543 20496 11552
rect 20444 11509 20453 11543
rect 20453 11509 20487 11543
rect 20487 11509 20496 11543
rect 20444 11500 20496 11509
rect 20536 11500 20588 11552
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 26608 11636 26660 11688
rect 30840 11772 30892 11824
rect 29000 11704 29052 11756
rect 31300 11704 31352 11756
rect 33140 11840 33192 11892
rect 34336 11840 34388 11892
rect 35440 11840 35492 11892
rect 33048 11772 33100 11824
rect 33600 11815 33652 11824
rect 33600 11781 33609 11815
rect 33609 11781 33643 11815
rect 33643 11781 33652 11815
rect 33600 11772 33652 11781
rect 34520 11772 34572 11824
rect 33416 11747 33468 11756
rect 33416 11713 33425 11747
rect 33425 11713 33459 11747
rect 33459 11713 33468 11747
rect 33416 11704 33468 11713
rect 34244 11704 34296 11756
rect 35716 11772 35768 11824
rect 30656 11636 30708 11688
rect 35072 11747 35124 11756
rect 35072 11713 35081 11747
rect 35081 11713 35115 11747
rect 35115 11713 35124 11747
rect 39028 11840 39080 11892
rect 40224 11883 40276 11892
rect 40224 11849 40233 11883
rect 40233 11849 40267 11883
rect 40267 11849 40276 11883
rect 40224 11840 40276 11849
rect 37096 11772 37148 11824
rect 35072 11704 35124 11713
rect 35440 11636 35492 11688
rect 36360 11704 36412 11756
rect 37280 11704 37332 11756
rect 39764 11772 39816 11824
rect 36452 11636 36504 11688
rect 39120 11704 39172 11756
rect 40684 11772 40736 11824
rect 27620 11543 27672 11552
rect 27620 11509 27629 11543
rect 27629 11509 27663 11543
rect 27663 11509 27672 11543
rect 27620 11500 27672 11509
rect 31392 11568 31444 11620
rect 34428 11568 34480 11620
rect 34152 11500 34204 11552
rect 36820 11500 36872 11552
rect 67640 11611 67692 11620
rect 67640 11577 67649 11611
rect 67649 11577 67683 11611
rect 67683 11577 67692 11611
rect 67640 11568 67692 11577
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 3976 11296 4028 11348
rect 6552 11296 6604 11348
rect 7012 11296 7064 11348
rect 7288 11296 7340 11348
rect 9680 11296 9732 11348
rect 10968 11296 11020 11348
rect 13176 11296 13228 11348
rect 13544 11296 13596 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 19984 11296 20036 11348
rect 20352 11296 20404 11348
rect 20720 11296 20772 11348
rect 5816 11228 5868 11280
rect 10324 11228 10376 11280
rect 15660 11228 15712 11280
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 7012 11160 7064 11212
rect 7196 11160 7248 11212
rect 5080 11092 5132 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 6920 11024 6972 11076
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 9772 11160 9824 11212
rect 8116 11092 8168 11101
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 8392 11024 8444 11076
rect 8760 11024 8812 11076
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 13268 11160 13320 11212
rect 16488 11203 16540 11212
rect 16488 11169 16497 11203
rect 16497 11169 16531 11203
rect 16531 11169 16540 11203
rect 16488 11160 16540 11169
rect 11060 11092 11112 11101
rect 9864 11024 9916 11076
rect 14280 11092 14332 11144
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 19432 11228 19484 11280
rect 24032 11296 24084 11348
rect 24216 11296 24268 11348
rect 25688 11296 25740 11348
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 19340 11160 19392 11212
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 18512 11092 18564 11144
rect 18972 11092 19024 11144
rect 23480 11228 23532 11280
rect 23848 11228 23900 11280
rect 13360 11067 13412 11076
rect 13360 11033 13369 11067
rect 13369 11033 13403 11067
rect 13403 11033 13412 11067
rect 13360 11024 13412 11033
rect 14832 11024 14884 11076
rect 19340 11024 19392 11076
rect 20536 11092 20588 11144
rect 20628 11135 20680 11144
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 23940 11160 23992 11212
rect 28540 11296 28592 11348
rect 29000 11339 29052 11348
rect 29000 11305 29009 11339
rect 29009 11305 29043 11339
rect 29043 11305 29052 11339
rect 29000 11296 29052 11305
rect 29920 11339 29972 11348
rect 29920 11305 29929 11339
rect 29929 11305 29963 11339
rect 29963 11305 29972 11339
rect 29920 11296 29972 11305
rect 31116 11339 31168 11348
rect 31116 11305 31125 11339
rect 31125 11305 31159 11339
rect 31159 11305 31168 11339
rect 31116 11296 31168 11305
rect 31300 11296 31352 11348
rect 35440 11296 35492 11348
rect 29644 11271 29696 11280
rect 29644 11237 29653 11271
rect 29653 11237 29687 11271
rect 29687 11237 29696 11271
rect 29644 11228 29696 11237
rect 31024 11228 31076 11280
rect 38936 11296 38988 11348
rect 37556 11271 37608 11280
rect 20628 11092 20680 11101
rect 20444 11024 20496 11076
rect 7564 10956 7616 11008
rect 10048 10956 10100 11008
rect 15936 10956 15988 11008
rect 18328 10956 18380 11008
rect 22376 10956 22428 11008
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 24216 11092 24268 11144
rect 24768 11092 24820 11144
rect 25320 11092 25372 11144
rect 27620 11092 27672 11144
rect 32128 11160 32180 11212
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 31208 11092 31260 11144
rect 31392 11135 31444 11144
rect 31392 11101 31401 11135
rect 31401 11101 31435 11135
rect 31435 11101 31444 11135
rect 31668 11135 31720 11144
rect 31392 11092 31444 11101
rect 31668 11101 31677 11135
rect 31677 11101 31711 11135
rect 31711 11101 31720 11135
rect 31668 11092 31720 11101
rect 32680 11135 32732 11144
rect 24032 11024 24084 11076
rect 24124 11024 24176 11076
rect 23940 10956 23992 11008
rect 31392 10956 31444 11008
rect 31576 11024 31628 11076
rect 32680 11101 32689 11135
rect 32689 11101 32723 11135
rect 32723 11101 32732 11135
rect 32680 11092 32732 11101
rect 33416 11092 33468 11144
rect 32496 11067 32548 11076
rect 32496 11033 32505 11067
rect 32505 11033 32539 11067
rect 32539 11033 32548 11067
rect 32496 11024 32548 11033
rect 34428 11092 34480 11144
rect 34704 11092 34756 11144
rect 37556 11237 37565 11271
rect 37565 11237 37599 11271
rect 37599 11237 37608 11271
rect 37556 11228 37608 11237
rect 39120 11160 39172 11212
rect 40408 11160 40460 11212
rect 37096 11135 37148 11144
rect 37096 11101 37105 11135
rect 37105 11101 37139 11135
rect 37139 11101 37148 11135
rect 37096 11092 37148 11101
rect 38844 11092 38896 11144
rect 40132 11135 40184 11144
rect 40132 11101 40141 11135
rect 40141 11101 40175 11135
rect 40175 11101 40184 11135
rect 40132 11092 40184 11101
rect 36728 11024 36780 11076
rect 36820 11067 36872 11076
rect 36820 11033 36838 11067
rect 36838 11033 36872 11067
rect 36820 11024 36872 11033
rect 40316 11135 40368 11144
rect 40316 11101 40325 11135
rect 40325 11101 40359 11135
rect 40359 11101 40368 11135
rect 40316 11092 40368 11101
rect 40500 11135 40552 11144
rect 40500 11101 40509 11135
rect 40509 11101 40543 11135
rect 40543 11101 40552 11135
rect 40500 11092 40552 11101
rect 35716 10956 35768 11008
rect 40224 10956 40276 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 1860 10752 1912 10804
rect 3148 10752 3200 10804
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 8116 10752 8168 10804
rect 9496 10752 9548 10804
rect 12532 10752 12584 10804
rect 18328 10752 18380 10804
rect 19524 10752 19576 10804
rect 20168 10752 20220 10804
rect 20628 10752 20680 10804
rect 1400 10727 1452 10736
rect 1400 10693 1409 10727
rect 1409 10693 1443 10727
rect 1443 10693 1452 10727
rect 1400 10684 1452 10693
rect 5264 10684 5316 10736
rect 6552 10684 6604 10736
rect 3148 10616 3200 10668
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4712 10659 4764 10668
rect 4712 10625 4746 10659
rect 4746 10625 4764 10659
rect 4712 10616 4764 10625
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 7012 10616 7064 10668
rect 8944 10684 8996 10736
rect 11704 10727 11756 10736
rect 11704 10693 11713 10727
rect 11713 10693 11747 10727
rect 11747 10693 11756 10727
rect 11704 10684 11756 10693
rect 13636 10684 13688 10736
rect 7564 10659 7616 10668
rect 7564 10625 7598 10659
rect 7598 10625 7616 10659
rect 7564 10616 7616 10625
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 11060 10616 11112 10668
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12440 10616 12492 10668
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 14188 10616 14240 10668
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 15936 10616 15988 10668
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 18236 10616 18288 10668
rect 18512 10616 18564 10668
rect 11336 10548 11388 10600
rect 15476 10548 15528 10600
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 23112 10684 23164 10736
rect 19524 10616 19576 10668
rect 19156 10548 19208 10600
rect 12072 10523 12124 10532
rect 12072 10489 12081 10523
rect 12081 10489 12115 10523
rect 12115 10489 12124 10523
rect 12072 10480 12124 10489
rect 12256 10480 12308 10532
rect 9036 10412 9088 10464
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 17040 10412 17092 10464
rect 19524 10480 19576 10532
rect 20076 10616 20128 10668
rect 20996 10616 21048 10668
rect 22376 10616 22428 10668
rect 23480 10752 23532 10804
rect 24676 10752 24728 10804
rect 27528 10752 27580 10804
rect 30012 10795 30064 10804
rect 30012 10761 30021 10795
rect 30021 10761 30055 10795
rect 30055 10761 30064 10795
rect 30012 10752 30064 10761
rect 30656 10752 30708 10804
rect 32128 10795 32180 10804
rect 26700 10684 26752 10736
rect 23756 10659 23808 10668
rect 23756 10625 23765 10659
rect 23765 10625 23799 10659
rect 23799 10625 23808 10659
rect 23756 10616 23808 10625
rect 23848 10616 23900 10668
rect 24676 10659 24728 10668
rect 24676 10625 24685 10659
rect 24685 10625 24719 10659
rect 24719 10625 24728 10659
rect 24676 10616 24728 10625
rect 24952 10659 25004 10668
rect 24952 10625 24961 10659
rect 24961 10625 24995 10659
rect 24995 10625 25004 10659
rect 24952 10616 25004 10625
rect 29552 10659 29604 10668
rect 29552 10625 29561 10659
rect 29561 10625 29595 10659
rect 29595 10625 29604 10659
rect 29552 10616 29604 10625
rect 32128 10761 32137 10795
rect 32137 10761 32171 10795
rect 32171 10761 32180 10795
rect 32128 10752 32180 10761
rect 31392 10727 31444 10736
rect 31392 10693 31401 10727
rect 31401 10693 31435 10727
rect 31435 10693 31444 10727
rect 32496 10727 32548 10736
rect 31392 10684 31444 10693
rect 32496 10693 32505 10727
rect 32505 10693 32539 10727
rect 32539 10693 32548 10727
rect 32496 10684 32548 10693
rect 31208 10659 31260 10668
rect 31208 10625 31217 10659
rect 31217 10625 31251 10659
rect 31251 10625 31260 10659
rect 31208 10616 31260 10625
rect 31300 10659 31352 10668
rect 31300 10625 31309 10659
rect 31309 10625 31343 10659
rect 31343 10625 31352 10659
rect 31300 10616 31352 10625
rect 32220 10616 32272 10668
rect 38660 10752 38712 10804
rect 40316 10752 40368 10804
rect 34336 10684 34388 10736
rect 34612 10684 34664 10736
rect 36360 10684 36412 10736
rect 37556 10684 37608 10736
rect 40132 10727 40184 10736
rect 40132 10693 40141 10727
rect 40141 10693 40175 10727
rect 40175 10693 40184 10727
rect 40132 10684 40184 10693
rect 33324 10659 33376 10668
rect 28448 10548 28500 10600
rect 29000 10548 29052 10600
rect 33324 10625 33333 10659
rect 33333 10625 33367 10659
rect 33367 10625 33376 10659
rect 33324 10616 33376 10625
rect 34152 10659 34204 10668
rect 34152 10625 34161 10659
rect 34161 10625 34195 10659
rect 34195 10625 34204 10659
rect 34152 10616 34204 10625
rect 34704 10616 34756 10668
rect 38936 10616 38988 10668
rect 39948 10616 40000 10668
rect 20812 10480 20864 10532
rect 20904 10480 20956 10532
rect 27620 10523 27672 10532
rect 27620 10489 27629 10523
rect 27629 10489 27663 10523
rect 27663 10489 27672 10523
rect 27620 10480 27672 10489
rect 31576 10480 31628 10532
rect 18144 10412 18196 10464
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 21088 10412 21140 10464
rect 24216 10412 24268 10464
rect 26700 10412 26752 10464
rect 30380 10412 30432 10464
rect 30656 10412 30708 10464
rect 36452 10548 36504 10600
rect 34428 10412 34480 10464
rect 36360 10412 36412 10464
rect 39764 10412 39816 10464
rect 67640 10455 67692 10464
rect 67640 10421 67649 10455
rect 67649 10421 67683 10455
rect 67683 10421 67692 10455
rect 67640 10412 67692 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 3148 10208 3200 10260
rect 7196 10208 7248 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 19432 10208 19484 10260
rect 20628 10251 20680 10260
rect 20628 10217 20637 10251
rect 20637 10217 20671 10251
rect 20671 10217 20680 10251
rect 20628 10208 20680 10217
rect 21824 10208 21876 10260
rect 29000 10251 29052 10260
rect 14096 10140 14148 10192
rect 29000 10217 29009 10251
rect 29009 10217 29043 10251
rect 29043 10217 29052 10251
rect 29000 10208 29052 10217
rect 29920 10208 29972 10260
rect 35716 10251 35768 10260
rect 35716 10217 35725 10251
rect 35725 10217 35759 10251
rect 35759 10217 35768 10251
rect 35716 10208 35768 10217
rect 1400 10004 1452 10056
rect 1860 10004 1912 10056
rect 2044 10004 2096 10056
rect 7012 10072 7064 10124
rect 8024 10072 8076 10124
rect 8944 10072 8996 10124
rect 5080 10004 5132 10056
rect 10048 10004 10100 10056
rect 8300 9936 8352 9988
rect 14280 10004 14332 10056
rect 15476 10047 15528 10056
rect 13452 9936 13504 9988
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 30564 10140 30616 10192
rect 31300 10140 31352 10192
rect 38292 10140 38344 10192
rect 40224 10140 40276 10192
rect 16396 10072 16448 10124
rect 17408 10072 17460 10124
rect 23940 10072 23992 10124
rect 24676 10115 24728 10124
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 27344 10115 27396 10124
rect 27344 10081 27353 10115
rect 27353 10081 27387 10115
rect 27387 10081 27396 10115
rect 27344 10072 27396 10081
rect 17040 10004 17092 10056
rect 17500 10047 17552 10056
rect 16120 9936 16172 9988
rect 17500 10013 17509 10047
rect 17509 10013 17543 10047
rect 17543 10013 17552 10047
rect 17500 10004 17552 10013
rect 19340 10004 19392 10056
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 21916 10004 21968 10056
rect 24032 10004 24084 10056
rect 25228 10004 25280 10056
rect 25688 10004 25740 10056
rect 26240 10047 26292 10056
rect 26240 10013 26249 10047
rect 26249 10013 26283 10047
rect 26283 10013 26292 10047
rect 26240 10004 26292 10013
rect 28356 10004 28408 10056
rect 28908 10072 28960 10124
rect 17960 9936 18012 9988
rect 21364 9936 21416 9988
rect 27252 9979 27304 9988
rect 2596 9868 2648 9920
rect 9588 9868 9640 9920
rect 13176 9868 13228 9920
rect 15016 9868 15068 9920
rect 18328 9868 18380 9920
rect 27252 9945 27261 9979
rect 27261 9945 27295 9979
rect 27295 9945 27304 9979
rect 27252 9936 27304 9945
rect 22560 9868 22612 9920
rect 23112 9868 23164 9920
rect 29460 10004 29512 10056
rect 29828 10047 29880 10056
rect 29828 10013 29837 10047
rect 29837 10013 29871 10047
rect 29871 10013 29880 10047
rect 29828 10004 29880 10013
rect 33140 10072 33192 10124
rect 31576 10004 31628 10056
rect 32312 10004 32364 10056
rect 37556 10004 37608 10056
rect 39764 10004 39816 10056
rect 40500 10047 40552 10056
rect 28632 9979 28684 9988
rect 28632 9945 28641 9979
rect 28641 9945 28675 9979
rect 28675 9945 28684 9979
rect 28632 9936 28684 9945
rect 29368 9936 29420 9988
rect 29736 9979 29788 9988
rect 29736 9945 29745 9979
rect 29745 9945 29779 9979
rect 29779 9945 29788 9979
rect 29736 9936 29788 9945
rect 34428 9936 34480 9988
rect 34888 9979 34940 9988
rect 34888 9945 34897 9979
rect 34897 9945 34931 9979
rect 34931 9945 34940 9979
rect 34888 9936 34940 9945
rect 35624 9979 35676 9988
rect 35624 9945 35633 9979
rect 35633 9945 35667 9979
rect 35667 9945 35676 9979
rect 35624 9936 35676 9945
rect 38936 9979 38988 9988
rect 38936 9945 38945 9979
rect 38945 9945 38979 9979
rect 38979 9945 38988 9979
rect 38936 9936 38988 9945
rect 40500 10013 40509 10047
rect 40509 10013 40543 10047
rect 40543 10013 40552 10047
rect 40500 10004 40552 10013
rect 29000 9868 29052 9920
rect 34796 9868 34848 9920
rect 39856 9911 39908 9920
rect 39856 9877 39865 9911
rect 39865 9877 39899 9911
rect 39899 9877 39908 9911
rect 39856 9868 39908 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 1400 9664 1452 9716
rect 2688 9664 2740 9716
rect 5264 9707 5316 9716
rect 5264 9673 5273 9707
rect 5273 9673 5307 9707
rect 5307 9673 5316 9707
rect 5264 9664 5316 9673
rect 11796 9664 11848 9716
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 19432 9664 19484 9716
rect 21916 9707 21968 9716
rect 21916 9673 21925 9707
rect 21925 9673 21959 9707
rect 21959 9673 21968 9707
rect 21916 9664 21968 9673
rect 1768 9596 1820 9648
rect 2044 9528 2096 9580
rect 7656 9596 7708 9648
rect 8760 9596 8812 9648
rect 3884 9571 3936 9580
rect 2596 9460 2648 9512
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 10876 9639 10928 9648
rect 10876 9605 10885 9639
rect 10885 9605 10919 9639
rect 10919 9605 10928 9639
rect 10876 9596 10928 9605
rect 11704 9639 11756 9648
rect 11704 9605 11713 9639
rect 11713 9605 11747 9639
rect 11747 9605 11756 9639
rect 11704 9596 11756 9605
rect 21456 9596 21508 9648
rect 22560 9596 22612 9648
rect 23664 9639 23716 9648
rect 23664 9605 23673 9639
rect 23673 9605 23707 9639
rect 23707 9605 23716 9639
rect 23664 9596 23716 9605
rect 9772 9528 9824 9580
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 11060 9528 11112 9580
rect 6828 9460 6880 9512
rect 4896 9392 4948 9444
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 12532 9528 12584 9580
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 13176 9528 13228 9580
rect 15016 9571 15068 9580
rect 15016 9537 15050 9571
rect 15050 9537 15068 9571
rect 15016 9528 15068 9537
rect 18328 9571 18380 9580
rect 18328 9537 18346 9571
rect 18346 9537 18380 9571
rect 18328 9528 18380 9537
rect 21088 9528 21140 9580
rect 21640 9528 21692 9580
rect 21732 9528 21784 9580
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 23756 9528 23808 9580
rect 28632 9596 28684 9648
rect 29736 9596 29788 9648
rect 27804 9571 27856 9580
rect 13544 9460 13596 9512
rect 14280 9460 14332 9512
rect 18604 9503 18656 9512
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 25504 9503 25556 9512
rect 25504 9469 25513 9503
rect 25513 9469 25547 9503
rect 25547 9469 25556 9503
rect 25504 9460 25556 9469
rect 27804 9537 27813 9571
rect 27813 9537 27847 9571
rect 27847 9537 27856 9571
rect 27804 9528 27856 9537
rect 27712 9460 27764 9512
rect 27988 9571 28040 9580
rect 27988 9537 27997 9571
rect 27997 9537 28031 9571
rect 28031 9537 28040 9571
rect 32404 9664 32456 9716
rect 32680 9664 32732 9716
rect 37556 9707 37608 9716
rect 37556 9673 37565 9707
rect 37565 9673 37599 9707
rect 37599 9673 37608 9707
rect 37556 9664 37608 9673
rect 39764 9707 39816 9716
rect 39764 9673 39773 9707
rect 39773 9673 39807 9707
rect 39807 9673 39816 9707
rect 39764 9664 39816 9673
rect 27988 9528 28040 9537
rect 28080 9460 28132 9512
rect 8852 9367 8904 9376
rect 8852 9333 8861 9367
rect 8861 9333 8895 9367
rect 8895 9333 8904 9367
rect 8852 9324 8904 9333
rect 9680 9324 9732 9376
rect 9956 9324 10008 9376
rect 10048 9324 10100 9376
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 16856 9324 16908 9376
rect 17224 9367 17276 9376
rect 17224 9333 17233 9367
rect 17233 9333 17267 9367
rect 17267 9333 17276 9367
rect 17224 9324 17276 9333
rect 27252 9392 27304 9444
rect 19892 9324 19944 9376
rect 20352 9324 20404 9376
rect 28264 9367 28316 9376
rect 28264 9333 28273 9367
rect 28273 9333 28307 9367
rect 28307 9333 28316 9367
rect 28264 9324 28316 9333
rect 33324 9528 33376 9580
rect 34060 9528 34112 9580
rect 34796 9596 34848 9648
rect 39856 9596 39908 9648
rect 31300 9503 31352 9512
rect 31300 9469 31309 9503
rect 31309 9469 31343 9503
rect 31343 9469 31352 9503
rect 31300 9460 31352 9469
rect 32588 9460 32640 9512
rect 34704 9528 34756 9580
rect 38844 9528 38896 9580
rect 35624 9460 35676 9512
rect 36728 9503 36780 9512
rect 36728 9469 36737 9503
rect 36737 9469 36771 9503
rect 36771 9469 36780 9503
rect 36728 9460 36780 9469
rect 34796 9324 34848 9376
rect 36360 9324 36412 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 11060 9120 11112 9172
rect 13728 9120 13780 9172
rect 15292 9120 15344 9172
rect 24860 9120 24912 9172
rect 27344 9120 27396 9172
rect 27804 9120 27856 9172
rect 28356 9120 28408 9172
rect 33692 9120 33744 9172
rect 34704 9163 34756 9172
rect 34704 9129 34713 9163
rect 34713 9129 34747 9163
rect 34747 9129 34756 9163
rect 34704 9120 34756 9129
rect 14372 9052 14424 9104
rect 21364 9052 21416 9104
rect 2044 8984 2096 9036
rect 2964 8984 3016 9036
rect 3240 8984 3292 9036
rect 3976 8984 4028 9036
rect 2688 8916 2740 8968
rect 3884 8916 3936 8968
rect 4896 8848 4948 8900
rect 5540 8916 5592 8968
rect 8760 8984 8812 9036
rect 8944 9027 8996 9036
rect 8944 8993 8953 9027
rect 8953 8993 8987 9027
rect 8987 8993 8996 9027
rect 8944 8984 8996 8993
rect 15200 8984 15252 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 16396 8984 16448 9036
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 8852 8916 8904 8968
rect 14464 8916 14516 8968
rect 3240 8780 3292 8832
rect 3332 8780 3384 8832
rect 9772 8848 9824 8900
rect 11244 8848 11296 8900
rect 17316 8916 17368 8968
rect 8208 8780 8260 8832
rect 9128 8780 9180 8832
rect 10876 8780 10928 8832
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 11888 8780 11940 8832
rect 16304 8848 16356 8900
rect 12992 8780 13044 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 15016 8780 15068 8832
rect 15384 8780 15436 8832
rect 15844 8823 15896 8832
rect 15844 8789 15853 8823
rect 15853 8789 15887 8823
rect 15887 8789 15896 8823
rect 15844 8780 15896 8789
rect 16028 8780 16080 8832
rect 18972 8848 19024 8900
rect 20168 8959 20220 8968
rect 20168 8925 20177 8959
rect 20177 8925 20211 8959
rect 20211 8925 20220 8959
rect 20168 8916 20220 8925
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 20904 8984 20956 9036
rect 20536 8959 20588 8968
rect 20536 8925 20545 8959
rect 20545 8925 20579 8959
rect 20579 8925 20588 8959
rect 22836 8984 22888 9036
rect 20536 8916 20588 8925
rect 21916 8916 21968 8968
rect 24492 8848 24544 8900
rect 20352 8780 20404 8832
rect 20812 8823 20864 8832
rect 20812 8789 20821 8823
rect 20821 8789 20855 8823
rect 20855 8789 20864 8823
rect 20812 8780 20864 8789
rect 24676 8959 24728 8968
rect 24676 8925 24685 8959
rect 24685 8925 24719 8959
rect 24719 8925 24728 8959
rect 24952 8959 25004 8968
rect 24676 8916 24728 8925
rect 24952 8925 24961 8959
rect 24961 8925 24995 8959
rect 24995 8925 25004 8959
rect 24952 8916 25004 8925
rect 25504 9052 25556 9104
rect 26608 9052 26660 9104
rect 27528 9052 27580 9104
rect 29552 9052 29604 9104
rect 27620 8984 27672 9036
rect 27804 8984 27856 9036
rect 28264 8984 28316 9036
rect 26240 8916 26292 8968
rect 29552 8959 29604 8968
rect 29552 8925 29561 8959
rect 29561 8925 29595 8959
rect 29595 8925 29604 8959
rect 29552 8916 29604 8925
rect 31300 8984 31352 9036
rect 31576 8959 31628 8968
rect 31576 8925 31585 8959
rect 31585 8925 31619 8959
rect 31619 8925 31628 8959
rect 31576 8916 31628 8925
rect 31944 8959 31996 8968
rect 31944 8925 31953 8959
rect 31953 8925 31987 8959
rect 31987 8925 31996 8959
rect 31944 8916 31996 8925
rect 32312 8916 32364 8968
rect 34796 8984 34848 9036
rect 33692 8916 33744 8968
rect 25688 8780 25740 8832
rect 27252 8848 27304 8900
rect 27620 8780 27672 8832
rect 31484 8848 31536 8900
rect 32772 8891 32824 8900
rect 32772 8857 32781 8891
rect 32781 8857 32815 8891
rect 32815 8857 32824 8891
rect 32772 8848 32824 8857
rect 29828 8780 29880 8832
rect 32496 8823 32548 8832
rect 32496 8789 32505 8823
rect 32505 8789 32539 8823
rect 32539 8789 32548 8823
rect 32496 8780 32548 8789
rect 32588 8780 32640 8832
rect 33968 8959 34020 8968
rect 33968 8925 33977 8959
rect 33977 8925 34011 8959
rect 34011 8925 34020 8959
rect 33968 8916 34020 8925
rect 34244 8916 34296 8968
rect 36728 8984 36780 9036
rect 68100 8959 68152 8968
rect 68100 8925 68109 8959
rect 68109 8925 68143 8959
rect 68143 8925 68152 8959
rect 68100 8916 68152 8925
rect 34612 8780 34664 8832
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4896 8576 4948 8628
rect 7748 8576 7800 8628
rect 8208 8576 8260 8628
rect 2044 8440 2096 8492
rect 3332 8508 3384 8560
rect 3148 8440 3200 8492
rect 3976 8508 4028 8560
rect 6828 8508 6880 8560
rect 7932 8508 7984 8560
rect 9588 8508 9640 8560
rect 7012 8440 7064 8492
rect 9680 8440 9732 8492
rect 10140 8508 10192 8560
rect 12532 8576 12584 8628
rect 14096 8576 14148 8628
rect 2596 8304 2648 8356
rect 5908 8304 5960 8356
rect 6184 8304 6236 8356
rect 9036 8347 9088 8356
rect 9036 8313 9045 8347
rect 9045 8313 9079 8347
rect 9079 8313 9088 8347
rect 9036 8304 9088 8313
rect 9220 8304 9272 8356
rect 10968 8304 11020 8356
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 14004 8483 14056 8492
rect 14004 8449 14022 8483
rect 14022 8449 14056 8483
rect 14004 8440 14056 8449
rect 14924 8576 14976 8628
rect 20260 8576 20312 8628
rect 21456 8576 21508 8628
rect 25780 8576 25832 8628
rect 29368 8619 29420 8628
rect 15844 8508 15896 8560
rect 20812 8508 20864 8560
rect 23848 8508 23900 8560
rect 24676 8508 24728 8560
rect 26424 8508 26476 8560
rect 29368 8585 29377 8619
rect 29377 8585 29411 8619
rect 29411 8585 29420 8619
rect 29368 8576 29420 8585
rect 29644 8576 29696 8628
rect 33968 8619 34020 8628
rect 33968 8585 33977 8619
rect 33977 8585 34011 8619
rect 34011 8585 34020 8619
rect 33968 8576 34020 8585
rect 34336 8576 34388 8628
rect 10600 8236 10652 8288
rect 11060 8236 11112 8288
rect 11152 8236 11204 8288
rect 12624 8372 12676 8424
rect 14280 8415 14332 8424
rect 14280 8381 14289 8415
rect 14289 8381 14323 8415
rect 14323 8381 14332 8415
rect 14280 8372 14332 8381
rect 14648 8372 14700 8424
rect 19156 8440 19208 8492
rect 21364 8440 21416 8492
rect 23940 8440 23992 8492
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 24768 8440 24820 8492
rect 25688 8440 25740 8492
rect 20168 8415 20220 8424
rect 13084 8236 13136 8288
rect 13636 8236 13688 8288
rect 16856 8304 16908 8356
rect 16948 8304 17000 8356
rect 17316 8304 17368 8356
rect 18696 8236 18748 8288
rect 20168 8381 20177 8415
rect 20177 8381 20211 8415
rect 20211 8381 20220 8415
rect 20168 8372 20220 8381
rect 25136 8372 25188 8424
rect 25504 8372 25556 8424
rect 26516 8440 26568 8492
rect 27252 8483 27304 8492
rect 27252 8449 27261 8483
rect 27261 8449 27295 8483
rect 27295 8449 27304 8483
rect 27252 8440 27304 8449
rect 27712 8440 27764 8492
rect 31576 8508 31628 8560
rect 28172 8372 28224 8424
rect 29092 8440 29144 8492
rect 24492 8304 24544 8356
rect 31760 8440 31812 8492
rect 32312 8483 32364 8492
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 30932 8372 30984 8424
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32772 8508 32824 8560
rect 35256 8508 35308 8560
rect 36360 8551 36412 8560
rect 36360 8517 36369 8551
rect 36369 8517 36403 8551
rect 36403 8517 36412 8551
rect 36360 8508 36412 8517
rect 32496 8440 32548 8449
rect 34152 8440 34204 8492
rect 35532 8483 35584 8492
rect 35532 8449 35541 8483
rect 35541 8449 35575 8483
rect 35575 8449 35584 8483
rect 35532 8440 35584 8449
rect 37280 8440 37332 8492
rect 38844 8440 38896 8492
rect 33968 8304 34020 8356
rect 25044 8236 25096 8288
rect 36268 8236 36320 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 3884 8032 3936 8084
rect 5540 7896 5592 7948
rect 2136 7760 2188 7812
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 2412 7692 2464 7744
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 5080 7692 5132 7744
rect 7380 7828 7432 7880
rect 10232 7828 10284 7880
rect 7840 7692 7892 7744
rect 8944 7692 8996 7744
rect 11888 7964 11940 8016
rect 14004 8032 14056 8084
rect 16764 8032 16816 8084
rect 14464 7964 14516 8016
rect 16304 7964 16356 8016
rect 17776 7964 17828 8016
rect 11060 7896 11112 7948
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 13084 7871 13136 7880
rect 10876 7760 10928 7812
rect 11152 7760 11204 7812
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 26056 8032 26108 8084
rect 26884 8032 26936 8084
rect 28540 8032 28592 8084
rect 29092 8032 29144 8084
rect 31024 8032 31076 8084
rect 33692 8032 33744 8084
rect 34520 8032 34572 8084
rect 35532 8032 35584 8084
rect 30472 7964 30524 8016
rect 20720 7896 20772 7948
rect 13544 7760 13596 7812
rect 14832 7760 14884 7812
rect 10784 7692 10836 7744
rect 12256 7692 12308 7744
rect 12532 7692 12584 7744
rect 14280 7692 14332 7744
rect 15660 7692 15712 7744
rect 17224 7692 17276 7744
rect 20168 7828 20220 7880
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 22008 7871 22060 7880
rect 21456 7828 21508 7837
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 22192 7871 22244 7880
rect 22192 7837 22201 7871
rect 22201 7837 22235 7871
rect 22235 7837 22244 7871
rect 22192 7828 22244 7837
rect 18420 7760 18472 7812
rect 17868 7692 17920 7744
rect 18236 7692 18288 7744
rect 24676 7735 24728 7744
rect 24676 7701 24685 7735
rect 24685 7701 24719 7735
rect 24719 7701 24728 7735
rect 24676 7692 24728 7701
rect 25136 7871 25188 7880
rect 25136 7837 25145 7871
rect 25145 7837 25179 7871
rect 25179 7837 25188 7871
rect 25136 7828 25188 7837
rect 25320 7871 25372 7880
rect 25320 7837 25329 7871
rect 25329 7837 25363 7871
rect 25363 7837 25372 7871
rect 26056 7871 26108 7880
rect 25320 7828 25372 7837
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 25228 7760 25280 7812
rect 26240 7871 26292 7880
rect 26240 7837 26249 7871
rect 26249 7837 26283 7871
rect 26283 7837 26292 7871
rect 27712 7896 27764 7948
rect 26240 7828 26292 7837
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 27988 7871 28040 7880
rect 27988 7837 27997 7871
rect 27997 7837 28031 7871
rect 28031 7837 28040 7871
rect 31024 7896 31076 7948
rect 27988 7828 28040 7837
rect 31668 7871 31720 7880
rect 31668 7837 31677 7871
rect 31677 7837 31711 7871
rect 31711 7837 31720 7871
rect 31668 7828 31720 7837
rect 32772 7896 32824 7948
rect 35624 7939 35676 7948
rect 34428 7828 34480 7880
rect 28080 7760 28132 7812
rect 25044 7692 25096 7744
rect 25688 7692 25740 7744
rect 28356 7692 28408 7744
rect 31852 7803 31904 7812
rect 31852 7769 31861 7803
rect 31861 7769 31895 7803
rect 31895 7769 31904 7803
rect 31852 7760 31904 7769
rect 32496 7760 32548 7812
rect 35624 7905 35633 7939
rect 35633 7905 35667 7939
rect 35667 7905 35676 7939
rect 35624 7896 35676 7905
rect 35900 7828 35952 7880
rect 36360 7964 36412 8016
rect 37280 8032 37332 8084
rect 40500 7964 40552 8016
rect 36268 7828 36320 7880
rect 68100 7871 68152 7880
rect 68100 7837 68109 7871
rect 68109 7837 68143 7871
rect 68143 7837 68152 7871
rect 68100 7828 68152 7837
rect 33232 7692 33284 7744
rect 36176 7692 36228 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 9312 7488 9364 7540
rect 10140 7488 10192 7540
rect 12900 7488 12952 7540
rect 14280 7488 14332 7540
rect 14832 7488 14884 7540
rect 18420 7488 18472 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 26240 7488 26292 7540
rect 27988 7488 28040 7540
rect 29092 7488 29144 7540
rect 36268 7488 36320 7540
rect 36360 7488 36412 7540
rect 8300 7420 8352 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 6460 7352 6512 7404
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 10600 7352 10652 7404
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 3056 7216 3108 7268
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 7196 7284 7248 7336
rect 23940 7463 23992 7472
rect 12532 7395 12584 7404
rect 12532 7361 12541 7395
rect 12541 7361 12575 7395
rect 12575 7361 12584 7395
rect 12532 7352 12584 7361
rect 13176 7352 13228 7404
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 14832 7352 14884 7404
rect 18236 7395 18288 7404
rect 18236 7361 18254 7395
rect 18254 7361 18288 7395
rect 18236 7352 18288 7361
rect 21272 7352 21324 7404
rect 23940 7429 23949 7463
rect 23949 7429 23983 7463
rect 23983 7429 23992 7463
rect 23940 7420 23992 7429
rect 26332 7420 26384 7472
rect 27620 7463 27672 7472
rect 27620 7429 27629 7463
rect 27629 7429 27663 7463
rect 27663 7429 27672 7463
rect 27620 7420 27672 7429
rect 31024 7420 31076 7472
rect 31944 7420 31996 7472
rect 32404 7420 32456 7472
rect 4620 7148 4672 7200
rect 15568 7216 15620 7268
rect 11520 7148 11572 7200
rect 16396 7148 16448 7200
rect 16764 7148 16816 7200
rect 17224 7148 17276 7200
rect 18604 7284 18656 7336
rect 18972 7284 19024 7336
rect 20720 7284 20772 7336
rect 22192 7352 22244 7404
rect 24860 7352 24912 7404
rect 26424 7352 26476 7404
rect 27252 7284 27304 7336
rect 31392 7352 31444 7404
rect 34520 7420 34572 7472
rect 34152 7352 34204 7404
rect 34612 7352 34664 7404
rect 35900 7395 35952 7404
rect 35900 7361 35909 7395
rect 35909 7361 35943 7395
rect 35943 7361 35952 7395
rect 35900 7352 35952 7361
rect 36084 7395 36136 7404
rect 36084 7361 36088 7395
rect 36088 7361 36122 7395
rect 36122 7361 36136 7395
rect 36084 7352 36136 7361
rect 31852 7216 31904 7268
rect 18788 7148 18840 7200
rect 20536 7148 20588 7200
rect 22744 7148 22796 7200
rect 24768 7148 24820 7200
rect 27804 7148 27856 7200
rect 28448 7148 28500 7200
rect 28540 7148 28592 7200
rect 30288 7191 30340 7200
rect 30288 7157 30297 7191
rect 30297 7157 30331 7191
rect 30331 7157 30340 7191
rect 30288 7148 30340 7157
rect 31024 7148 31076 7200
rect 32312 7148 32364 7200
rect 33508 7148 33560 7200
rect 36084 7216 36136 7268
rect 38844 7395 38896 7404
rect 38844 7361 38853 7395
rect 38853 7361 38887 7395
rect 38887 7361 38896 7395
rect 38844 7352 38896 7361
rect 39028 7395 39080 7404
rect 39028 7361 39037 7395
rect 39037 7361 39071 7395
rect 39071 7361 39080 7395
rect 39028 7352 39080 7361
rect 35624 7148 35676 7200
rect 36544 7191 36596 7200
rect 36544 7157 36553 7191
rect 36553 7157 36587 7191
rect 36587 7157 36596 7191
rect 36544 7148 36596 7157
rect 38384 7191 38436 7200
rect 38384 7157 38393 7191
rect 38393 7157 38427 7191
rect 38427 7157 38436 7191
rect 38384 7148 38436 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 4436 6944 4488 6996
rect 10048 6944 10100 6996
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 3240 6808 3292 6860
rect 5172 6808 5224 6860
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 10416 6876 10468 6928
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 9772 6808 9824 6860
rect 10232 6808 10284 6860
rect 4620 6740 4672 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 8208 6783 8260 6792
rect 5448 6740 5500 6749
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 9680 6740 9732 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 2504 6672 2556 6724
rect 1952 6604 2004 6656
rect 4712 6604 4764 6656
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 5540 6672 5592 6724
rect 6552 6604 6604 6656
rect 7472 6604 7524 6656
rect 8300 6604 8352 6656
rect 8484 6604 8536 6656
rect 9128 6604 9180 6656
rect 10968 6944 11020 6996
rect 12532 6944 12584 6996
rect 20260 6944 20312 6996
rect 23848 6987 23900 6996
rect 23848 6953 23857 6987
rect 23857 6953 23891 6987
rect 23891 6953 23900 6987
rect 23848 6944 23900 6953
rect 26424 6944 26476 6996
rect 31116 6944 31168 6996
rect 32404 6987 32456 6996
rect 32404 6953 32413 6987
rect 32413 6953 32447 6987
rect 32447 6953 32456 6987
rect 32404 6944 32456 6953
rect 38844 6944 38896 6996
rect 11336 6876 11388 6928
rect 12440 6876 12492 6928
rect 14832 6876 14884 6928
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11152 6808 11204 6860
rect 14280 6808 14332 6860
rect 15108 6876 15160 6928
rect 36268 6919 36320 6928
rect 36268 6885 36277 6919
rect 36277 6885 36311 6919
rect 36311 6885 36320 6919
rect 36268 6876 36320 6885
rect 17224 6851 17276 6860
rect 10968 6604 11020 6656
rect 11152 6604 11204 6656
rect 12624 6740 12676 6792
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 14464 6740 14516 6792
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 17224 6817 17233 6851
rect 17233 6817 17267 6851
rect 17267 6817 17276 6851
rect 17224 6808 17276 6817
rect 18604 6808 18656 6860
rect 35532 6808 35584 6860
rect 35992 6808 36044 6860
rect 11428 6647 11480 6656
rect 11428 6613 11437 6647
rect 11437 6613 11471 6647
rect 11471 6613 11480 6647
rect 11428 6604 11480 6613
rect 12716 6604 12768 6656
rect 14096 6604 14148 6656
rect 17592 6740 17644 6792
rect 18052 6740 18104 6792
rect 18236 6749 18245 6770
rect 18245 6749 18279 6770
rect 18279 6749 18288 6770
rect 18236 6718 18288 6749
rect 18512 6783 18564 6792
rect 16028 6604 16080 6656
rect 16304 6604 16356 6656
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 23480 6740 23532 6792
rect 23940 6740 23992 6792
rect 25688 6783 25740 6792
rect 25688 6749 25722 6783
rect 25722 6749 25740 6783
rect 25688 6740 25740 6749
rect 28356 6783 28408 6792
rect 28356 6749 28374 6783
rect 28374 6749 28408 6783
rect 28632 6783 28684 6792
rect 28356 6740 28408 6749
rect 28632 6749 28641 6783
rect 28641 6749 28675 6783
rect 28675 6749 28684 6783
rect 29552 6783 29604 6792
rect 28632 6740 28684 6749
rect 29552 6749 29561 6783
rect 29561 6749 29595 6783
rect 29595 6749 29604 6783
rect 29552 6740 29604 6749
rect 21640 6672 21692 6724
rect 24676 6672 24728 6724
rect 24768 6715 24820 6724
rect 24768 6681 24777 6715
rect 24777 6681 24811 6715
rect 24811 6681 24820 6715
rect 24768 6672 24820 6681
rect 25044 6672 25096 6724
rect 30748 6740 30800 6792
rect 30932 6740 30984 6792
rect 38660 6740 38712 6792
rect 30564 6672 30616 6724
rect 31392 6715 31444 6724
rect 31392 6681 31401 6715
rect 31401 6681 31435 6715
rect 31435 6681 31444 6715
rect 31392 6672 31444 6681
rect 31576 6715 31628 6724
rect 31576 6681 31585 6715
rect 31585 6681 31619 6715
rect 31619 6681 31628 6715
rect 31576 6672 31628 6681
rect 32956 6672 33008 6724
rect 18512 6604 18564 6656
rect 20812 6604 20864 6656
rect 27620 6604 27672 6656
rect 30472 6604 30524 6656
rect 31852 6604 31904 6656
rect 32220 6604 32272 6656
rect 36544 6672 36596 6724
rect 37280 6672 37332 6724
rect 38752 6715 38804 6724
rect 38752 6681 38761 6715
rect 38761 6681 38795 6715
rect 38795 6681 38804 6715
rect 38752 6672 38804 6681
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 2228 6400 2280 6452
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 3976 6400 4028 6452
rect 4804 6400 4856 6452
rect 3240 6332 3292 6384
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 5724 6264 5776 6316
rect 7564 6332 7616 6384
rect 9312 6400 9364 6452
rect 10048 6332 10100 6384
rect 6276 6264 6328 6316
rect 9128 6264 9180 6316
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 12256 6400 12308 6452
rect 14832 6400 14884 6452
rect 17776 6400 17828 6452
rect 20904 6400 20956 6452
rect 21364 6400 21416 6452
rect 24952 6400 25004 6452
rect 25688 6400 25740 6452
rect 26884 6400 26936 6452
rect 30564 6443 30616 6452
rect 30564 6409 30573 6443
rect 30573 6409 30607 6443
rect 30607 6409 30616 6443
rect 30564 6400 30616 6409
rect 32312 6400 32364 6452
rect 32956 6443 33008 6452
rect 11888 6332 11940 6384
rect 14096 6332 14148 6384
rect 18696 6332 18748 6384
rect 10416 6264 10468 6316
rect 11428 6264 11480 6316
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 14556 6264 14608 6316
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 4068 6196 4120 6248
rect 5448 6196 5500 6248
rect 5632 6196 5684 6248
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 4988 6128 5040 6180
rect 4436 6103 4488 6112
rect 4436 6069 4445 6103
rect 4445 6069 4479 6103
rect 4479 6069 4488 6103
rect 4436 6060 4488 6069
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 5724 6060 5776 6112
rect 8024 6128 8076 6180
rect 11060 6128 11112 6180
rect 6736 6060 6788 6112
rect 8300 6060 8352 6112
rect 10232 6060 10284 6112
rect 10416 6060 10468 6112
rect 11152 6060 11204 6112
rect 11980 6060 12032 6112
rect 13820 6196 13872 6248
rect 17868 6264 17920 6316
rect 17684 6239 17736 6248
rect 17684 6205 17693 6239
rect 17693 6205 17727 6239
rect 17727 6205 17736 6239
rect 17684 6196 17736 6205
rect 17776 6196 17828 6248
rect 20536 6332 20588 6384
rect 20260 6264 20312 6316
rect 20812 6313 20864 6316
rect 20812 6279 20816 6313
rect 20816 6279 20850 6313
rect 20850 6279 20864 6313
rect 20812 6264 20864 6279
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 23480 6264 23532 6316
rect 24492 6307 24544 6316
rect 24492 6273 24526 6307
rect 24526 6273 24544 6307
rect 24492 6264 24544 6273
rect 25412 6264 25464 6316
rect 20076 6239 20128 6248
rect 20076 6205 20085 6239
rect 20085 6205 20119 6239
rect 20119 6205 20128 6239
rect 20076 6196 20128 6205
rect 24216 6239 24268 6248
rect 24216 6205 24225 6239
rect 24225 6205 24259 6239
rect 24259 6205 24268 6239
rect 24216 6196 24268 6205
rect 26332 6264 26384 6316
rect 27988 6307 28040 6316
rect 27988 6273 27997 6307
rect 27997 6273 28031 6307
rect 28031 6273 28040 6307
rect 27988 6264 28040 6273
rect 30380 6264 30432 6316
rect 30840 6307 30892 6316
rect 30840 6273 30849 6307
rect 30849 6273 30883 6307
rect 30883 6273 30892 6307
rect 30840 6264 30892 6273
rect 17592 6128 17644 6180
rect 20260 6128 20312 6180
rect 28632 6128 28684 6180
rect 16488 6060 16540 6112
rect 17500 6060 17552 6112
rect 17776 6060 17828 6112
rect 18604 6060 18656 6112
rect 19432 6060 19484 6112
rect 31024 6307 31076 6316
rect 31024 6273 31033 6307
rect 31033 6273 31067 6307
rect 31067 6273 31076 6307
rect 31024 6264 31076 6273
rect 32956 6409 32965 6443
rect 32965 6409 32999 6443
rect 32999 6409 33008 6443
rect 32956 6400 33008 6409
rect 32772 6332 32824 6384
rect 33232 6332 33284 6384
rect 32680 6307 32732 6316
rect 32680 6273 32689 6307
rect 32689 6273 32723 6307
rect 32723 6273 32732 6307
rect 33508 6307 33560 6316
rect 32680 6264 32732 6273
rect 33508 6273 33517 6307
rect 33517 6273 33551 6307
rect 33551 6273 33560 6307
rect 33508 6264 33560 6273
rect 35624 6307 35676 6316
rect 35624 6273 35633 6307
rect 35633 6273 35667 6307
rect 35667 6273 35676 6307
rect 35624 6264 35676 6273
rect 35992 6264 36044 6316
rect 39028 6264 39080 6316
rect 37188 6196 37240 6248
rect 33140 6128 33192 6180
rect 34060 6128 34112 6180
rect 67640 6171 67692 6180
rect 67640 6137 67649 6171
rect 67649 6137 67683 6171
rect 67683 6137 67692 6171
rect 67640 6128 67692 6137
rect 31668 6060 31720 6112
rect 32772 6060 32824 6112
rect 34612 6060 34664 6112
rect 35532 6060 35584 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 4896 5856 4948 5908
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 8116 5856 8168 5908
rect 13728 5856 13780 5908
rect 15200 5856 15252 5908
rect 17960 5856 18012 5908
rect 18236 5856 18288 5908
rect 5448 5788 5500 5840
rect 1860 5720 1912 5772
rect 2320 5720 2372 5772
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 7932 5788 7984 5840
rect 8300 5788 8352 5840
rect 10876 5788 10928 5840
rect 11060 5788 11112 5840
rect 12532 5788 12584 5840
rect 12716 5831 12768 5840
rect 12716 5797 12725 5831
rect 12725 5797 12759 5831
rect 12759 5797 12768 5831
rect 12716 5788 12768 5797
rect 13544 5788 13596 5840
rect 9404 5720 9456 5772
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 11520 5720 11572 5772
rect 3148 5652 3200 5704
rect 5632 5652 5684 5704
rect 7104 5695 7156 5704
rect 2780 5584 2832 5636
rect 4160 5584 4212 5636
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 8668 5584 8720 5636
rect 1952 5516 2004 5568
rect 4068 5516 4120 5568
rect 5172 5516 5224 5568
rect 7012 5516 7064 5568
rect 8300 5516 8352 5568
rect 9312 5652 9364 5704
rect 14556 5763 14608 5772
rect 14556 5729 14565 5763
rect 14565 5729 14599 5763
rect 14599 5729 14608 5763
rect 14556 5720 14608 5729
rect 13268 5652 13320 5704
rect 14096 5695 14148 5704
rect 9128 5584 9180 5636
rect 10692 5516 10744 5568
rect 11612 5584 11664 5636
rect 12072 5584 12124 5636
rect 13176 5584 13228 5636
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 18328 5788 18380 5840
rect 19156 5788 19208 5840
rect 23664 5856 23716 5908
rect 24492 5856 24544 5908
rect 26332 5899 26384 5908
rect 26332 5865 26341 5899
rect 26341 5865 26375 5899
rect 26375 5865 26384 5899
rect 26332 5856 26384 5865
rect 26700 5856 26752 5908
rect 27344 5856 27396 5908
rect 27896 5856 27948 5908
rect 29460 5856 29512 5908
rect 30748 5856 30800 5908
rect 17132 5720 17184 5772
rect 17684 5720 17736 5772
rect 20076 5720 20128 5772
rect 24216 5788 24268 5840
rect 28356 5788 28408 5840
rect 28632 5788 28684 5840
rect 20904 5720 20956 5772
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 18052 5652 18104 5704
rect 19340 5652 19392 5704
rect 21640 5695 21692 5704
rect 15292 5584 15344 5636
rect 16304 5584 16356 5636
rect 16856 5584 16908 5636
rect 18696 5627 18748 5636
rect 18696 5593 18705 5627
rect 18705 5593 18739 5627
rect 18739 5593 18748 5627
rect 18696 5584 18748 5593
rect 20260 5584 20312 5636
rect 21640 5661 21649 5695
rect 21649 5661 21683 5695
rect 21683 5661 21692 5695
rect 21640 5652 21692 5661
rect 24584 5652 24636 5704
rect 25596 5720 25648 5772
rect 27896 5720 27948 5772
rect 30932 5763 30984 5772
rect 25136 5652 25188 5704
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 28172 5695 28224 5704
rect 28172 5661 28176 5695
rect 28176 5661 28210 5695
rect 28210 5661 28224 5695
rect 28172 5652 28224 5661
rect 30932 5729 30941 5763
rect 30941 5729 30975 5763
rect 30975 5729 30984 5763
rect 30932 5720 30984 5729
rect 31852 5695 31904 5704
rect 31852 5661 31866 5695
rect 31866 5661 31900 5695
rect 31900 5661 31904 5695
rect 31852 5652 31904 5661
rect 33140 5652 33192 5704
rect 38660 5856 38712 5908
rect 35624 5720 35676 5772
rect 34060 5652 34112 5704
rect 34244 5652 34296 5704
rect 25872 5627 25924 5636
rect 25872 5593 25881 5627
rect 25881 5593 25915 5627
rect 25915 5593 25924 5627
rect 25872 5584 25924 5593
rect 26976 5584 27028 5636
rect 27896 5584 27948 5636
rect 38384 5652 38436 5704
rect 35072 5627 35124 5636
rect 35072 5593 35081 5627
rect 35081 5593 35115 5627
rect 35115 5593 35124 5627
rect 35072 5584 35124 5593
rect 35348 5584 35400 5636
rect 37280 5584 37332 5636
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 16672 5516 16724 5568
rect 19984 5516 20036 5568
rect 20076 5516 20128 5568
rect 20812 5516 20864 5568
rect 23020 5516 23072 5568
rect 27252 5516 27304 5568
rect 28264 5516 28316 5568
rect 31300 5516 31352 5568
rect 31668 5516 31720 5568
rect 34520 5516 34572 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4160 5312 4212 5364
rect 4988 5312 5040 5364
rect 5540 5312 5592 5364
rect 8668 5355 8720 5364
rect 8668 5321 8677 5355
rect 8677 5321 8711 5355
rect 8711 5321 8720 5355
rect 8668 5312 8720 5321
rect 9036 5355 9088 5364
rect 9036 5321 9045 5355
rect 9045 5321 9079 5355
rect 9079 5321 9088 5355
rect 9036 5312 9088 5321
rect 9312 5312 9364 5364
rect 14924 5312 14976 5364
rect 15016 5312 15068 5364
rect 16304 5312 16356 5364
rect 19340 5312 19392 5364
rect 23020 5312 23072 5364
rect 10876 5244 10928 5296
rect 11520 5287 11572 5296
rect 11520 5253 11529 5287
rect 11529 5253 11563 5287
rect 11563 5253 11572 5287
rect 11520 5244 11572 5253
rect 11612 5244 11664 5296
rect 12348 5244 12400 5296
rect 13544 5244 13596 5296
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 5448 5176 5500 5228
rect 5816 5176 5868 5228
rect 6368 5176 6420 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 8024 5176 8076 5228
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 9772 5176 9824 5228
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 4804 5151 4856 5160
rect 4804 5117 4813 5151
rect 4813 5117 4847 5151
rect 4847 5117 4856 5151
rect 4804 5108 4856 5117
rect 9312 5151 9364 5160
rect 8852 5040 8904 5092
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 7380 4972 7432 5024
rect 7472 4972 7524 5024
rect 8944 4972 8996 5024
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 10048 5108 10100 5160
rect 12900 5176 12952 5228
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 15384 5244 15436 5296
rect 17132 5287 17184 5296
rect 17132 5253 17141 5287
rect 17141 5253 17175 5287
rect 17175 5253 17184 5287
rect 17132 5244 17184 5253
rect 20444 5244 20496 5296
rect 24768 5312 24820 5364
rect 25596 5312 25648 5364
rect 27252 5312 27304 5364
rect 27988 5312 28040 5364
rect 34796 5312 34848 5364
rect 35072 5312 35124 5364
rect 37188 5312 37240 5364
rect 12808 5108 12860 5160
rect 13176 5108 13228 5160
rect 13544 5108 13596 5160
rect 15016 5176 15068 5228
rect 16580 5176 16632 5228
rect 19248 5176 19300 5228
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 20076 5176 20128 5228
rect 21180 5176 21232 5228
rect 23480 5176 23532 5228
rect 23664 5219 23716 5228
rect 23664 5185 23673 5219
rect 23673 5185 23707 5219
rect 23707 5185 23716 5219
rect 23664 5176 23716 5185
rect 10232 4972 10284 5024
rect 11612 5015 11664 5024
rect 11612 4981 11621 5015
rect 11621 4981 11655 5015
rect 11655 4981 11664 5015
rect 11612 4972 11664 4981
rect 11980 4972 12032 5024
rect 12348 5040 12400 5092
rect 16856 5108 16908 5160
rect 19156 5108 19208 5160
rect 14648 5040 14700 5092
rect 14740 4972 14792 5024
rect 15200 5040 15252 5092
rect 15292 5040 15344 5092
rect 17776 5040 17828 5092
rect 20536 5108 20588 5160
rect 25872 5244 25924 5296
rect 26608 5244 26660 5296
rect 25136 5176 25188 5228
rect 26976 5219 27028 5228
rect 26976 5185 26985 5219
rect 26985 5185 27019 5219
rect 27019 5185 27028 5219
rect 26976 5176 27028 5185
rect 29460 5244 29512 5296
rect 30932 5244 30984 5296
rect 32680 5244 32732 5296
rect 33508 5244 33560 5296
rect 33968 5287 34020 5296
rect 27344 5219 27396 5228
rect 27344 5185 27353 5219
rect 27353 5185 27387 5219
rect 27387 5185 27396 5219
rect 28080 5219 28132 5228
rect 27344 5176 27396 5185
rect 28080 5185 28089 5219
rect 28089 5185 28123 5219
rect 28123 5185 28132 5219
rect 28080 5176 28132 5185
rect 28172 5176 28224 5228
rect 31300 5219 31352 5228
rect 31300 5185 31318 5219
rect 31318 5185 31352 5219
rect 31576 5219 31628 5228
rect 31300 5176 31352 5185
rect 31576 5185 31585 5219
rect 31585 5185 31619 5219
rect 31619 5185 31628 5219
rect 31576 5176 31628 5185
rect 17684 4972 17736 5024
rect 28724 5040 28776 5092
rect 30472 5040 30524 5092
rect 33968 5253 33977 5287
rect 33977 5253 34011 5287
rect 34011 5253 34020 5287
rect 33968 5244 34020 5253
rect 34060 5244 34112 5296
rect 34612 5244 34664 5296
rect 34244 5176 34296 5228
rect 35624 5244 35676 5296
rect 35992 5219 36044 5228
rect 34060 5108 34112 5160
rect 35992 5185 36001 5219
rect 36001 5185 36035 5219
rect 36035 5185 36044 5219
rect 35992 5176 36044 5185
rect 38292 5287 38344 5296
rect 38292 5253 38301 5287
rect 38301 5253 38335 5287
rect 38335 5253 38344 5287
rect 38292 5244 38344 5253
rect 35624 5108 35676 5160
rect 36360 5219 36412 5228
rect 36360 5185 36369 5219
rect 36369 5185 36403 5219
rect 36403 5185 36412 5219
rect 36360 5176 36412 5185
rect 36820 5176 36872 5228
rect 38752 5176 38804 5228
rect 58808 5108 58860 5160
rect 59268 5040 59320 5092
rect 19432 4972 19484 5024
rect 19984 4972 20036 5024
rect 20352 4972 20404 5024
rect 20904 4972 20956 5024
rect 27344 4972 27396 5024
rect 27620 5015 27672 5024
rect 27620 4981 27629 5015
rect 27629 4981 27663 5015
rect 27663 4981 27672 5015
rect 27620 4972 27672 4981
rect 35348 5015 35400 5024
rect 35348 4981 35357 5015
rect 35357 4981 35391 5015
rect 35391 4981 35400 5015
rect 35348 4972 35400 4981
rect 36636 5015 36688 5024
rect 36636 4981 36645 5015
rect 36645 4981 36679 5015
rect 36679 4981 36688 5015
rect 36636 4972 36688 4981
rect 58716 4972 58768 5024
rect 67640 5015 67692 5024
rect 67640 4981 67649 5015
rect 67649 4981 67683 5015
rect 67683 4981 67692 5015
rect 67640 4972 67692 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 9956 4768 10008 4820
rect 10416 4811 10468 4820
rect 10416 4777 10425 4811
rect 10425 4777 10459 4811
rect 10459 4777 10468 4811
rect 10416 4768 10468 4777
rect 12900 4768 12952 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 21180 4811 21232 4820
rect 21180 4777 21189 4811
rect 21189 4777 21223 4811
rect 21223 4777 21232 4811
rect 21180 4768 21232 4777
rect 23664 4768 23716 4820
rect 30748 4768 30800 4820
rect 33232 4768 33284 4820
rect 34796 4768 34848 4820
rect 38292 4768 38344 4820
rect 6460 4700 6512 4752
rect 11980 4700 12032 4752
rect 6920 4632 6972 4684
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 4620 4564 4672 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 8852 4632 8904 4684
rect 9588 4632 9640 4684
rect 10508 4632 10560 4684
rect 4712 4564 4764 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 10876 4632 10928 4684
rect 11336 4632 11388 4684
rect 11428 4632 11480 4684
rect 11888 4632 11940 4684
rect 13544 4700 13596 4752
rect 14924 4700 14976 4752
rect 20076 4700 20128 4752
rect 12256 4675 12308 4684
rect 12256 4641 12265 4675
rect 12265 4641 12299 4675
rect 12299 4641 12308 4675
rect 12256 4632 12308 4641
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 11980 4564 12032 4616
rect 13636 4564 13688 4616
rect 17684 4632 17736 4684
rect 15016 4564 15068 4616
rect 15292 4564 15344 4616
rect 15568 4607 15620 4616
rect 15568 4573 15577 4607
rect 15577 4573 15611 4607
rect 15611 4573 15620 4607
rect 15568 4564 15620 4573
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17132 4564 17184 4616
rect 17500 4564 17552 4616
rect 20076 4564 20128 4616
rect 20260 4632 20312 4684
rect 21640 4675 21692 4684
rect 21640 4641 21649 4675
rect 21649 4641 21683 4675
rect 21683 4641 21692 4675
rect 21640 4632 21692 4641
rect 24216 4632 24268 4684
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 57244 4700 57296 4752
rect 58256 4700 58308 4752
rect 36636 4632 36688 4684
rect 26516 4564 26568 4616
rect 29000 4564 29052 4616
rect 31576 4564 31628 4616
rect 35164 4564 35216 4616
rect 2504 4428 2556 4480
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 11428 4496 11480 4548
rect 12348 4496 12400 4548
rect 14004 4496 14056 4548
rect 2780 4428 2832 4437
rect 7012 4428 7064 4480
rect 8116 4428 8168 4480
rect 8760 4428 8812 4480
rect 11704 4428 11756 4480
rect 13360 4471 13412 4480
rect 13360 4437 13369 4471
rect 13369 4437 13403 4471
rect 13403 4437 13412 4471
rect 13360 4428 13412 4437
rect 18972 4496 19024 4548
rect 19248 4496 19300 4548
rect 25228 4496 25280 4548
rect 25872 4496 25924 4548
rect 28172 4496 28224 4548
rect 30840 4496 30892 4548
rect 15752 4471 15804 4480
rect 15752 4437 15761 4471
rect 15761 4437 15795 4471
rect 15795 4437 15804 4471
rect 15752 4428 15804 4437
rect 16672 4471 16724 4480
rect 16672 4437 16681 4471
rect 16681 4437 16715 4471
rect 16715 4437 16724 4471
rect 16672 4428 16724 4437
rect 17500 4428 17552 4480
rect 17868 4471 17920 4480
rect 17868 4437 17877 4471
rect 17877 4437 17911 4471
rect 17911 4437 17920 4471
rect 17868 4428 17920 4437
rect 19616 4428 19668 4480
rect 20352 4428 20404 4480
rect 25688 4428 25740 4480
rect 28540 4428 28592 4480
rect 35348 4496 35400 4548
rect 34060 4471 34112 4480
rect 34060 4437 34069 4471
rect 34069 4437 34103 4471
rect 34103 4437 34112 4471
rect 34060 4428 34112 4437
rect 35532 4564 35584 4616
rect 37280 4607 37332 4616
rect 37280 4573 37289 4607
rect 37289 4573 37323 4607
rect 37323 4573 37332 4607
rect 37280 4564 37332 4573
rect 58900 4632 58952 4684
rect 57152 4564 57204 4616
rect 57612 4564 57664 4616
rect 36820 4471 36872 4480
rect 36820 4437 36829 4471
rect 36829 4437 36863 4471
rect 36863 4437 36872 4471
rect 36820 4428 36872 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 2136 4224 2188 4276
rect 7748 4224 7800 4276
rect 8852 4267 8904 4276
rect 8852 4233 8861 4267
rect 8861 4233 8895 4267
rect 8895 4233 8904 4267
rect 8852 4224 8904 4233
rect 8944 4267 8996 4276
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 9864 4224 9916 4276
rect 10416 4224 10468 4276
rect 10692 4267 10744 4276
rect 10692 4233 10717 4267
rect 10717 4233 10744 4267
rect 10876 4267 10928 4276
rect 10692 4224 10744 4233
rect 10876 4233 10885 4267
rect 10885 4233 10919 4267
rect 10919 4233 10928 4267
rect 10876 4224 10928 4233
rect 11428 4224 11480 4276
rect 12072 4224 12124 4276
rect 12348 4224 12400 4276
rect 13268 4224 13320 4276
rect 16856 4224 16908 4276
rect 17960 4224 18012 4276
rect 21640 4224 21692 4276
rect 26608 4224 26660 4276
rect 29000 4224 29052 4276
rect 33968 4224 34020 4276
rect 36268 4224 36320 4276
rect 2780 4156 2832 4208
rect 8760 4156 8812 4208
rect 10508 4199 10560 4208
rect 3148 4088 3200 4140
rect 4712 4088 4764 4140
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 7564 4088 7616 4140
rect 7748 4088 7800 4140
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 8116 4088 8168 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 2136 3884 2188 3936
rect 8760 4020 8812 4072
rect 9128 4020 9180 4072
rect 9680 4020 9732 4072
rect 10508 4165 10517 4199
rect 10517 4165 10551 4199
rect 10551 4165 10560 4199
rect 10508 4156 10560 4165
rect 11888 4156 11940 4208
rect 18236 4156 18288 4208
rect 20812 4199 20864 4208
rect 10600 4088 10652 4140
rect 12348 4088 12400 4140
rect 13452 4088 13504 4140
rect 14648 4088 14700 4140
rect 15292 4088 15344 4140
rect 16120 4088 16172 4140
rect 17500 4131 17552 4140
rect 17500 4097 17509 4131
rect 17509 4097 17543 4131
rect 17543 4097 17552 4131
rect 17500 4088 17552 4097
rect 17684 4131 17736 4140
rect 17684 4097 17693 4131
rect 17693 4097 17727 4131
rect 17727 4097 17736 4131
rect 17684 4088 17736 4097
rect 18788 4131 18840 4140
rect 11980 4020 12032 4072
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 20812 4165 20821 4199
rect 20821 4165 20855 4199
rect 20855 4165 20864 4199
rect 20812 4156 20864 4165
rect 20904 4199 20956 4208
rect 20904 4165 20913 4199
rect 20913 4165 20947 4199
rect 20947 4165 20956 4199
rect 20904 4156 20956 4165
rect 23480 4156 23532 4208
rect 19616 4131 19668 4140
rect 7748 3952 7800 4004
rect 9588 3952 9640 4004
rect 4804 3884 4856 3936
rect 6828 3884 6880 3936
rect 8208 3884 8260 3936
rect 12256 3952 12308 4004
rect 12900 3952 12952 4004
rect 17500 3952 17552 4004
rect 19340 4020 19392 4072
rect 19616 4097 19625 4131
rect 19625 4097 19659 4131
rect 19659 4097 19668 4131
rect 19616 4088 19668 4097
rect 21180 4088 21232 4140
rect 27620 4156 27672 4208
rect 31484 4156 31536 4208
rect 36820 4156 36872 4208
rect 19800 4020 19852 4072
rect 20444 4020 20496 4072
rect 20536 4020 20588 4072
rect 19524 3952 19576 4004
rect 20168 3952 20220 4004
rect 20812 3952 20864 4004
rect 24676 4088 24728 4140
rect 25412 4088 25464 4140
rect 25596 4131 25648 4140
rect 25596 4097 25605 4131
rect 25605 4097 25639 4131
rect 25639 4097 25648 4131
rect 25596 4088 25648 4097
rect 25688 4134 25740 4140
rect 25688 4100 25697 4134
rect 25697 4100 25731 4134
rect 25731 4100 25740 4134
rect 25688 4088 25740 4100
rect 26976 4088 27028 4140
rect 28356 4131 28408 4140
rect 28356 4097 28365 4131
rect 28365 4097 28399 4131
rect 28399 4097 28408 4131
rect 28356 4088 28408 4097
rect 28724 4088 28776 4140
rect 29000 4088 29052 4140
rect 31576 4088 31628 4140
rect 34520 4088 34572 4140
rect 35164 4131 35216 4140
rect 35164 4097 35173 4131
rect 35173 4097 35207 4131
rect 35207 4097 35216 4131
rect 35164 4088 35216 4097
rect 57980 4088 58032 4140
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 59176 4020 59228 4072
rect 11796 3884 11848 3936
rect 13268 3884 13320 3936
rect 13636 3884 13688 3936
rect 15016 3884 15068 3936
rect 18880 3884 18932 3936
rect 19340 3884 19392 3936
rect 20996 3884 21048 3936
rect 57520 3952 57572 4004
rect 58624 3952 58676 4004
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 56140 3884 56192 3936
rect 56324 3884 56376 3936
rect 56968 3884 57020 3936
rect 58072 3884 58124 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 2596 3680 2648 3732
rect 1860 3612 1912 3664
rect 4712 3680 4764 3732
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 7380 3680 7432 3732
rect 3240 3655 3292 3664
rect 3240 3621 3249 3655
rect 3249 3621 3283 3655
rect 3283 3621 3292 3655
rect 3240 3612 3292 3621
rect 1768 3544 1820 3596
rect 4804 3612 4856 3664
rect 5356 3612 5408 3664
rect 6368 3612 6420 3664
rect 9680 3612 9732 3664
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 7104 3544 7156 3596
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 7748 3544 7800 3596
rect 9312 3544 9364 3596
rect 9956 3612 10008 3664
rect 13084 3680 13136 3732
rect 14556 3680 14608 3732
rect 14648 3680 14700 3732
rect 12532 3612 12584 3664
rect 17868 3680 17920 3732
rect 18512 3612 18564 3664
rect 12072 3544 12124 3596
rect 12716 3544 12768 3596
rect 14188 3544 14240 3596
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 19616 3680 19668 3732
rect 19892 3680 19944 3732
rect 21180 3723 21232 3732
rect 21180 3689 21189 3723
rect 21189 3689 21223 3723
rect 21223 3689 21232 3723
rect 21180 3680 21232 3689
rect 29000 3723 29052 3732
rect 29000 3689 29009 3723
rect 29009 3689 29043 3723
rect 29043 3689 29052 3723
rect 29000 3680 29052 3689
rect 57796 3680 57848 3732
rect 58072 3680 58124 3732
rect 41144 3612 41196 3664
rect 56508 3612 56560 3664
rect 58348 3612 58400 3664
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 2964 3476 3016 3528
rect 3148 3476 3200 3528
rect 7564 3519 7616 3528
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 4896 3408 4948 3460
rect 5264 3408 5316 3460
rect 5540 3408 5592 3460
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 8208 3476 8260 3528
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 10324 3476 10376 3528
rect 11244 3519 11296 3528
rect 5724 3408 5776 3460
rect 6644 3408 6696 3460
rect 7840 3408 7892 3460
rect 6276 3340 6328 3392
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 9680 3340 9732 3392
rect 10140 3340 10192 3392
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 10692 3408 10744 3460
rect 10784 3451 10836 3460
rect 10784 3417 10793 3451
rect 10793 3417 10827 3451
rect 10827 3417 10836 3451
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 11888 3476 11940 3528
rect 13268 3476 13320 3528
rect 14372 3476 14424 3528
rect 14740 3476 14792 3528
rect 15752 3476 15804 3528
rect 16672 3476 16724 3528
rect 10784 3408 10836 3417
rect 12624 3408 12676 3460
rect 14004 3408 14056 3460
rect 19432 3544 19484 3596
rect 19984 3544 20036 3596
rect 20260 3544 20312 3596
rect 28264 3544 28316 3596
rect 11336 3340 11388 3392
rect 11612 3340 11664 3392
rect 11796 3340 11848 3392
rect 13084 3340 13136 3392
rect 13728 3340 13780 3392
rect 14556 3340 14608 3392
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 17224 3340 17276 3392
rect 17960 3340 18012 3392
rect 20168 3476 20220 3528
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 21824 3476 21876 3528
rect 22652 3476 22704 3528
rect 23480 3476 23532 3528
rect 24308 3476 24360 3528
rect 25136 3476 25188 3528
rect 25964 3476 26016 3528
rect 26792 3476 26844 3528
rect 27620 3476 27672 3528
rect 27896 3476 27948 3528
rect 28540 3519 28592 3528
rect 28540 3485 28549 3519
rect 28549 3485 28583 3519
rect 28583 3485 28592 3519
rect 28540 3476 28592 3485
rect 55772 3544 55824 3596
rect 56784 3544 56836 3596
rect 58992 3544 59044 3596
rect 28724 3519 28776 3528
rect 28724 3485 28733 3519
rect 28733 3485 28767 3519
rect 28767 3485 28776 3519
rect 28724 3476 28776 3485
rect 29828 3476 29880 3528
rect 30656 3476 30708 3528
rect 31484 3476 31536 3528
rect 32312 3476 32364 3528
rect 33140 3476 33192 3528
rect 39212 3476 39264 3528
rect 40040 3476 40092 3528
rect 40868 3476 40920 3528
rect 42524 3476 42576 3528
rect 43076 3476 43128 3528
rect 45008 3476 45060 3528
rect 45284 3476 45336 3528
rect 46112 3476 46164 3528
rect 46940 3476 46992 3528
rect 47768 3476 47820 3528
rect 48872 3476 48924 3528
rect 50160 3476 50212 3528
rect 50804 3476 50856 3528
rect 51356 3476 51408 3528
rect 52736 3476 52788 3528
rect 53012 3476 53064 3528
rect 54668 3476 54720 3528
rect 55496 3476 55548 3528
rect 56232 3476 56284 3528
rect 57336 3476 57388 3528
rect 60464 3519 60516 3528
rect 60464 3485 60473 3519
rect 60473 3485 60507 3519
rect 60507 3485 60516 3519
rect 60464 3476 60516 3485
rect 68100 3519 68152 3528
rect 68100 3485 68109 3519
rect 68109 3485 68143 3519
rect 68143 3485 68152 3519
rect 68100 3476 68152 3485
rect 19340 3451 19392 3460
rect 19340 3417 19349 3451
rect 19349 3417 19383 3451
rect 19383 3417 19392 3451
rect 19340 3408 19392 3417
rect 19432 3340 19484 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4620 3136 4672 3188
rect 4160 3068 4212 3120
rect 3148 3000 3200 3052
rect 7196 3136 7248 3188
rect 7656 3136 7708 3188
rect 7840 3136 7892 3188
rect 11428 3136 11480 3188
rect 12164 3136 12216 3188
rect 1768 2932 1820 2984
rect 2596 2932 2648 2984
rect 5540 2932 5592 2984
rect 6460 3000 6512 3052
rect 10232 3068 10284 3120
rect 11612 3068 11664 3120
rect 12624 3068 12676 3120
rect 13728 3068 13780 3120
rect 8300 3000 8352 3052
rect 8484 3043 8536 3052
rect 8484 3009 8518 3043
rect 8518 3009 8536 3043
rect 8484 3000 8536 3009
rect 12256 3000 12308 3052
rect 12440 3000 12492 3052
rect 14096 3136 14148 3188
rect 20904 3136 20956 3188
rect 55956 3136 56008 3188
rect 58072 3136 58124 3188
rect 14556 3068 14608 3120
rect 15936 3068 15988 3120
rect 16764 3000 16816 3052
rect 17316 3000 17368 3052
rect 57704 3068 57756 3120
rect 60464 3068 60516 3120
rect 20168 3000 20220 3052
rect 21732 3000 21784 3052
rect 58164 3000 58216 3052
rect 10600 2975 10652 2984
rect 4804 2907 4856 2916
rect 4804 2873 4813 2907
rect 4813 2873 4847 2907
rect 4847 2873 4856 2907
rect 4804 2864 4856 2873
rect 2596 2796 2648 2848
rect 10600 2941 10609 2975
rect 10609 2941 10643 2975
rect 10643 2941 10652 2975
rect 10600 2932 10652 2941
rect 12164 2975 12216 2984
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 11888 2864 11940 2916
rect 12256 2907 12308 2916
rect 12256 2873 12265 2907
rect 12265 2873 12299 2907
rect 12299 2873 12308 2907
rect 12256 2864 12308 2873
rect 12532 2864 12584 2916
rect 13452 2864 13504 2916
rect 14556 2975 14608 2984
rect 14556 2941 14565 2975
rect 14565 2941 14599 2975
rect 14599 2941 14608 2975
rect 14556 2932 14608 2941
rect 20260 2932 20312 2984
rect 21272 2932 21324 2984
rect 37280 2932 37332 2984
rect 44732 2932 44784 2984
rect 48596 2932 48648 2984
rect 52460 2932 52512 2984
rect 53564 2932 53616 2984
rect 55220 2932 55272 2984
rect 56692 2932 56744 2984
rect 8392 2796 8444 2848
rect 11980 2796 12032 2848
rect 14832 2864 14884 2916
rect 15660 2864 15712 2916
rect 20444 2864 20496 2916
rect 38384 2864 38436 2916
rect 39764 2864 39816 2916
rect 42248 2864 42300 2916
rect 43628 2864 43680 2916
rect 47492 2864 47544 2916
rect 49424 2864 49476 2916
rect 50620 2864 50672 2916
rect 53288 2864 53340 2916
rect 54392 2864 54444 2916
rect 55680 2864 55732 2916
rect 57060 2864 57112 2916
rect 58440 2932 58492 2984
rect 14004 2839 14056 2848
rect 14004 2805 14013 2839
rect 14013 2805 14047 2839
rect 14047 2805 14056 2839
rect 14004 2796 14056 2805
rect 14188 2796 14240 2848
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 15844 2796 15896 2848
rect 18696 2796 18748 2848
rect 20720 2796 20772 2848
rect 21548 2796 21600 2848
rect 22928 2796 22980 2848
rect 23756 2796 23808 2848
rect 24032 2796 24084 2848
rect 24860 2796 24912 2848
rect 25688 2796 25740 2848
rect 26240 2796 26292 2848
rect 27068 2796 27120 2848
rect 28172 2796 28224 2848
rect 28724 2796 28776 2848
rect 29276 2796 29328 2848
rect 30104 2796 30156 2848
rect 30380 2796 30432 2848
rect 31208 2796 31260 2848
rect 32036 2796 32088 2848
rect 32864 2839 32916 2848
rect 32864 2805 32873 2839
rect 32873 2805 32907 2839
rect 32907 2805 32916 2839
rect 32864 2796 32916 2805
rect 33692 2796 33744 2848
rect 34244 2796 34296 2848
rect 34520 2796 34572 2848
rect 35348 2796 35400 2848
rect 36176 2796 36228 2848
rect 36728 2796 36780 2848
rect 37832 2796 37884 2848
rect 38936 2796 38988 2848
rect 40316 2796 40368 2848
rect 41696 2796 41748 2848
rect 42800 2796 42852 2848
rect 44180 2796 44232 2848
rect 45560 2796 45612 2848
rect 46664 2796 46716 2848
rect 48044 2796 48096 2848
rect 49976 2796 50028 2848
rect 51908 2796 51960 2848
rect 53840 2796 53892 2848
rect 55404 2796 55456 2848
rect 56048 2796 56100 2848
rect 59360 2864 59412 2916
rect 59452 2796 59504 2848
rect 60464 2839 60516 2848
rect 60464 2805 60473 2839
rect 60473 2805 60507 2839
rect 60507 2805 60516 2839
rect 60464 2796 60516 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 4620 2592 4672 2644
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 6644 2592 6696 2644
rect 8300 2592 8352 2644
rect 11244 2592 11296 2644
rect 12256 2592 12308 2644
rect 15016 2592 15068 2644
rect 17132 2592 17184 2644
rect 8116 2524 8168 2576
rect 10784 2524 10836 2576
rect 12440 2524 12492 2576
rect 14464 2524 14516 2576
rect 2504 2456 2556 2508
rect 12164 2456 12216 2508
rect 14096 2456 14148 2508
rect 14556 2456 14608 2508
rect 1492 2388 1544 2440
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 4988 2388 5040 2440
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 5908 2388 5960 2440
rect 6184 2388 6236 2440
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 8024 2388 8076 2440
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 10508 2388 10560 2440
rect 11520 2388 11572 2440
rect 11980 2388 12032 2440
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 13084 2388 13136 2440
rect 16028 2431 16080 2440
rect 11060 2320 11112 2372
rect 12164 2320 12216 2372
rect 14556 2363 14608 2372
rect 14556 2329 14565 2363
rect 14565 2329 14599 2363
rect 14599 2329 14608 2363
rect 14556 2320 14608 2329
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 18236 2567 18288 2576
rect 18236 2533 18245 2567
rect 18245 2533 18279 2567
rect 18279 2533 18288 2567
rect 18236 2524 18288 2533
rect 19984 2592 20036 2644
rect 21732 2592 21784 2644
rect 21916 2592 21968 2644
rect 55220 2592 55272 2644
rect 57428 2592 57480 2644
rect 20536 2524 20588 2576
rect 22100 2524 22152 2576
rect 23204 2524 23256 2576
rect 27344 2524 27396 2576
rect 29000 2524 29052 2576
rect 30932 2524 30984 2576
rect 40592 2524 40644 2576
rect 44456 2524 44508 2576
rect 48320 2524 48372 2576
rect 52184 2524 52236 2576
rect 55864 2524 55916 2576
rect 58072 2524 58124 2576
rect 17868 2456 17920 2508
rect 21916 2456 21968 2508
rect 22008 2456 22060 2508
rect 26516 2456 26568 2508
rect 37004 2456 37056 2508
rect 38108 2456 38160 2508
rect 41420 2456 41472 2508
rect 43352 2456 43404 2508
rect 46388 2456 46440 2508
rect 49148 2456 49200 2508
rect 51080 2456 51132 2508
rect 54944 2456 54996 2508
rect 63684 2499 63736 2508
rect 20996 2388 21048 2440
rect 22376 2388 22428 2440
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 3884 2295 3936 2304
rect 3884 2261 3893 2295
rect 3893 2261 3927 2295
rect 3927 2261 3936 2295
rect 3884 2252 3936 2261
rect 10324 2252 10376 2304
rect 13728 2252 13780 2304
rect 22008 2320 22060 2372
rect 25412 2388 25464 2440
rect 24584 2320 24636 2372
rect 28448 2388 28500 2440
rect 29552 2388 29604 2440
rect 27896 2320 27948 2372
rect 32588 2388 32640 2440
rect 33416 2388 33468 2440
rect 33968 2388 34020 2440
rect 34796 2388 34848 2440
rect 35072 2388 35124 2440
rect 35624 2388 35676 2440
rect 35900 2388 35952 2440
rect 36452 2388 36504 2440
rect 37556 2388 37608 2440
rect 38660 2388 38712 2440
rect 31760 2320 31812 2372
rect 39488 2320 39540 2372
rect 41972 2388 42024 2440
rect 43904 2320 43956 2372
rect 45836 2388 45888 2440
rect 47216 2320 47268 2372
rect 49700 2388 49752 2440
rect 51632 2388 51684 2440
rect 54116 2320 54168 2372
rect 56416 2388 56468 2440
rect 17592 2252 17644 2304
rect 56876 2252 56928 2304
rect 63684 2465 63693 2499
rect 63693 2465 63727 2499
rect 63727 2465 63736 2499
rect 63684 2456 63736 2465
rect 61752 2431 61804 2440
rect 61752 2397 61761 2431
rect 61761 2397 61795 2431
rect 61795 2397 61804 2431
rect 61752 2388 61804 2397
rect 63040 2431 63092 2440
rect 63040 2397 63049 2431
rect 63049 2397 63083 2431
rect 63083 2397 63092 2431
rect 63040 2388 63092 2397
rect 66996 2431 67048 2440
rect 66996 2397 67005 2431
rect 67005 2397 67039 2431
rect 67039 2397 67048 2431
rect 66996 2388 67048 2397
rect 67548 2388 67600 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 6644 2048 6696 2100
rect 11244 2048 11296 2100
rect 3884 1980 3936 2032
rect 11980 1980 12032 2032
rect 14556 2048 14608 2100
rect 18788 2048 18840 2100
rect 19800 2048 19852 2100
rect 58072 2048 58124 2100
rect 61752 2048 61804 2100
rect 17592 1980 17644 2032
rect 24676 1980 24728 2032
rect 59084 1980 59136 2032
rect 63684 1980 63736 2032
rect 5080 1912 5132 1964
rect 14648 1912 14700 1964
rect 58532 1912 58584 1964
rect 63040 1912 63092 1964
rect 5632 1844 5684 1896
rect 12716 1844 12768 1896
rect 3240 1776 3292 1828
rect 12624 1776 12676 1828
rect 9680 1708 9732 1760
rect 8116 1640 8168 1692
rect 10048 1640 10100 1692
rect 9772 1572 9824 1624
rect 10692 1572 10744 1624
rect 10324 1436 10376 1488
rect 10140 1368 10192 1420
rect 10876 1368 10928 1420
rect 12440 1368 12492 1420
rect 12716 1368 12768 1420
rect 14280 1436 14332 1488
rect 15016 1436 15068 1488
rect 12900 1300 12952 1352
rect 12992 1300 13044 1352
rect 12716 1232 12768 1284
rect 13728 1368 13780 1420
rect 14188 1368 14240 1420
rect 14832 1368 14884 1420
rect 19524 1300 19576 1352
rect 20352 1300 20404 1352
rect 12808 1164 12860 1216
rect 15660 1164 15712 1216
rect 56784 1164 56836 1216
rect 57060 1164 57112 1216
rect 12348 1096 12400 1148
rect 19340 1096 19392 1148
rect 19708 1096 19760 1148
rect 12256 892 12308 944
rect 57060 1028 57112 1080
rect 59452 1028 59504 1080
<< metal2 >>
rect 5170 59200 5226 60000
rect 15106 59200 15162 60000
rect 25042 59200 25098 60000
rect 34978 59200 35034 60000
rect 44914 59200 44970 60000
rect 54850 59200 54906 60000
rect 64786 59200 64842 60000
rect 67546 59256 67602 59265
rect 5184 57458 5212 59200
rect 15120 57882 15148 59200
rect 15120 57854 15240 57882
rect 15212 57458 15240 57854
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 25056 57458 25084 59200
rect 34992 57458 35020 59200
rect 44928 57458 44956 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 54864 57458 54892 59200
rect 64800 57458 64828 59200
rect 67546 59191 67602 59200
rect 66994 57896 67050 57905
rect 66994 57831 67050 57840
rect 67008 57458 67036 57831
rect 67560 57458 67588 59191
rect 5172 57452 5224 57458
rect 5172 57394 5224 57400
rect 15200 57452 15252 57458
rect 15200 57394 15252 57400
rect 25044 57452 25096 57458
rect 25044 57394 25096 57400
rect 34980 57452 35032 57458
rect 34980 57394 35032 57400
rect 44916 57452 44968 57458
rect 44916 57394 44968 57400
rect 54852 57452 54904 57458
rect 54852 57394 54904 57400
rect 64788 57452 64840 57458
rect 64788 57394 64840 57400
rect 66996 57452 67048 57458
rect 66996 57394 67048 57400
rect 67548 57452 67600 57458
rect 67548 57394 67600 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 68100 56840 68152 56846
rect 68100 56782 68152 56788
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 68112 56545 68140 56782
rect 68098 56536 68154 56545
rect 68098 56471 68154 56480
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 67638 55176 67694 55185
rect 67638 55111 67640 55120
rect 67692 55111 67694 55120
rect 67640 55082 67692 55088
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 67548 53984 67600 53990
rect 67548 53926 67600 53932
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 67560 53825 67588 53926
rect 67546 53816 67602 53825
rect 67546 53751 67602 53760
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 68100 52488 68152 52494
rect 68098 52456 68100 52465
rect 68152 52456 68154 52465
rect 68098 52391 68154 52400
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 68100 51400 68152 51406
rect 68100 51342 68152 51348
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 68112 51105 68140 51342
rect 68098 51096 68154 51105
rect 68098 51031 68154 51040
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 67640 49768 67692 49774
rect 67638 49736 67640 49745
rect 67692 49736 67694 49745
rect 67638 49671 67694 49680
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 67640 48544 67692 48550
rect 67640 48486 67692 48492
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 67652 48385 67680 48486
rect 67638 48376 67694 48385
rect 67638 48311 67694 48320
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 68100 47048 68152 47054
rect 68098 47016 68100 47025
rect 68152 47016 68154 47025
rect 68098 46951 68154 46960
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 68100 45960 68152 45966
rect 68100 45902 68152 45908
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 68112 45665 68140 45902
rect 68098 45656 68154 45665
rect 68098 45591 68154 45600
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 67638 44296 67694 44305
rect 67638 44231 67640 44240
rect 67692 44231 67694 44240
rect 67640 44202 67692 44208
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 67640 43104 67692 43110
rect 67640 43046 67692 43052
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 67652 42945 67680 43046
rect 67638 42936 67694 42945
rect 67638 42871 67694 42880
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 68100 41608 68152 41614
rect 68098 41576 68100 41585
rect 68152 41576 68154 41585
rect 68098 41511 68154 41520
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 68100 40520 68152 40526
rect 68100 40462 68152 40468
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 68112 40225 68140 40462
rect 68098 40216 68154 40225
rect 68098 40151 68154 40160
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 67638 38856 67694 38865
rect 67638 38791 67640 38800
rect 67692 38791 67694 38800
rect 67640 38762 67692 38768
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 67640 37664 67692 37670
rect 67640 37606 67692 37612
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 67652 37505 67680 37606
rect 67638 37496 67694 37505
rect 67638 37431 67694 37440
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 68100 36168 68152 36174
rect 68098 36136 68100 36145
rect 68152 36136 68154 36145
rect 68098 36071 68154 36080
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 68100 35080 68152 35086
rect 68100 35022 68152 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 68112 34785 68140 35022
rect 68098 34776 68154 34785
rect 68098 34711 68154 34720
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 67638 33416 67694 33425
rect 67638 33351 67640 33360
rect 67692 33351 67694 33360
rect 67640 33322 67692 33328
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 67640 32224 67692 32230
rect 67640 32166 67692 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 67652 32065 67680 32166
rect 67638 32056 67694 32065
rect 67638 31991 67694 32000
rect 15108 31748 15160 31754
rect 15108 31690 15160 31696
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 7840 31408 7892 31414
rect 7840 31350 7892 31356
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 7852 30394 7880 31350
rect 8392 31340 8444 31346
rect 8392 31282 8444 31288
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 13176 31340 13228 31346
rect 13228 31300 13308 31328
rect 13176 31282 13228 31288
rect 8404 30734 8432 31282
rect 9404 31136 9456 31142
rect 9404 31078 9456 31084
rect 9312 30932 9364 30938
rect 9312 30874 9364 30880
rect 9324 30734 9352 30874
rect 8392 30728 8444 30734
rect 8392 30670 8444 30676
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 8208 30660 8260 30666
rect 8208 30602 8260 30608
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 3792 30252 3844 30258
rect 3792 30194 3844 30200
rect 3804 29714 3832 30194
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3792 29708 3844 29714
rect 3792 29650 3844 29656
rect 3332 29572 3384 29578
rect 3332 29514 3384 29520
rect 1768 28484 1820 28490
rect 1768 28426 1820 28432
rect 3240 28484 3292 28490
rect 3240 28426 3292 28432
rect 1780 28082 1808 28426
rect 2228 28416 2280 28422
rect 2228 28358 2280 28364
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1780 26314 1808 28018
rect 2240 27470 2268 28358
rect 3252 28218 3280 28426
rect 3240 28212 3292 28218
rect 3240 28154 3292 28160
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2332 27334 2360 28018
rect 2596 27600 2648 27606
rect 2596 27542 2648 27548
rect 2608 27470 2636 27542
rect 2884 27538 2912 28018
rect 3344 27606 3372 29514
rect 5172 29504 5224 29510
rect 5172 29446 5224 29452
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5184 28694 5212 29446
rect 6736 29300 6788 29306
rect 6736 29242 6788 29248
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6656 28762 6684 29106
rect 6644 28756 6696 28762
rect 6644 28698 6696 28704
rect 5172 28688 5224 28694
rect 5172 28630 5224 28636
rect 3424 28552 3476 28558
rect 3424 28494 3476 28500
rect 3332 27600 3384 27606
rect 3332 27542 3384 27548
rect 2872 27532 2924 27538
rect 2872 27474 2924 27480
rect 2596 27464 2648 27470
rect 2596 27406 2648 27412
rect 2320 27328 2372 27334
rect 2320 27270 2372 27276
rect 2332 26994 2360 27270
rect 2320 26988 2372 26994
rect 2320 26930 2372 26936
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 1768 26308 1820 26314
rect 1768 26250 1820 26256
rect 1780 25974 1808 26250
rect 1768 25968 1820 25974
rect 1768 25910 1820 25916
rect 1780 24886 1808 25910
rect 2332 25906 2360 26930
rect 2516 26586 2544 26930
rect 2504 26580 2556 26586
rect 2504 26522 2556 26528
rect 2320 25900 2372 25906
rect 2320 25842 2372 25848
rect 2332 25294 2360 25842
rect 2320 25288 2372 25294
rect 2320 25230 2372 25236
rect 1768 24880 1820 24886
rect 1768 24822 1820 24828
rect 1780 24410 1808 24822
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 2332 23730 2360 25230
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2320 23724 2372 23730
rect 2320 23666 2372 23672
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 1596 21554 1624 23054
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 2148 22030 2176 22578
rect 2332 22234 2360 23054
rect 2516 22982 2544 24074
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 2320 22228 2372 22234
rect 2320 22170 2372 22176
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 1768 21956 1820 21962
rect 1768 21898 1820 21904
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1688 21554 1716 21830
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1596 20466 1624 21490
rect 1780 20874 1808 21898
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 1768 20868 1820 20874
rect 1768 20810 1820 20816
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 19854 1624 20198
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1780 19446 1808 20810
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2240 20466 2268 20742
rect 2332 20466 2360 21354
rect 2516 20942 2544 22918
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2320 20460 2372 20466
rect 2320 20402 2372 20408
rect 2056 19854 2084 20402
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 1768 19440 1820 19446
rect 1768 19382 1820 19388
rect 2056 18834 2084 19790
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2148 18290 2176 20334
rect 2332 19990 2360 20402
rect 2320 19984 2372 19990
rect 2320 19926 2372 19932
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2044 17672 2096 17678
rect 2148 17660 2176 18226
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2240 17814 2268 18158
rect 2228 17808 2280 17814
rect 2228 17750 2280 17756
rect 2096 17632 2176 17660
rect 2044 17614 2096 17620
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1596 15434 1624 17138
rect 2056 16658 2084 17614
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2056 16114 2084 16594
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2056 15502 2084 16050
rect 2240 16046 2268 17750
rect 2332 17338 2360 18226
rect 2424 17354 2452 19722
rect 2516 19514 2544 19790
rect 2608 19700 2636 27406
rect 2884 26926 2912 27474
rect 3436 26994 3464 28494
rect 5184 28422 5212 28630
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5172 28416 5224 28422
rect 5172 28358 5224 28364
rect 5368 28082 5396 28494
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 28150 5488 28358
rect 5448 28144 5500 28150
rect 5448 28086 5500 28092
rect 6748 28082 6776 29242
rect 6840 29238 6868 30126
rect 6828 29232 6880 29238
rect 6828 29174 6880 29180
rect 7288 28960 7340 28966
rect 7288 28902 7340 28908
rect 7300 28558 7328 28902
rect 7852 28558 7880 30330
rect 8220 30054 8248 30602
rect 9128 30592 9180 30598
rect 9128 30534 9180 30540
rect 9140 30326 9168 30534
rect 9128 30320 9180 30326
rect 9128 30262 9180 30268
rect 9416 30258 9444 31078
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 9692 30666 9720 30738
rect 9772 30728 9824 30734
rect 9770 30696 9772 30705
rect 9824 30696 9826 30705
rect 9680 30660 9732 30666
rect 9770 30631 9826 30640
rect 9680 30602 9732 30608
rect 9692 30326 9720 30602
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 9680 30320 9732 30326
rect 9680 30262 9732 30268
rect 10416 30320 10468 30326
rect 10416 30262 10468 30268
rect 9404 30252 9456 30258
rect 9404 30194 9456 30200
rect 8208 30048 8260 30054
rect 8208 29990 8260 29996
rect 8116 28688 8168 28694
rect 8116 28630 8168 28636
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7840 28552 7892 28558
rect 7840 28494 7892 28500
rect 7024 28218 7052 28494
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 5644 27674 5672 28018
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 5632 27668 5684 27674
rect 5632 27610 5684 27616
rect 6552 27396 6604 27402
rect 6552 27338 6604 27344
rect 6564 27130 6592 27338
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 3424 26988 3476 26994
rect 6840 26976 6868 27814
rect 7012 26988 7064 26994
rect 6840 26948 7012 26976
rect 3424 26930 3476 26936
rect 7012 26930 7064 26936
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 2884 25906 2912 26862
rect 3436 26450 3464 26930
rect 3700 26784 3752 26790
rect 3700 26726 3752 26732
rect 3712 26518 3740 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5172 26580 5224 26586
rect 5172 26522 5224 26528
rect 3700 26512 3752 26518
rect 3700 26454 3752 26460
rect 3424 26444 3476 26450
rect 3424 26386 3476 26392
rect 3792 26444 3844 26450
rect 3792 26386 3844 26392
rect 3240 26308 3292 26314
rect 3240 26250 3292 26256
rect 3252 26042 3280 26250
rect 3240 26036 3292 26042
rect 3240 25978 3292 25984
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2884 25294 2912 25842
rect 3804 25362 3832 26386
rect 5184 25974 5212 26522
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 5724 26240 5776 26246
rect 5724 26182 5776 26188
rect 5172 25968 5224 25974
rect 5172 25910 5224 25916
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 5736 25498 5764 26182
rect 6840 26042 6868 26318
rect 6920 26308 6972 26314
rect 6920 26250 6972 26256
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 6828 25900 6880 25906
rect 6828 25842 6880 25848
rect 5724 25492 5776 25498
rect 5724 25434 5776 25440
rect 3792 25356 3844 25362
rect 3792 25298 3844 25304
rect 2872 25288 2924 25294
rect 2924 25248 3004 25276
rect 2872 25230 2924 25236
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 24954 2912 25094
rect 2872 24948 2924 24954
rect 2872 24890 2924 24896
rect 2976 24410 3004 25248
rect 2964 24404 3016 24410
rect 2964 24346 3016 24352
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 2872 24132 2924 24138
rect 2792 24092 2872 24120
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2700 23050 2728 24006
rect 2688 23044 2740 23050
rect 2688 22986 2740 22992
rect 2700 21350 2728 22986
rect 2792 21894 2820 24092
rect 2872 24074 2924 24080
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2976 21978 3004 23054
rect 2976 21950 3096 21978
rect 3068 21894 3096 21950
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 2792 21486 2820 21830
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 3068 20806 3096 21830
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2688 19712 2740 19718
rect 2608 19672 2688 19700
rect 2688 19654 2740 19660
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2608 18873 2636 19450
rect 2594 18864 2650 18873
rect 2594 18799 2650 18808
rect 2700 17678 2728 19654
rect 2976 19446 3004 19654
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 3160 18834 3188 23462
rect 3344 23186 3372 24142
rect 3804 23730 3832 25298
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4724 24614 4752 24754
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3804 23186 3832 23666
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3804 22710 3832 23122
rect 3988 22778 4016 24142
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4448 23798 4476 24006
rect 4436 23792 4488 23798
rect 4436 23734 4488 23740
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4632 22778 4660 22986
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 3792 22704 3844 22710
rect 3792 22646 3844 22652
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3252 21690 3280 22578
rect 3804 22166 3832 22646
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 4632 22098 4660 22714
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3344 20448 3372 21830
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 3436 20602 3464 20810
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3424 20460 3476 20466
rect 3344 20420 3424 20448
rect 3424 20402 3476 20408
rect 3896 19378 3924 20878
rect 4632 20602 4660 21898
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3160 18630 3188 18770
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2502 17368 2558 17377
rect 2320 17332 2372 17338
rect 2424 17326 2502 17354
rect 2502 17303 2558 17312
rect 2320 17274 2372 17280
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 1584 15428 1636 15434
rect 1584 15370 1636 15376
rect 1676 15428 1728 15434
rect 1676 15370 1728 15376
rect 1596 14278 1624 15370
rect 1688 14890 1716 15370
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13326 1624 14214
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 12238 1440 12582
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 10742 1440 12174
rect 1780 11762 1808 13874
rect 1964 13530 1992 13874
rect 2240 13870 2268 14894
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2332 12850 2360 14214
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 11762 2268 12038
rect 2424 11898 2452 12106
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1400 10736 1452 10742
rect 1400 10678 1452 10684
rect 1412 10062 1440 10678
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9722 1440 9998
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1780 9654 1808 10406
rect 1872 10062 1900 10746
rect 2056 10062 2084 11698
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 2056 9586 2084 9998
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2056 9042 2084 9522
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2056 8498 2084 8978
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1504 2446 1532 7686
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 6322 1992 6598
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1780 5234 1808 6190
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1780 3602 1808 5170
rect 1872 4078 1900 5714
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1964 5234 1992 5510
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 2148 4282 2176 7754
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 6458 2268 7346
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 5778 2360 6802
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 1860 4072 1912 4078
rect 2148 4049 2176 4218
rect 1860 4014 1912 4020
rect 2134 4040 2190 4049
rect 1872 3670 1900 4014
rect 2134 3975 2190 3984
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 1860 3664 1912 3670
rect 1860 3606 1912 3612
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 2990 1808 3538
rect 2148 3534 2176 3878
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 2424 2446 2452 7686
rect 2516 6730 2544 17303
rect 2608 17270 2636 17478
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2700 17202 2728 17478
rect 2792 17338 2820 17546
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 16114 2820 16390
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2596 15972 2648 15978
rect 2596 15914 2648 15920
rect 2608 15502 2636 15914
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 14958 2636 15438
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2792 14006 2820 14962
rect 2780 14000 2832 14006
rect 2700 13960 2780 13988
rect 2700 13462 2728 13960
rect 2780 13942 2832 13948
rect 2792 13877 2820 13942
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2608 12102 2636 13262
rect 2792 12374 2820 13738
rect 2884 12434 2912 16662
rect 2976 15706 3004 17546
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3068 16998 3096 17138
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3160 16726 3188 18566
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3252 16726 3280 18226
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3620 17746 3648 18158
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3620 17202 3648 17682
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3344 16250 3372 16730
rect 3528 16590 3556 17070
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3804 16289 3832 18566
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3790 16280 3846 16289
rect 3332 16244 3384 16250
rect 3790 16215 3846 16224
rect 3332 16186 3384 16192
rect 3804 16182 3832 16215
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 4528 16108 4580 16114
rect 4632 16096 4660 17138
rect 4580 16068 4660 16096
rect 4528 16050 4580 16056
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 3160 15026 3188 15302
rect 3712 15026 3740 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2976 13870 3004 14894
rect 3804 14482 3832 15438
rect 3988 15366 4016 15438
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3896 14618 3924 14962
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 4080 14414 4108 15438
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14414 4660 14758
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3068 12986 3096 13874
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3896 12850 3924 13670
rect 4080 13394 4108 14350
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 12986 4108 13330
rect 4632 13326 4660 13806
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 2884 12406 3004 12434
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11830 2636 12038
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2608 9926 2636 11766
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2700 10282 2728 11698
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2884 11218 2912 11630
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2700 10254 2820 10282
rect 2792 10010 2820 10254
rect 2700 9982 2820 10010
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 9518 2636 9862
rect 2700 9722 2728 9982
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 8362 2636 9454
rect 2700 8974 2728 9658
rect 2976 9042 3004 12406
rect 3804 12306 3832 12786
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12434 4752 24550
rect 4816 22094 4844 24618
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 5184 23594 5212 24210
rect 5644 23866 5672 25230
rect 5736 24750 5764 25434
rect 5724 24744 5776 24750
rect 5724 24686 5776 24692
rect 6656 24614 6684 25842
rect 6840 25498 6868 25842
rect 6932 25702 6960 26250
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 6920 25696 6972 25702
rect 6920 25638 6972 25644
rect 6828 25492 6880 25498
rect 6828 25434 6880 25440
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6644 24608 6696 24614
rect 6644 24550 6696 24556
rect 6656 24342 6684 24550
rect 6644 24336 6696 24342
rect 6644 24278 6696 24284
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 5632 23860 5684 23866
rect 5632 23802 5684 23808
rect 5644 23712 5672 23802
rect 5644 23684 5764 23712
rect 5172 23588 5224 23594
rect 5172 23530 5224 23536
rect 5632 23588 5684 23594
rect 5632 23530 5684 23536
rect 5184 22438 5212 23530
rect 5644 23322 5672 23530
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 22778 5488 22918
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 4816 22066 4936 22094
rect 4804 21412 4856 21418
rect 4804 21354 4856 21360
rect 4816 20534 4844 21354
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4908 18630 4936 22066
rect 5460 21622 5488 22714
rect 5448 21616 5500 21622
rect 5448 21558 5500 21564
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5092 19378 5120 20198
rect 5448 19848 5500 19854
rect 5552 19825 5580 23054
rect 5644 22030 5672 23258
rect 5736 23118 5764 23684
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5920 21350 5948 22510
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21554 6592 21830
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 5736 20262 5764 20742
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5448 19790 5500 19796
rect 5538 19816 5594 19825
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4807 16108 4859 16114
rect 4807 16050 4859 16056
rect 4816 15094 4844 16050
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4816 14414 4844 15030
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4724 12406 4844 12434
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3068 11626 3096 12106
rect 3252 11898 3280 12174
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 3160 10810 3188 11630
rect 3988 11354 4016 12242
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3988 10674 4016 11290
rect 4724 10674 4752 12038
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 3160 10266 3188 10610
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3884 9580 3936 9586
rect 3988 9568 4016 10610
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3936 9540 4016 9568
rect 3884 9522 3936 9528
rect 3988 9042 4016 9540
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 3252 8838 3280 8978
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 3160 8090 3188 8434
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2792 5642 2820 6394
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2516 2514 2544 4422
rect 2608 3738 2636 4558
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4214 2820 4422
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2964 3528 3016 3534
rect 2962 3496 2964 3505
rect 3016 3496 3018 3505
rect 2962 3431 3018 3440
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2608 2854 2636 2926
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 3068 2446 3096 7210
rect 3160 5710 3188 7278
rect 3252 6866 3280 8774
rect 3344 8566 3372 8774
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3896 8090 3924 8910
rect 3988 8566 4016 8978
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3160 4146 3188 5646
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3160 3534 3188 4082
rect 3252 3670 3280 6326
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3436 4321 3464 4966
rect 3422 4312 3478 4321
rect 3422 4247 3478 4256
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3148 3528 3200 3534
rect 3896 3505 3924 7686
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3148 3470 3200 3476
rect 3882 3496 3938 3505
rect 3160 3058 3188 3470
rect 3882 3431 3938 3440
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3988 2774 4016 6394
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4080 5574 4108 6190
rect 4448 6118 4476 6938
rect 4632 6798 4660 7142
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4172 5370 4200 5578
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4724 4729 4752 6598
rect 4816 6458 4844 12406
rect 5092 11150 5120 19314
rect 5276 18630 5304 19722
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5184 15706 5212 16186
rect 5276 15994 5304 18566
rect 5368 18154 5396 19110
rect 5460 18737 5488 19790
rect 5538 19751 5594 19760
rect 5552 19718 5580 19751
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5446 18728 5502 18737
rect 5446 18663 5502 18672
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5368 17746 5396 18090
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5460 17542 5488 18022
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5368 16114 5396 16662
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5276 15966 5396 15994
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5184 15094 5212 15642
rect 5276 15502 5304 15846
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5368 12986 5396 15966
rect 5460 15910 5488 17478
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5552 14074 5580 19654
rect 5828 19514 5856 20266
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5828 14074 5856 18158
rect 5920 17241 5948 21286
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6460 20256 6512 20262
rect 6460 20198 6512 20204
rect 6472 19854 6500 20198
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6196 19446 6224 19654
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 6472 19174 6500 19790
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6564 18698 6592 20402
rect 6656 19446 6684 24074
rect 6748 24070 6776 24754
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6748 23712 6776 24006
rect 6828 23724 6880 23730
rect 6748 23684 6828 23712
rect 6748 22642 6776 23684
rect 6828 23666 6880 23672
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6828 23248 6880 23254
rect 6828 23190 6880 23196
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6748 22234 6776 22578
rect 6736 22228 6788 22234
rect 6736 22170 6788 22176
rect 6748 21010 6776 22170
rect 6840 22098 6868 23190
rect 6932 23118 6960 23462
rect 7024 23118 7052 25842
rect 7116 25226 7144 27950
rect 7300 26994 7328 28494
rect 7380 28484 7432 28490
rect 7380 28426 7432 28432
rect 7392 27334 7420 28426
rect 8128 28218 8156 28630
rect 8116 28212 8168 28218
rect 8116 28154 8168 28160
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7944 27470 7972 27814
rect 7748 27464 7800 27470
rect 7748 27406 7800 27412
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 7380 27328 7432 27334
rect 7380 27270 7432 27276
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 7104 25220 7156 25226
rect 7104 25162 7156 25168
rect 7116 24682 7144 25162
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 7116 23866 7144 24618
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7116 22574 7144 22986
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6748 19854 6776 20198
rect 7116 19990 7144 22510
rect 7196 21956 7248 21962
rect 7196 21898 7248 21904
rect 7208 21865 7236 21898
rect 7194 21856 7250 21865
rect 7194 21791 7250 21800
rect 7208 20534 7236 21791
rect 7196 20528 7248 20534
rect 7196 20470 7248 20476
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 19440 6696 19446
rect 6642 19408 6644 19417
rect 6696 19408 6698 19417
rect 6642 19343 6698 19352
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6932 18970 6960 19246
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 5906 17232 5962 17241
rect 5906 17167 5962 17176
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6196 14550 6224 14962
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 6196 14414 6224 14486
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6472 14074 6500 14282
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6564 13870 6592 18634
rect 6932 18426 6960 18702
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 7300 18222 7328 26930
rect 7392 26926 7420 27270
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7392 25838 7420 26862
rect 7484 26586 7512 26862
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7760 25906 7788 27406
rect 8036 27334 8064 27406
rect 8024 27328 8076 27334
rect 8024 27270 8076 27276
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 7392 24682 7420 25774
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7380 24676 7432 24682
rect 7380 24618 7432 24624
rect 7392 23186 7420 24618
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7484 23322 7512 23666
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7576 23202 7604 24686
rect 7760 23254 7788 24686
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7748 23248 7800 23254
rect 7380 23180 7432 23186
rect 7576 23174 7696 23202
rect 7748 23190 7800 23196
rect 7380 23122 7432 23128
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7484 19922 7512 23054
rect 7564 22568 7616 22574
rect 7564 22510 7616 22516
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7484 18748 7512 19722
rect 7576 18902 7604 22510
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7564 18760 7616 18766
rect 7484 18720 7564 18748
rect 7564 18702 7616 18708
rect 7576 18290 7604 18702
rect 7668 18358 7696 23174
rect 7760 22574 7788 23190
rect 7852 23118 7880 24142
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7932 22500 7984 22506
rect 7932 22442 7984 22448
rect 7944 22030 7972 22442
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7852 20874 7880 21490
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 7760 20602 7788 20810
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 7944 20466 7972 20538
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6656 15706 6684 16050
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6748 15026 6776 17478
rect 6840 17338 6868 17614
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6840 14958 6868 16050
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7024 15434 7052 15506
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 7024 15026 7052 15370
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14414 6868 14894
rect 7116 14414 7144 17682
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7300 17202 7328 17614
rect 7576 17542 7604 18226
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7392 16425 7420 16458
rect 7378 16416 7434 16425
rect 7378 16351 7434 16360
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7392 15502 7420 15846
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7300 15094 7328 15370
rect 7484 15162 7512 17138
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7300 14414 7328 15030
rect 7576 14550 7604 17138
rect 7654 15736 7710 15745
rect 7654 15671 7656 15680
rect 7708 15671 7710 15680
rect 7656 15642 7708 15648
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7116 13938 7144 14214
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5368 11898 5396 12922
rect 6932 12850 6960 13126
rect 7208 12850 7236 13942
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6656 12238 6684 12582
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5828 11286 5856 11698
rect 6564 11354 6592 12174
rect 7208 11898 7236 12786
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 5092 10062 5120 11086
rect 5828 10810 5856 11222
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6564 10742 6592 11290
rect 6932 11082 6960 11494
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7024 11218 7052 11290
rect 7208 11218 7236 11834
rect 7300 11354 7328 14010
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11898 7512 12038
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 5264 10736 5316 10742
rect 6552 10736 6604 10742
rect 5264 10678 5316 10684
rect 5630 10704 5686 10713
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5276 9722 5304 10678
rect 6552 10678 6604 10684
rect 5630 10639 5686 10648
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4908 8906 4936 9386
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4908 8634 4936 8842
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5552 7954 5580 8910
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5000 6662 5028 7278
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5000 6186 5028 6598
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4724 4622 4752 4655
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3126 4200 3334
rect 4632 3194 4660 4558
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4724 3738 4752 4082
rect 4816 3942 4844 5102
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4724 3602 4752 3674
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4618 3088 4674 3097
rect 4618 3023 4674 3032
rect 3988 2746 4108 2774
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1964 1873 1992 2246
rect 1950 1864 2006 1873
rect 1950 1799 2006 1808
rect 2424 1737 2452 2382
rect 3068 2145 3096 2382
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3054 2136 3110 2145
rect 3054 2071 3110 2080
rect 3252 1834 3280 2246
rect 3896 2038 3924 2246
rect 3884 2032 3936 2038
rect 4080 2009 4108 2746
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 3023
rect 4816 2922 4844 3606
rect 4908 3466 4936 5850
rect 5000 5370 5028 6122
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4988 2440 5040 2446
rect 5092 2428 5120 7686
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5184 6118 5212 6802
rect 5460 6798 5488 7278
rect 5644 6866 5672 10639
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9178 6868 9454
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6840 8566 6868 9114
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5574 5212 6054
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5368 3670 5396 6734
rect 5460 6254 5488 6734
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5460 5846 5488 6190
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5460 5234 5488 5782
rect 5552 5370 5580 6666
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5736 6202 5764 6258
rect 5644 5710 5672 6190
rect 5736 6174 5856 6202
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5644 4826 5672 5646
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5736 3466 5764 6054
rect 5828 5234 5856 6174
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5814 4040 5870 4049
rect 5814 3975 5870 3984
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5040 2400 5120 2428
rect 4988 2382 5040 2388
rect 3884 1974 3936 1980
rect 4066 2000 4122 2009
rect 5092 1970 5120 2400
rect 5172 2440 5224 2446
rect 5276 2417 5304 3402
rect 5552 2990 5580 3402
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5828 2650 5856 3975
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5920 2446 5948 8298
rect 6196 2446 6224 8298
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 5914 6316 6258
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6380 3670 6408 5170
rect 6472 4842 6500 7346
rect 6552 6656 6604 6662
rect 6604 6616 6684 6644
rect 6552 6598 6604 6604
rect 6656 5234 6684 6616
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6748 5778 6776 6054
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6472 4814 6592 4842
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 3097 6316 3334
rect 6274 3088 6330 3097
rect 6472 3058 6500 4694
rect 6274 3023 6330 3032
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6564 2774 6592 4814
rect 6656 3466 6684 5170
rect 6932 4690 6960 11018
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7024 10130 7052 10610
rect 7208 10266 7236 11154
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10674 7604 10950
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7024 8498 7052 10066
rect 7668 9654 7696 14214
rect 7760 14074 7788 17750
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7852 17202 7880 17274
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7852 15570 7880 16934
rect 7944 16250 7972 20402
rect 8036 17814 8064 23054
rect 8128 22438 8156 28154
rect 8220 28082 8248 29990
rect 10428 29850 10456 30262
rect 10140 29844 10192 29850
rect 10140 29786 10192 29792
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 9588 29096 9640 29102
rect 9588 29038 9640 29044
rect 9128 28484 9180 28490
rect 9128 28426 9180 28432
rect 8944 28416 8996 28422
rect 8944 28358 8996 28364
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8220 26586 8248 27270
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 8220 25294 8248 26522
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 8220 22642 8248 22918
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 8864 21962 8892 23054
rect 8852 21956 8904 21962
rect 8852 21898 8904 21904
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8220 20466 8248 20742
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8128 19922 8156 20402
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8864 18358 8892 21898
rect 8956 20602 8984 28358
rect 9140 28082 9168 28426
rect 9600 28218 9628 29038
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9692 28694 9720 28902
rect 9680 28688 9732 28694
rect 9680 28630 9732 28636
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 9692 26994 9720 28630
rect 10152 28082 10180 29786
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10520 29034 10548 29582
rect 11348 29578 11376 30534
rect 11900 30394 11928 30738
rect 11980 30728 12032 30734
rect 11978 30696 11980 30705
rect 12032 30696 12034 30705
rect 11978 30631 12034 30640
rect 11888 30388 11940 30394
rect 11888 30330 11940 30336
rect 11992 29850 12020 30631
rect 12084 30258 12112 31282
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 11336 29572 11388 29578
rect 11336 29514 11388 29520
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 10508 29028 10560 29034
rect 10508 28970 10560 28976
rect 10520 28490 10548 28970
rect 11072 28490 11100 29446
rect 11796 29232 11848 29238
rect 12084 29186 12112 30194
rect 12162 29336 12218 29345
rect 12162 29271 12164 29280
rect 12216 29271 12218 29280
rect 12164 29242 12216 29248
rect 12256 29232 12308 29238
rect 11848 29180 11928 29186
rect 11796 29174 11928 29180
rect 11336 29164 11388 29170
rect 11808 29158 11928 29174
rect 12084 29170 12204 29186
rect 12256 29174 12308 29180
rect 11336 29106 11388 29112
rect 10508 28484 10560 28490
rect 10508 28426 10560 28432
rect 11060 28484 11112 28490
rect 11060 28426 11112 28432
rect 10324 28144 10376 28150
rect 10244 28104 10324 28132
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10244 28014 10272 28104
rect 10324 28086 10376 28092
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 10244 27130 10272 27950
rect 10324 27940 10376 27946
rect 10324 27882 10376 27888
rect 10336 27849 10364 27882
rect 10322 27840 10378 27849
rect 10322 27775 10378 27784
rect 10336 27606 10364 27775
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10140 27056 10192 27062
rect 10140 26998 10192 27004
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 9128 26852 9180 26858
rect 9128 26794 9180 26800
rect 9496 26852 9548 26858
rect 9496 26794 9548 26800
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 9140 19854 9168 26794
rect 9508 23118 9536 26794
rect 10152 26330 10180 26998
rect 10428 26790 10456 28018
rect 10520 27470 10548 28426
rect 11348 28422 11376 29106
rect 11900 28966 11928 29158
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 12084 29164 12216 29170
rect 12084 29158 12164 29164
rect 11888 28960 11940 28966
rect 11808 28920 11888 28948
rect 11808 28490 11836 28920
rect 11888 28902 11940 28908
rect 11796 28484 11848 28490
rect 11796 28426 11848 28432
rect 11336 28416 11388 28422
rect 11336 28358 11388 28364
rect 11152 28144 11204 28150
rect 11152 28086 11204 28092
rect 10782 27704 10838 27713
rect 10782 27639 10784 27648
rect 10836 27639 10838 27648
rect 10784 27610 10836 27616
rect 10508 27464 10560 27470
rect 10508 27406 10560 27412
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10416 26784 10468 26790
rect 10416 26726 10468 26732
rect 10152 26314 10456 26330
rect 10152 26308 10468 26314
rect 10152 26302 10416 26308
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9600 24206 9628 24550
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9600 23730 9628 24142
rect 10152 24138 10180 26302
rect 10416 26250 10468 26256
rect 10232 25764 10284 25770
rect 10232 25706 10284 25712
rect 10244 24206 10272 25706
rect 10520 25362 10548 27406
rect 10888 27130 10916 27406
rect 11164 27402 11192 28086
rect 11348 27674 11376 28358
rect 11808 28150 11836 28426
rect 11992 28200 12020 29106
rect 11900 28172 12020 28200
rect 11796 28144 11848 28150
rect 11796 28086 11848 28092
rect 11900 28014 11928 28172
rect 11888 28008 11940 28014
rect 11888 27950 11940 27956
rect 11336 27668 11388 27674
rect 11336 27610 11388 27616
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 11152 27396 11204 27402
rect 11152 27338 11204 27344
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10692 26988 10744 26994
rect 10612 26948 10692 26976
rect 10612 26382 10640 26948
rect 10692 26930 10744 26936
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10508 25356 10560 25362
rect 10508 25298 10560 25304
rect 10612 24206 10640 26318
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10704 25974 10732 26250
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 10152 23730 10180 24074
rect 10612 23730 10640 24142
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10152 23186 10180 23666
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10612 23118 10640 23666
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9324 22098 9352 22442
rect 9508 22166 9536 23054
rect 10612 22642 10640 23054
rect 11164 22642 11192 24006
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 22166 11008 22510
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9678 21992 9734 22001
rect 9678 21927 9734 21936
rect 9402 21856 9458 21865
rect 9402 21791 9458 21800
rect 9416 21690 9444 21791
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9496 21616 9548 21622
rect 9310 21584 9366 21593
rect 9366 21542 9444 21570
rect 9310 21519 9366 21528
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9310 21448 9366 21457
rect 9232 21350 9260 21422
rect 9310 21383 9366 21392
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9324 20942 9352 21383
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9220 20528 9272 20534
rect 9324 20516 9352 20878
rect 9416 20534 9444 21542
rect 9488 21564 9496 21604
rect 9488 21558 9548 21564
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9488 21468 9516 21558
rect 9488 21440 9536 21468
rect 9600 21457 9628 21558
rect 9272 20488 9352 20516
rect 9404 20528 9456 20534
rect 9220 20470 9272 20476
rect 9404 20470 9456 20476
rect 9508 20346 9536 21440
rect 9586 21448 9642 21457
rect 9586 21383 9642 21392
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9416 20318 9536 20346
rect 9416 20058 9444 20318
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9508 19854 9536 20198
rect 9600 20058 9628 21286
rect 9692 20874 9720 21927
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10244 20942 10272 21626
rect 10612 21593 10640 21626
rect 10598 21584 10654 21593
rect 10598 21519 10654 21528
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 8942 19408 8998 19417
rect 8942 19343 8998 19352
rect 8956 18970 8984 19343
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8128 17882 8156 18226
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7944 15706 7972 16186
rect 8036 16114 8064 16934
rect 8128 16794 8156 17206
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8116 16584 8168 16590
rect 8312 16572 8340 16934
rect 9140 16726 9168 19790
rect 9600 19446 9628 19994
rect 10048 19984 10100 19990
rect 10048 19926 10100 19932
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9600 18290 9628 19382
rect 10060 18698 10088 19926
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10244 19394 10272 20878
rect 10520 20398 10548 20878
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10520 19854 10548 20334
rect 10704 19990 10732 20946
rect 10692 19984 10744 19990
rect 10692 19926 10744 19932
rect 10508 19848 10560 19854
rect 10692 19848 10744 19854
rect 10508 19790 10560 19796
rect 10598 19816 10654 19825
rect 10152 19174 10180 19382
rect 10244 19378 10456 19394
rect 10244 19372 10468 19378
rect 10244 19366 10416 19372
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9232 17746 9260 18022
rect 9600 17746 9628 18226
rect 9692 18154 9720 18634
rect 10152 18426 10180 19110
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10244 18290 10272 19366
rect 10416 19314 10468 19320
rect 10520 18902 10548 19790
rect 10692 19790 10744 19796
rect 10968 19848 11020 19854
rect 11020 19808 11100 19836
rect 10968 19790 11020 19796
rect 10598 19751 10654 19760
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 18426 10364 18702
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9600 17202 9628 17682
rect 10060 17678 10088 18022
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9876 17542 9904 17614
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9416 16658 9444 16934
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 8116 16526 8168 16532
rect 8220 16544 8340 16572
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7852 12170 7880 15370
rect 8036 15094 8064 15438
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 8128 14618 8156 16526
rect 8220 15434 8248 16544
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8312 15026 8340 16390
rect 9692 16182 9720 16594
rect 9784 16590 9812 17478
rect 10060 16794 10088 17614
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9770 16280 9826 16289
rect 9770 16215 9772 16224
rect 9824 16215 9826 16224
rect 9772 16186 9824 16192
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 8390 16008 8446 16017
rect 8390 15943 8446 15952
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8404 14906 8432 15943
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8956 15502 8984 15846
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8220 14890 8432 14906
rect 8208 14884 8432 14890
rect 8260 14878 8432 14884
rect 8208 14826 8260 14832
rect 8956 14618 8984 15302
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8036 13530 8064 13874
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12374 7972 13262
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8036 12986 8064 13194
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7668 8401 7696 9590
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7654 8392 7710 8401
rect 7654 8327 7710 8336
rect 7852 8242 7880 12106
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 11150 7972 11494
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8036 10130 8064 12922
rect 8128 12850 8156 14554
rect 8956 14414 8984 14554
rect 9140 14414 9168 15370
rect 9324 14414 9352 15438
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8312 14006 8340 14282
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8312 13394 8340 13942
rect 9140 13938 9168 14350
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8312 12918 8340 13194
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8208 12436 8260 12442
rect 8312 12434 8340 12854
rect 8404 12850 8432 13194
rect 8772 12850 8800 13670
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 9416 12434 9444 15642
rect 9496 15632 9548 15638
rect 9494 15600 9496 15609
rect 9548 15600 9550 15609
rect 9494 15535 9550 15544
rect 9692 14346 9720 16118
rect 10336 16114 10364 16662
rect 10612 16590 10640 19751
rect 10704 19310 10732 19790
rect 11072 19514 11100 19808
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 17678 10916 18566
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10336 15026 10364 16050
rect 10428 15162 10456 16050
rect 10508 15972 10560 15978
rect 10508 15914 10560 15920
rect 10520 15162 10548 15914
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9692 12918 9720 14282
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 8312 12406 8432 12434
rect 8208 12378 8260 12384
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10810 8156 11086
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8220 8838 8248 12378
rect 8404 11082 8432 12406
rect 9232 12406 9444 12434
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8634 8248 8774
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7760 8214 7880 8242
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7546 7420 7822
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7760 7410 7788 8214
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7546 7880 7686
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7944 7426 7972 8502
rect 8312 7698 8340 9930
rect 8772 9654 8800 11018
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8956 10130 8984 10678
rect 9048 10470 9076 11698
rect 9140 11558 9168 11698
rect 9232 11626 9260 12406
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9600 11830 9628 12310
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9324 11694 9352 11766
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9586 11656 9642 11665
rect 9220 11620 9272 11626
rect 9692 11626 9720 11698
rect 9586 11591 9642 11600
rect 9680 11620 9732 11626
rect 9220 11562 9272 11568
rect 9600 11558 9628 11591
rect 9680 11562 9732 11568
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9692 11150 9720 11290
rect 9784 11218 9812 14962
rect 10520 14550 10548 15098
rect 10612 15008 10640 16526
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10980 16250 11008 16458
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10692 15020 10744 15026
rect 10612 14980 10692 15008
rect 10692 14962 10744 14968
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10796 13938 10824 14418
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 9876 13190 9904 13874
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9876 12986 9904 13126
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 10152 12434 10180 13262
rect 10612 12646 10640 13874
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10152 12406 10272 12434
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9508 10810 9536 11086
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8772 9042 8800 9590
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8864 8974 8892 9318
rect 8956 9042 8984 10066
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 9140 8838 9168 9522
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9600 8566 9628 9862
rect 9692 9382 9720 10610
rect 9784 9586 9812 11154
rect 9876 11082 9904 12106
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9692 8498 9720 9318
rect 9784 8906 9812 9522
rect 9876 9194 9904 11018
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10060 10062 10088 10950
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9382 9996 9522
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9876 9166 9996 9194
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7852 7398 7972 7426
rect 8128 7670 8340 7698
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7024 4486 7052 5510
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6734 3768 6790 3777
rect 6734 3703 6736 3712
rect 6788 3703 6790 3712
rect 6736 3674 6788 3680
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6840 3233 6868 3878
rect 7116 3602 7144 5646
rect 7208 4146 7236 7278
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 5030 7512 6598
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7392 3738 7420 4966
rect 7576 4146 7604 6326
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7760 4146 7788 4218
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7852 4026 7880 7398
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7944 4146 7972 5782
rect 8036 5234 8064 6122
rect 8128 5914 8156 7670
rect 8298 7576 8354 7585
rect 8298 7511 8354 7520
rect 8312 7478 8340 7511
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8128 4622 8156 5170
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4146 8156 4422
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7748 4004 7800 4010
rect 7852 3998 8064 4026
rect 7748 3946 7800 3952
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7562 3632 7618 3641
rect 7104 3596 7156 3602
rect 7760 3602 7788 3946
rect 7562 3567 7618 3576
rect 7656 3596 7708 3602
rect 7104 3538 7156 3544
rect 7576 3534 7604 3567
rect 7656 3538 7708 3544
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 6826 3224 6882 3233
rect 7208 3194 7236 3334
rect 7668 3194 7696 3538
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 3194 7880 3402
rect 6826 3159 6882 3168
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 6564 2746 6684 2774
rect 6656 2650 6684 2746
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 8036 2446 8064 3998
rect 8220 3942 8248 6734
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8312 6118 8340 6598
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5846 8340 5877
rect 8300 5840 8352 5846
rect 8298 5808 8300 5817
rect 8352 5808 8354 5817
rect 8298 5743 8354 5752
rect 8312 5710 8340 5743
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8220 2774 8248 3470
rect 8312 3058 8340 5510
rect 8496 3058 8524 6598
rect 8956 5710 8984 7686
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8680 5370 8708 5578
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8864 4690 8892 5034
rect 8956 5030 8984 5646
rect 9048 5370 9076 8298
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 6322 9168 6598
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5642 9168 6258
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8942 4448 8998 4457
rect 8772 4214 8800 4422
rect 8942 4383 8998 4392
rect 8850 4312 8906 4321
rect 8956 4282 8984 4383
rect 8850 4247 8852 4256
rect 8904 4247 8906 4256
rect 8944 4276 8996 4282
rect 8852 4218 8904 4224
rect 8944 4218 8996 4224
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8772 4078 8800 4150
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8864 3369 8892 4218
rect 8956 3777 8984 4218
rect 8942 3768 8998 3777
rect 8942 3703 8998 3712
rect 8850 3360 8906 3369
rect 8850 3295 8906 3304
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8220 2746 8340 2774
rect 8312 2650 8340 2746
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 5632 2440 5684 2446
rect 5172 2382 5224 2388
rect 5262 2408 5318 2417
rect 5184 2281 5212 2382
rect 5632 2382 5684 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 5262 2343 5318 2352
rect 5170 2272 5226 2281
rect 5170 2207 5226 2216
rect 4066 1935 4122 1944
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 5644 1902 5672 2382
rect 6656 2106 6684 2382
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 3240 1828 3292 1834
rect 3240 1770 3292 1776
rect 2410 1728 2466 1737
rect 8128 1698 8156 2518
rect 8404 2446 8432 2790
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 2410 1663 2466 1672
rect 8116 1692 8168 1698
rect 8116 1634 8168 1640
rect 9048 1601 9076 5306
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9140 3505 9168 4014
rect 9232 3534 9260 8298
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9324 6866 9352 7482
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9324 5710 9352 6394
rect 9692 6322 9720 6734
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9416 5778 9444 6190
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 5370 9352 5646
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9310 5264 9366 5273
rect 9784 5234 9812 6802
rect 9310 5199 9366 5208
rect 9772 5228 9824 5234
rect 9324 5166 9352 5199
rect 9772 5170 9824 5176
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9324 3602 9352 5102
rect 9968 4826 9996 9166
rect 10060 7002 10088 9318
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10152 7546 10180 8502
rect 10244 7886 10272 12406
rect 10796 12238 10824 13874
rect 10888 13841 10916 14010
rect 10874 13832 10930 13841
rect 10874 13767 10930 13776
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 11286 10364 11698
rect 10600 11552 10652 11558
rect 10598 11520 10600 11529
rect 10652 11520 10654 11529
rect 10598 11455 10654 11464
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10888 9654 10916 13670
rect 10980 13326 11008 14962
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11072 12918 11100 13194
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10980 11762 11008 12174
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10980 11354 11008 11698
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11072 11150 11100 12854
rect 11256 12646 11284 27542
rect 11348 18970 11376 27610
rect 11900 27470 11928 27950
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11900 26858 11928 27406
rect 12084 27334 12112 29158
rect 12164 29106 12216 29112
rect 12268 29034 12296 29174
rect 12256 29028 12308 29034
rect 12256 28970 12308 28976
rect 12452 28694 12480 30194
rect 12636 30054 12664 31282
rect 12912 30190 12940 31282
rect 13280 30870 13308 31300
rect 13544 31136 13596 31142
rect 13544 31078 13596 31084
rect 13268 30864 13320 30870
rect 13268 30806 13320 30812
rect 12900 30184 12952 30190
rect 12900 30126 12952 30132
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12440 28688 12492 28694
rect 12440 28630 12492 28636
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12164 28144 12216 28150
rect 12164 28086 12216 28092
rect 12176 27713 12204 28086
rect 12256 27872 12308 27878
rect 12544 27849 12572 28494
rect 12256 27814 12308 27820
rect 12530 27840 12586 27849
rect 12162 27704 12218 27713
rect 12162 27639 12218 27648
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 12164 26580 12216 26586
rect 12164 26522 12216 26528
rect 11888 26512 11940 26518
rect 11888 26454 11940 26460
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11532 23050 11560 24006
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 11532 22094 11560 22986
rect 11440 22066 11560 22094
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11348 16250 11376 18906
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 15706 11376 16186
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11440 13530 11468 22066
rect 11624 22030 11652 23462
rect 11716 22030 11744 25298
rect 11900 23730 11928 26454
rect 12176 24818 12204 26522
rect 12268 25430 12296 27814
rect 12530 27775 12586 27784
rect 12636 26518 12664 29990
rect 12912 29646 12940 30126
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12728 29306 12756 29582
rect 12716 29300 12768 29306
rect 12716 29242 12768 29248
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12728 28082 12756 28494
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12820 27713 12848 28358
rect 12806 27704 12862 27713
rect 12806 27639 12862 27648
rect 12912 27554 12940 29582
rect 13280 29578 13308 30806
rect 13556 30326 13584 31078
rect 15120 30938 15148 31690
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15108 30932 15160 30938
rect 15108 30874 15160 30880
rect 15120 30734 15148 30874
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 14924 30592 14976 30598
rect 14924 30534 14976 30540
rect 13544 30320 13596 30326
rect 13544 30262 13596 30268
rect 14004 30184 14056 30190
rect 14004 30126 14056 30132
rect 14016 29714 14044 30126
rect 14004 29708 14056 29714
rect 14004 29650 14056 29656
rect 13268 29572 13320 29578
rect 13268 29514 13320 29520
rect 13280 28082 13308 29514
rect 14016 29238 14044 29650
rect 14004 29232 14056 29238
rect 14004 29174 14056 29180
rect 14936 29170 14964 30534
rect 15212 29306 15240 31282
rect 15304 30598 15332 31350
rect 17420 31346 17448 31622
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 17776 31408 17828 31414
rect 17776 31350 17828 31356
rect 16672 31340 16724 31346
rect 16672 31282 16724 31288
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17408 31340 17460 31346
rect 17408 31282 17460 31288
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 16580 31204 16632 31210
rect 16580 31146 16632 31152
rect 15384 31136 15436 31142
rect 15384 31078 15436 31084
rect 15396 30734 15424 31078
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15292 30592 15344 30598
rect 15292 30534 15344 30540
rect 15304 30258 15332 30534
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15304 29238 15332 30194
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 14924 29164 14976 29170
rect 14924 29106 14976 29112
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 14648 28688 14700 28694
rect 14648 28630 14700 28636
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 14096 28008 14148 28014
rect 14096 27950 14148 27956
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 12820 27526 12940 27554
rect 12820 26586 12848 27526
rect 13004 27470 13032 27814
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12912 26790 12940 27338
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 12624 26512 12676 26518
rect 12624 26454 12676 26460
rect 12820 26382 12848 26522
rect 12912 26382 12940 26726
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12452 26042 12480 26182
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12544 25838 12572 26318
rect 12624 26240 12676 26246
rect 13004 26194 13032 27406
rect 14108 27334 14136 27950
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14108 26994 14136 27270
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 12624 26182 12676 26188
rect 12636 25906 12664 26182
rect 12912 26166 13032 26194
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12256 25424 12308 25430
rect 12256 25366 12308 25372
rect 12636 25226 12664 25842
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 11992 24410 12020 24754
rect 12176 24698 12204 24754
rect 12360 24750 12388 25162
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12084 24670 12204 24698
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 12084 23322 12112 24670
rect 12452 24206 12480 25094
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12164 23588 12216 23594
rect 12164 23530 12216 23536
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 12176 22710 12204 23530
rect 12164 22704 12216 22710
rect 12084 22664 12164 22692
rect 12084 22166 12112 22664
rect 12164 22646 12216 22652
rect 12360 22642 12388 23666
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11532 20942 11560 21490
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11716 20534 11744 20742
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 11992 20330 12020 21898
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11532 19514 11560 20198
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11716 17882 11744 18838
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 11624 14958 11652 16390
rect 11716 15162 11744 16730
rect 11808 15502 11836 19450
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11992 18086 12020 18294
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 17882 12020 18022
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14550 11560 14758
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11532 13394 11560 13942
rect 11624 13938 11652 14894
rect 11716 14278 11744 14894
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11532 12442 11560 13330
rect 11716 13326 11744 13874
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11716 12918 11744 13262
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11532 11830 11560 12378
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11060 11144 11112 11150
rect 11058 11112 11060 11121
rect 11112 11112 11114 11121
rect 11058 11047 11114 11056
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10888 8838 10916 9590
rect 11072 9586 11100 10610
rect 11348 10606 11376 11698
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11348 10266 11376 10542
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 9178 11100 9522
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10152 7410 10180 7482
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10244 6866 10272 7822
rect 10612 7410 10640 8230
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10416 6928 10468 6934
rect 10468 6888 10548 6916
rect 10416 6870 10468 6876
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6390 10088 6734
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10428 6202 10456 6258
rect 10336 6174 10456 6202
rect 10232 6112 10284 6118
rect 10336 6066 10364 6174
rect 10284 6060 10364 6066
rect 10232 6054 10364 6060
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10244 6038 10364 6054
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9600 4010 9628 4626
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 4321 9720 4558
rect 9678 4312 9734 4321
rect 9678 4247 9734 4256
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9876 4146 9904 4218
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9680 4072 9732 4078
rect 9732 4032 9812 4060
rect 9680 4014 9732 4020
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9220 3528 9272 3534
rect 9126 3496 9182 3505
rect 9220 3470 9272 3476
rect 9126 3431 9182 3440
rect 9692 3398 9720 3606
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 1766 9720 2382
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 9784 1630 9812 4032
rect 9956 3664 10008 3670
rect 10060 3641 10088 5102
rect 10152 4049 10180 5170
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10138 4040 10194 4049
rect 10138 3975 10194 3984
rect 9956 3606 10008 3612
rect 10046 3632 10102 3641
rect 9968 3534 9996 3606
rect 10046 3567 10102 3576
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10060 1698 10088 3567
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10048 1692 10100 1698
rect 10048 1634 10100 1640
rect 9772 1624 9824 1630
rect 9034 1592 9090 1601
rect 9772 1566 9824 1572
rect 9034 1527 9090 1536
rect 10152 1426 10180 3334
rect 10244 3126 10272 4966
rect 10336 3534 10364 6038
rect 10428 5778 10456 6054
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10520 4865 10548 6888
rect 10506 4856 10562 4865
rect 10416 4820 10468 4826
rect 10506 4791 10562 4800
rect 10416 4762 10468 4768
rect 10428 4593 10456 4762
rect 10520 4690 10548 4791
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10414 4584 10470 4593
rect 10414 4519 10470 4528
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10428 3398 10456 4218
rect 10508 4208 10560 4214
rect 10506 4176 10508 4185
rect 10560 4176 10562 4185
rect 10612 4146 10640 7346
rect 10692 6792 10744 6798
rect 10690 6760 10692 6769
rect 10744 6760 10746 6769
rect 10690 6695 10746 6704
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10704 4282 10732 5510
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10506 4111 10562 4120
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10598 3904 10654 3913
rect 10598 3839 10654 3848
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10506 3088 10562 3097
rect 10506 3023 10562 3032
rect 10414 2816 10470 2825
rect 10414 2751 10470 2760
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 1494 10364 2246
rect 10324 1488 10376 1494
rect 10324 1430 10376 1436
rect 10428 1442 10456 2751
rect 10520 2446 10548 3023
rect 10612 2990 10640 3839
rect 10690 3768 10746 3777
rect 10690 3703 10746 3712
rect 10704 3466 10732 3703
rect 10796 3466 10824 7686
rect 10888 6474 10916 7754
rect 10980 7002 11008 8298
rect 11072 8294 11100 8774
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11072 7585 11100 7890
rect 11164 7818 11192 8230
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11058 7576 11114 7585
rect 11058 7511 11114 7520
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10966 6896 11022 6905
rect 11164 6866 11192 7754
rect 10966 6831 11022 6840
rect 11152 6860 11204 6866
rect 10980 6662 11008 6831
rect 11152 6802 11204 6808
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 10888 6446 11008 6474
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10888 5302 10916 5782
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10888 4282 10916 4626
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10874 3496 10930 3505
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10784 3460 10836 3466
rect 10874 3431 10930 3440
rect 10784 3402 10836 3408
rect 10600 2984 10652 2990
rect 10598 2952 10600 2961
rect 10652 2952 10654 2961
rect 10598 2887 10654 2896
rect 10888 2825 10916 3431
rect 10874 2816 10930 2825
rect 10874 2751 10930 2760
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10692 1624 10744 1630
rect 10692 1566 10744 1572
rect 10140 1420 10192 1426
rect 10428 1414 10640 1442
rect 10140 1362 10192 1368
rect 10612 800 10640 1414
rect 10704 800 10732 1566
rect 10796 800 10824 2518
rect 10876 1420 10928 1426
rect 10876 1362 10928 1368
rect 10888 800 10916 1362
rect 10980 800 11008 6446
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5846 11100 6122
rect 11164 6118 11192 6598
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11164 4622 11192 6054
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11256 3534 11284 8842
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11348 4690 11376 6870
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11440 6322 11468 6598
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11532 5896 11560 7142
rect 11440 5868 11560 5896
rect 11440 4690 11468 5868
rect 11624 5828 11652 12106
rect 11716 11830 11744 12854
rect 11808 12850 11836 14486
rect 11900 14006 11928 16934
rect 12084 16182 12112 18226
rect 12176 17882 12204 20878
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12084 14414 12112 16118
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11992 13308 12020 13874
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11900 13280 12020 13308
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11900 12782 11928 13280
rect 12084 12918 12112 13398
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11900 12238 11928 12718
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11716 10742 11744 11766
rect 11900 11694 11928 12174
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11716 9654 11744 10678
rect 11900 10674 11928 11630
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11808 9722 11836 10610
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11900 9586 11928 10610
rect 12070 10568 12126 10577
rect 12070 10503 12072 10512
rect 12124 10503 12126 10512
rect 12072 10474 12124 10480
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8022 11928 8774
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 11900 7886 11928 7958
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11624 5800 11836 5828
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11532 5302 11560 5714
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11624 5302 11652 5578
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11624 5030 11652 5238
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11610 4720 11666 4729
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11428 4684 11480 4690
rect 11610 4655 11666 4664
rect 11428 4626 11480 4632
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11440 4282 11468 4490
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11256 2774 11284 3470
rect 11624 3398 11652 4655
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11164 2746 11284 2774
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 11072 800 11100 2314
rect 11164 800 11192 2746
rect 11242 2680 11298 2689
rect 11242 2615 11244 2624
rect 11296 2615 11298 2624
rect 11244 2586 11296 2592
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 11256 800 11284 2042
rect 11348 800 11376 3334
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11440 800 11468 3130
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11532 800 11560 2382
rect 11624 800 11652 3062
rect 11716 800 11744 4422
rect 11808 4049 11836 5800
rect 11900 4690 11928 6326
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5030 12020 6054
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11980 4752 12032 4758
rect 11978 4720 11980 4729
rect 12032 4720 12034 4729
rect 11888 4684 11940 4690
rect 11978 4655 12034 4664
rect 11888 4626 11940 4632
rect 11900 4214 11928 4626
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11794 4040 11850 4049
rect 11794 3975 11850 3984
rect 11808 3942 11836 3975
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11900 3534 11928 4150
rect 11992 4078 12020 4558
rect 12084 4282 12112 5578
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 2774 11836 3334
rect 11900 2922 11928 3470
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11992 2854 12020 4014
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11808 2746 11928 2774
rect 11900 800 11928 2746
rect 11992 2446 12020 2790
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 11992 800 12020 1974
rect 12084 800 12112 3538
rect 12176 3194 12204 12922
rect 12268 10538 12296 22102
rect 12360 22030 12388 22578
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12452 18766 12480 24142
rect 12636 24138 12664 25162
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12532 23520 12584 23526
rect 12530 23488 12532 23497
rect 12584 23488 12586 23497
rect 12530 23423 12586 23432
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12544 21350 12572 22102
rect 12912 22094 12940 26166
rect 13096 26042 13124 26454
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 13004 23186 13032 25774
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13648 25106 13676 26862
rect 13924 26314 13952 26862
rect 14016 26382 14044 26930
rect 14108 26586 14136 26930
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14004 26376 14056 26382
rect 14004 26318 14056 26324
rect 13912 26308 13964 26314
rect 13912 26250 13964 26256
rect 13820 25152 13872 25158
rect 13648 25100 13820 25106
rect 13648 25094 13872 25100
rect 13464 24886 13492 25094
rect 13648 25078 13860 25094
rect 13452 24880 13504 24886
rect 13452 24822 13504 24828
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13372 24206 13400 24686
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 12992 23180 13044 23186
rect 13044 23140 13124 23168
rect 12992 23122 13044 23128
rect 12912 22066 13032 22094
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12728 19514 12756 19994
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12622 18864 12678 18873
rect 12622 18799 12678 18808
rect 12636 18766 12664 18799
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12728 17678 12756 18226
rect 12820 18154 12848 19178
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12622 17232 12678 17241
rect 12622 17167 12678 17176
rect 12636 16114 12664 17167
rect 12728 16658 12756 17614
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12820 16590 12848 18090
rect 12912 17270 12940 20946
rect 13004 20942 13032 22066
rect 13096 21622 13124 23140
rect 13188 22710 13216 24074
rect 13372 23730 13400 24142
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 13280 22438 13308 22918
rect 13372 22710 13400 22918
rect 13464 22710 13492 24822
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13556 22778 13584 23666
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 13452 22704 13504 22710
rect 13452 22646 13504 22652
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13096 20856 13124 21558
rect 13268 21548 13320 21554
rect 13372 21536 13400 22646
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13464 21894 13492 21966
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13320 21508 13400 21536
rect 13544 21548 13596 21554
rect 13268 21490 13320 21496
rect 13544 21490 13596 21496
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13176 20868 13228 20874
rect 13096 20828 13176 20856
rect 13096 18698 13124 20828
rect 13176 20810 13228 20816
rect 13280 20618 13308 21286
rect 13464 21146 13492 21354
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13452 20936 13504 20942
rect 13556 20924 13584 21490
rect 13504 20896 13584 20924
rect 13452 20878 13504 20884
rect 13464 20618 13492 20878
rect 13280 20590 13492 20618
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15094 12480 15846
rect 12636 15366 12664 16050
rect 13004 16046 13032 17614
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12544 14346 12572 14826
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12636 14226 12664 15302
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12912 14482 12940 15030
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 13004 14385 13032 14486
rect 12990 14376 13046 14385
rect 12990 14311 13046 14320
rect 12544 14198 12664 14226
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12346 12744 12402 12753
rect 12346 12679 12348 12688
rect 12400 12679 12402 12688
rect 12348 12650 12400 12656
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11694 12480 12038
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12544 10810 12572 14198
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12268 7750 12296 8434
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12452 6934 12480 10610
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12544 8634 12572 9522
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12544 7886 12572 8570
rect 12636 8430 12664 13670
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12728 7886 12756 14214
rect 13004 13938 13032 14311
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12808 13728 12860 13734
rect 12806 13696 12808 13705
rect 12860 13696 12862 13705
rect 12806 13631 12862 13640
rect 12912 13433 12940 13806
rect 12898 13424 12954 13433
rect 13096 13394 13124 18634
rect 13188 17202 13216 20198
rect 13372 18766 13400 20590
rect 13450 19544 13506 19553
rect 13450 19479 13452 19488
rect 13504 19479 13506 19488
rect 13452 19450 13504 19456
rect 13464 19378 13492 19450
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16794 13308 17138
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 12898 13359 12954 13368
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13372 12986 13400 18702
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13464 16726 13492 17546
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13464 15994 13492 16662
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13556 16114 13584 16526
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13464 15966 13584 15994
rect 13450 15464 13506 15473
rect 13450 15399 13452 15408
rect 13504 15399 13506 15408
rect 13452 15370 13504 15376
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12442 13032 12582
rect 13082 12472 13138 12481
rect 12992 12436 13044 12442
rect 13082 12407 13138 12416
rect 12992 12378 13044 12384
rect 13096 12306 13124 12407
rect 13174 12336 13230 12345
rect 13084 12300 13136 12306
rect 13174 12271 13230 12280
rect 13084 12242 13136 12248
rect 13188 12238 13216 12271
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 9586 12940 12038
rect 13188 11354 13216 12174
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13280 11218 13308 12786
rect 13556 12442 13584 15966
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13372 11082 13400 11698
rect 13556 11354 13584 12378
rect 13648 11898 13676 25078
rect 13924 24954 13952 26250
rect 14016 25906 14044 26318
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 14004 25764 14056 25770
rect 14004 25706 14056 25712
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13740 24410 13768 24754
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13924 24138 13952 24890
rect 13912 24132 13964 24138
rect 13912 24074 13964 24080
rect 13924 23798 13952 24074
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 20058 13768 21286
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13832 19990 13860 20810
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13726 19816 13782 19825
rect 13726 19751 13728 19760
rect 13780 19751 13782 19760
rect 13728 19722 13780 19728
rect 13832 19718 13860 19926
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13740 18290 13768 18566
rect 13832 18426 13860 19654
rect 13924 19378 13952 20742
rect 14016 19378 14044 25706
rect 14200 24750 14228 27406
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14384 24206 14412 25094
rect 14476 24614 14504 25230
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14476 23254 14504 24550
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14568 23322 14596 24278
rect 14660 23866 14688 28630
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14752 27674 14780 28018
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 15028 26382 15056 28902
rect 15304 28558 15332 29174
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15304 28218 15332 28494
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15488 27946 15516 31146
rect 16592 30802 16620 31146
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16212 30728 16264 30734
rect 16212 30670 16264 30676
rect 16396 30728 16448 30734
rect 16396 30670 16448 30676
rect 16224 30394 16252 30670
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 16408 30054 16436 30670
rect 16396 30048 16448 30054
rect 16396 29990 16448 29996
rect 16212 29572 16264 29578
rect 16212 29514 16264 29520
rect 15568 29504 15620 29510
rect 15568 29446 15620 29452
rect 15580 28490 15608 29446
rect 16224 28762 16252 29514
rect 16212 28756 16264 28762
rect 16212 28698 16264 28704
rect 16592 28558 16620 30738
rect 16684 30666 16712 31282
rect 17236 30938 17264 31282
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17420 30870 17448 31282
rect 17788 31210 17816 31350
rect 20548 31346 20576 31690
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 22744 31408 22796 31414
rect 22744 31350 22796 31356
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20904 31340 20956 31346
rect 20904 31282 20956 31288
rect 17776 31204 17828 31210
rect 17776 31146 17828 31152
rect 17408 30864 17460 30870
rect 17460 30824 17540 30852
rect 17408 30806 17460 30812
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 17224 30660 17276 30666
rect 17224 30602 17276 30608
rect 17236 30546 17264 30602
rect 17144 30518 17264 30546
rect 17144 30054 17172 30518
rect 17316 30320 17368 30326
rect 17316 30262 17368 30268
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 15568 28484 15620 28490
rect 15568 28426 15620 28432
rect 15476 27940 15528 27946
rect 15476 27882 15528 27888
rect 15580 27538 15608 28426
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15568 27532 15620 27538
rect 15568 27474 15620 27480
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 15212 26790 15240 27406
rect 15948 26994 15976 28018
rect 16592 28014 16620 28494
rect 16684 28422 16712 29446
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16580 28008 16632 28014
rect 16580 27950 16632 27956
rect 16592 27538 16620 27950
rect 16580 27532 16632 27538
rect 16580 27474 16632 27480
rect 16304 27464 16356 27470
rect 16304 27406 16356 27412
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 14936 25888 14964 26318
rect 15948 26042 15976 26930
rect 16316 26926 16344 27406
rect 16580 27396 16632 27402
rect 16580 27338 16632 27344
rect 16592 27130 16620 27338
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16304 26920 16356 26926
rect 16304 26862 16356 26868
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 16040 25974 16068 26726
rect 16316 26246 16344 26862
rect 16776 26382 16804 29786
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 16028 25968 16080 25974
rect 16028 25910 16080 25916
rect 15016 25900 15068 25906
rect 14936 25860 15016 25888
rect 15016 25842 15068 25848
rect 14832 25832 14884 25838
rect 14832 25774 14884 25780
rect 14844 25226 14872 25774
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14844 24410 14872 24754
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14936 24410 14964 24686
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14464 23248 14516 23254
rect 14464 23190 14516 23196
rect 14188 22160 14240 22166
rect 14188 22102 14240 22108
rect 14200 21078 14228 22102
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 14200 20602 14228 21014
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14384 19378 14412 21898
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14476 21146 14504 21422
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13924 16114 13952 18770
rect 14016 18290 14044 19178
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13372 10674 13400 11018
rect 13648 10742 13676 11834
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 9586 13216 9862
rect 13464 9722 13492 9930
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12544 7410 12572 7686
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12544 7002 12572 7346
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12544 6769 12572 6938
rect 12624 6792 12676 6798
rect 12530 6760 12586 6769
rect 12624 6734 12676 6740
rect 12530 6695 12586 6704
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12268 4690 12296 6394
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12360 5098 12388 5238
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12346 4856 12402 4865
rect 12346 4791 12402 4800
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12268 4010 12296 4626
rect 12360 4554 12388 4791
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12348 4276 12400 4282
rect 12400 4236 12480 4264
rect 12348 4218 12400 4224
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12268 3058 12296 3946
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12176 2514 12204 2926
rect 12256 2916 12308 2922
rect 12256 2858 12308 2864
rect 12268 2650 12296 2858
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12176 1034 12204 2314
rect 12360 1154 12388 4082
rect 12452 3058 12480 4236
rect 12544 3670 12572 5782
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 2582 12480 2994
rect 12544 2922 12572 3606
rect 12636 3466 12664 6734
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 5846 12756 6598
rect 12912 6322 12940 7482
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12820 5166 12848 5510
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12912 4826 12940 5170
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12714 3904 12770 3913
rect 12714 3839 12770 3848
rect 12728 3602 12756 3839
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12636 3126 12664 3402
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12636 1834 12664 3062
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 12624 1828 12676 1834
rect 12624 1770 12676 1776
rect 12622 1728 12678 1737
rect 12622 1663 12678 1672
rect 12440 1420 12492 1426
rect 12440 1362 12492 1368
rect 12348 1148 12400 1154
rect 12348 1090 12400 1096
rect 12176 1006 12388 1034
rect 12256 944 12308 950
rect 12256 886 12308 892
rect 12268 800 12296 886
rect 12360 800 12388 1006
rect 12452 800 12480 1362
rect 12636 800 12664 1663
rect 12728 1426 12756 1838
rect 12912 1442 12940 3946
rect 13004 2446 13032 8774
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13096 7886 13124 8230
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13096 3738 13124 7822
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13188 6798 13216 7346
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 5642 13216 6734
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13280 5234 13308 5646
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13188 4729 13216 5102
rect 13174 4720 13230 4729
rect 13174 4655 13230 4664
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13082 3632 13138 3641
rect 13082 3567 13138 3576
rect 13096 3398 13124 3567
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13188 2836 13216 4655
rect 13280 4282 13308 5170
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13268 3936 13320 3942
rect 13266 3904 13268 3913
rect 13320 3904 13322 3913
rect 13266 3839 13322 3848
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13280 2961 13308 3470
rect 13266 2952 13322 2961
rect 13266 2887 13322 2896
rect 13188 2808 13308 2836
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13096 2009 13124 2382
rect 13174 2136 13230 2145
rect 13174 2071 13230 2080
rect 13082 2000 13138 2009
rect 13082 1935 13138 1944
rect 12716 1420 12768 1426
rect 12912 1414 13124 1442
rect 12716 1362 12768 1368
rect 12900 1352 12952 1358
rect 12900 1294 12952 1300
rect 12992 1352 13044 1358
rect 12992 1294 13044 1300
rect 12716 1284 12768 1290
rect 12716 1226 12768 1232
rect 12728 800 12756 1226
rect 12808 1216 12860 1222
rect 12808 1158 12860 1164
rect 12820 800 12848 1158
rect 12912 800 12940 1294
rect 13004 800 13032 1294
rect 13096 800 13124 1414
rect 13188 800 13216 2071
rect 13280 800 13308 2808
rect 13372 800 13400 4422
rect 13464 4146 13492 8774
rect 13556 7818 13584 9454
rect 13740 9178 13768 15914
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13556 7342 13584 7754
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13556 5302 13584 5782
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13556 5166 13584 5238
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 4758 13584 5102
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13648 4622 13676 8230
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13452 4140 13504 4146
rect 13504 4100 13584 4128
rect 13452 4082 13504 4088
rect 13450 2952 13506 2961
rect 13450 2887 13452 2896
rect 13504 2887 13506 2896
rect 13452 2858 13504 2864
rect 13450 2816 13506 2825
rect 13450 2751 13506 2760
rect 13464 800 13492 2751
rect 13556 800 13584 4100
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13648 800 13676 3878
rect 13740 3641 13768 5850
rect 13832 4457 13860 6190
rect 13818 4448 13874 4457
rect 13818 4383 13874 4392
rect 13924 3913 13952 13874
rect 14016 13394 14044 18226
rect 14108 18086 14136 18226
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14200 15706 14228 19178
rect 14384 18290 14412 19314
rect 14660 19310 14688 21966
rect 15028 21962 15056 25842
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16224 25294 16252 25638
rect 16316 25294 16344 26182
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16408 25106 16436 25638
rect 16316 25078 16436 25106
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15212 23866 15240 24142
rect 15200 23860 15252 23866
rect 15200 23802 15252 23808
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 15212 23610 15240 23802
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15212 23582 15424 23610
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23118 15240 23462
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15212 21554 15240 21626
rect 15396 21554 15424 23582
rect 15488 22642 15516 23666
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15488 21962 15516 22034
rect 15948 22030 15976 22374
rect 16040 22030 16068 23802
rect 16132 23662 16160 24686
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16132 23526 16160 23598
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 16132 23186 16160 23462
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 16316 22574 16344 25078
rect 16500 24342 16528 26250
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16684 25498 16712 25842
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16776 25226 16804 26318
rect 16856 25968 16908 25974
rect 16856 25910 16908 25916
rect 16868 25294 16896 25910
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16488 24336 16540 24342
rect 16488 24278 16540 24284
rect 16776 23730 16804 25162
rect 16868 24818 16896 25230
rect 16960 24886 16988 28358
rect 17144 28150 17172 29990
rect 17328 29850 17356 30262
rect 17316 29844 17368 29850
rect 17316 29786 17368 29792
rect 17316 29164 17368 29170
rect 17316 29106 17368 29112
rect 17328 28694 17356 29106
rect 17408 28960 17460 28966
rect 17408 28902 17460 28908
rect 17316 28688 17368 28694
rect 17316 28630 17368 28636
rect 17132 28144 17184 28150
rect 17132 28086 17184 28092
rect 17420 28082 17448 28902
rect 17408 28076 17460 28082
rect 17408 28018 17460 28024
rect 17512 27674 17540 30824
rect 17788 30122 17816 31146
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 20260 31136 20312 31142
rect 20260 31078 20312 31084
rect 18064 30326 18092 31078
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 18052 30320 18104 30326
rect 18052 30262 18104 30268
rect 17776 30116 17828 30122
rect 17776 30058 17828 30064
rect 17592 29504 17644 29510
rect 17592 29446 17644 29452
rect 17604 29306 17632 29446
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17500 27668 17552 27674
rect 17500 27610 17552 27616
rect 17788 27538 17816 30058
rect 18340 29850 18368 30534
rect 18328 29844 18380 29850
rect 18328 29786 18380 29792
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 18064 28558 18092 29582
rect 18432 29578 18460 30738
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 20272 30326 20300 31078
rect 20732 30938 20760 31282
rect 20720 30932 20772 30938
rect 20720 30874 20772 30880
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20260 30320 20312 30326
rect 20260 30262 20312 30268
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18892 29646 18920 30194
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 20640 29238 20668 30602
rect 20732 30054 20760 30670
rect 20720 30048 20772 30054
rect 20720 29990 20772 29996
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 17868 28484 17920 28490
rect 17868 28426 17920 28432
rect 17880 28218 17908 28426
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17972 28150 18000 28494
rect 17960 28144 18012 28150
rect 17960 28086 18012 28092
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17972 27470 18000 28086
rect 18064 27878 18092 28494
rect 20088 28422 20116 29106
rect 20260 29028 20312 29034
rect 20260 28970 20312 28976
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17604 25294 17632 27338
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 17880 26450 17908 26862
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 16948 24880 17000 24886
rect 16948 24822 17000 24828
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17512 24274 17540 24686
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 16856 24132 16908 24138
rect 16856 24074 16908 24080
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16396 22500 16448 22506
rect 16396 22442 16448 22448
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 15476 21956 15528 21962
rect 15476 21898 15528 21904
rect 15488 21622 15516 21898
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15476 21616 15528 21622
rect 15476 21558 15528 21564
rect 15764 21554 15792 21830
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15292 21072 15344 21078
rect 15292 21014 15344 21020
rect 15200 20936 15252 20942
rect 15304 20924 15332 21014
rect 15396 20942 15424 21286
rect 15856 21146 15884 21490
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 15252 20896 15332 20924
rect 15200 20878 15252 20884
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 14752 19446 14780 19790
rect 15028 19718 15056 19790
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 15212 19310 15240 19722
rect 15304 19446 15332 20896
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15580 20466 15608 21082
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 17814 14412 18226
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14200 13938 14228 15642
rect 14278 15192 14334 15201
rect 14278 15127 14334 15136
rect 14292 14618 14320 15127
rect 14384 14958 14412 17070
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14476 14278 14504 19110
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 15028 18426 15056 18634
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14752 17678 14780 18158
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14660 16522 14688 16934
rect 14844 16794 14872 17818
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14844 16130 14872 16730
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14752 16102 14872 16130
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14476 14006 14504 14214
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14108 12374 14136 13738
rect 14292 13462 14320 13738
rect 14568 13734 14596 15302
rect 14660 14006 14688 16050
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14752 13870 14780 16102
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14844 15026 14872 15982
rect 15028 15978 15056 18362
rect 15304 18290 15332 19382
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14936 14618 14964 15846
rect 15028 15162 15056 15914
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14936 14414 14964 14554
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14556 13728 14608 13734
rect 14370 13696 14426 13705
rect 14556 13670 14608 13676
rect 14646 13696 14702 13705
rect 14370 13631 14426 13640
rect 14280 13456 14332 13462
rect 14200 13416 14280 13444
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14200 12306 14228 13416
rect 14280 13398 14332 13404
rect 14384 12646 14412 13631
rect 14568 13394 14596 13670
rect 14646 13631 14702 13640
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14372 12640 14424 12646
rect 14476 12617 14504 12718
rect 14568 12714 14596 13330
rect 14660 12850 14688 13631
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14372 12582 14424 12588
rect 14462 12608 14518 12617
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14200 11762 14228 12242
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14292 11506 14320 12582
rect 14660 12594 14688 12786
rect 14462 12543 14518 12552
rect 14568 12566 14688 12594
rect 14568 11898 14596 12566
rect 14936 12434 14964 14350
rect 15120 12986 15148 18226
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15212 17270 15240 17478
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15396 15706 15424 19450
rect 15488 19378 15516 19654
rect 15580 19446 15608 20402
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 19922 15792 20198
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15580 18834 15608 19382
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15488 17882 15516 18702
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18358 15608 18566
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15856 18290 15884 18838
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15488 17270 15516 17818
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15580 16794 15608 18158
rect 15672 17954 15700 18226
rect 15672 17926 15792 17954
rect 15764 17882 15792 17926
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15948 17678 15976 19450
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16040 17746 16068 18158
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15212 12434 15240 15302
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 12714 15332 13874
rect 15396 13394 15424 15030
rect 15488 14074 15516 15370
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15382 12880 15438 12889
rect 15488 12850 15516 13806
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15382 12815 15438 12824
rect 15476 12844 15528 12850
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15396 12646 15424 12815
rect 15476 12786 15528 12792
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 14752 12406 14964 12434
rect 15120 12406 15240 12434
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14200 11478 14320 11506
rect 14200 10674 14228 11478
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14108 10198 14136 10610
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14108 8634 14136 10134
rect 14292 10062 14320 11086
rect 14370 10704 14426 10713
rect 14370 10639 14372 10648
rect 14424 10639 14426 10648
rect 14372 10610 14424 10616
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14292 9518 14320 9998
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14016 8090 14044 8434
rect 14292 8430 14320 9454
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14292 7750 14320 8366
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7546 14320 7686
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6390 14136 6598
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14108 5710 14136 6326
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 14016 4457 14044 4490
rect 14002 4448 14058 4457
rect 14002 4383 14058 4392
rect 13910 3904 13966 3913
rect 13910 3839 13966 3848
rect 13726 3632 13782 3641
rect 14188 3596 14240 3602
rect 13726 3567 13782 3576
rect 13924 3556 14136 3584
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3126 13768 3334
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13818 2816 13874 2825
rect 13818 2751 13874 2760
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13740 1426 13768 2246
rect 13728 1420 13780 1426
rect 13728 1362 13780 1368
rect 13832 800 13860 2751
rect 13924 800 13952 3556
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 14016 2854 14044 3402
rect 14108 3194 14136 3556
rect 14188 3538 14240 3544
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14200 2854 14228 3538
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14108 800 14136 2450
rect 14292 1494 14320 6802
rect 14384 3618 14412 9046
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14476 8022 14504 8910
rect 14568 8242 14596 11698
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14660 8430 14688 8774
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14568 8214 14688 8242
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14476 6798 14504 7958
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14568 5778 14596 6258
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14660 5658 14688 8214
rect 14568 5630 14688 5658
rect 14568 3738 14596 5630
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14660 4826 14688 5034
rect 14752 5030 14780 12406
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14844 10470 14872 11018
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15028 9586 15056 9862
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14844 7546 14872 7754
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14844 7410 14872 7482
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14844 6934 14872 7346
rect 14832 6928 14884 6934
rect 14936 6905 14964 8570
rect 14832 6870 14884 6876
rect 14922 6896 14978 6905
rect 14922 6831 14978 6840
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14844 6458 14872 6734
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 15028 5370 15056 8774
rect 15120 6934 15148 12406
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15212 5914 15240 8978
rect 15304 7886 15332 9114
rect 15396 8838 15424 12582
rect 15488 12102 15516 12786
rect 15672 12442 15700 12854
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15764 11830 15792 17002
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 14890 16160 16050
rect 16224 15910 16252 21082
rect 16302 19952 16358 19961
rect 16302 19887 16358 19896
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 16316 14550 16344 19887
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 15856 14074 15884 14214
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15856 13977 15884 14010
rect 15842 13968 15898 13977
rect 15842 13903 15844 13912
rect 15896 13903 15898 13912
rect 15844 13874 15896 13880
rect 15856 13843 15884 13874
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15488 10062 15516 10542
rect 15672 10062 15700 11222
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10674 15976 10950
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15488 9042 15516 9998
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15856 8566 15884 8774
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14936 5250 14964 5306
rect 14936 5234 15056 5250
rect 14936 5228 15068 5234
rect 14936 5222 15016 5228
rect 15016 5170 15068 5176
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 4842 14780 4966
rect 14648 4820 14700 4826
rect 14752 4814 14964 4842
rect 14648 4762 14700 4768
rect 14936 4758 14964 4814
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15028 4622 15056 5170
rect 15212 5098 15240 5646
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5098 15332 5578
rect 15396 5302 15424 5646
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15304 4622 15332 5034
rect 15580 4622 15608 7210
rect 15016 4616 15068 4622
rect 14922 4584 14978 4593
rect 15016 4558 15068 4564
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 14922 4519 14978 4528
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14660 3738 14688 4082
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14384 3590 14504 3618
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14384 3233 14412 3470
rect 14370 3224 14426 3233
rect 14370 3159 14426 3168
rect 14280 1488 14332 1494
rect 14280 1430 14332 1436
rect 14188 1420 14240 1426
rect 14188 1362 14240 1368
rect 14200 800 14228 1362
rect 14384 800 14412 3159
rect 14476 2774 14504 3590
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14556 3392 14608 3398
rect 14648 3392 14700 3398
rect 14556 3334 14608 3340
rect 14646 3360 14648 3369
rect 14700 3360 14702 3369
rect 14568 3126 14596 3334
rect 14646 3295 14702 3304
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 14556 2984 14608 2990
rect 14554 2952 14556 2961
rect 14608 2952 14610 2961
rect 14554 2887 14610 2896
rect 14476 2746 14596 2774
rect 14464 2576 14516 2582
rect 14464 2518 14516 2524
rect 14476 800 14504 2518
rect 14568 2514 14596 2746
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14568 2106 14596 2314
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 14660 800 14688 1906
rect 14752 800 14780 3470
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14844 1426 14872 2858
rect 14936 2854 14964 4519
rect 15028 3942 15056 4558
rect 15106 4312 15162 4321
rect 15106 4247 15162 4256
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 15120 2774 15148 4247
rect 15304 4146 15332 4558
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15672 3602 15700 7686
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15764 3534 15792 4422
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15948 3126 15976 10610
rect 16040 8838 16068 12106
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16132 9382 16160 9930
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15120 2746 15332 2774
rect 15014 2680 15070 2689
rect 15014 2615 15016 2624
rect 15068 2615 15070 2624
rect 15016 2586 15068 2592
rect 15016 1488 15068 1494
rect 15016 1430 15068 1436
rect 14832 1420 14884 1426
rect 14832 1362 14884 1368
rect 15028 800 15056 1430
rect 15304 800 15332 2746
rect 15566 2272 15622 2281
rect 15566 2207 15622 2216
rect 15580 800 15608 2207
rect 15672 1222 15700 2858
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15660 1216 15712 1222
rect 15660 1158 15712 1164
rect 15856 800 15884 2790
rect 16040 2446 16068 6598
rect 16132 4146 16160 9318
rect 16316 8906 16344 14214
rect 16408 11354 16436 22442
rect 16580 21616 16632 21622
rect 16578 21584 16580 21593
rect 16632 21584 16634 21593
rect 16578 21519 16634 21528
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16592 14618 16620 21286
rect 16684 20942 16712 23258
rect 16776 23118 16804 23666
rect 16868 23322 16896 24074
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 17420 22642 17448 23666
rect 17512 23594 17540 24210
rect 17604 24206 17632 25230
rect 17880 24750 17908 26386
rect 17972 26382 18000 27406
rect 18064 26790 18092 27814
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 18156 27062 18184 27542
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18052 26784 18104 26790
rect 18052 26726 18104 26732
rect 18248 26382 18276 27270
rect 18524 26518 18552 27406
rect 18512 26512 18564 26518
rect 18512 26454 18564 26460
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 17972 24818 18000 26318
rect 18788 26240 18840 26246
rect 18788 26182 18840 26188
rect 18800 25430 18828 26182
rect 18604 25424 18656 25430
rect 18604 25366 18656 25372
rect 18788 25424 18840 25430
rect 18788 25366 18840 25372
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18156 24818 18184 25094
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17972 24206 18000 24754
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 18156 24070 18184 24618
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 17604 23730 17632 24006
rect 18248 23730 18276 24074
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17512 23186 17540 23530
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17604 22778 17632 23054
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17592 22772 17644 22778
rect 17592 22714 17644 22720
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17604 22234 17632 22714
rect 17696 22710 17724 22918
rect 17684 22704 17736 22710
rect 17684 22646 17736 22652
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16868 20602 16896 20810
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 17788 19990 17816 23258
rect 18248 23118 18276 23666
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 18328 23044 18380 23050
rect 18328 22986 18380 22992
rect 18340 22778 18368 22986
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17972 20466 18000 20810
rect 18064 20534 18092 21422
rect 18052 20528 18104 20534
rect 18052 20470 18104 20476
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16868 19310 16896 19722
rect 17328 19378 17356 19790
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16684 17814 16712 19110
rect 17328 18970 17356 19314
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17328 18290 17356 18906
rect 17420 18426 17448 19314
rect 18156 18630 18184 22714
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18524 21146 18552 21830
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18248 19553 18276 20878
rect 18512 20800 18564 20806
rect 18510 20768 18512 20777
rect 18564 20768 18566 20777
rect 18510 20703 18566 20712
rect 18234 19544 18290 19553
rect 18234 19479 18290 19488
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16868 17610 16896 18226
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16868 17270 16896 17546
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16684 15026 16712 16118
rect 16776 16046 16804 16594
rect 16868 16182 16896 17206
rect 16960 16590 16988 17614
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16856 16176 16908 16182
rect 16856 16118 16908 16124
rect 16960 16046 16988 16526
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16776 15502 16804 15846
rect 16960 15502 16988 15982
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 17052 15026 17080 15506
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16684 14414 16712 14758
rect 17144 14618 17172 18022
rect 17236 17678 17264 18022
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17328 17202 17356 18226
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17604 17678 17632 18022
rect 17696 17882 17724 18294
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16590 17540 16934
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17604 16436 17632 17614
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 17696 16590 17724 16662
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17788 16522 17816 17546
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18064 16794 18092 17138
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17512 16408 17632 16436
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17420 13530 17448 13942
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17130 13016 17186 13025
rect 17130 12951 17132 12960
rect 17184 12951 17186 12960
rect 17132 12922 17184 12928
rect 17512 12238 17540 16408
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15570 17632 15846
rect 17788 15638 17816 16458
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 13977 17632 14350
rect 17590 13968 17646 13977
rect 17590 13903 17646 13912
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17604 12986 17632 13194
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17696 12918 17724 15370
rect 17880 14890 17908 15438
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 15094 18000 15302
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 18156 14822 18184 16730
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17408 12232 17460 12238
rect 16578 12200 16634 12209
rect 17408 12174 17460 12180
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 16578 12135 16634 12144
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16486 11248 16542 11257
rect 16486 11183 16488 11192
rect 16540 11183 16542 11192
rect 16488 11154 16540 11160
rect 16592 11150 16620 12135
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 17314 10976 17370 10985
rect 17314 10911 17370 10920
rect 17222 10704 17278 10713
rect 17328 10674 17356 10911
rect 17222 10639 17278 10648
rect 17316 10668 17368 10674
rect 17236 10606 17264 10639
rect 17316 10610 17368 10616
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9042 16436 10066
rect 17052 10062 17080 10406
rect 17420 10130 17448 12174
rect 17512 11694 17540 12174
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17604 11150 17632 11766
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17512 9466 17540 9998
rect 17788 9674 17816 14214
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17866 13016 17922 13025
rect 17866 12951 17922 12960
rect 17880 12850 17908 12951
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17972 12434 18000 13738
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12850 18092 13126
rect 18432 12850 18460 13262
rect 18052 12844 18104 12850
rect 18236 12844 18288 12850
rect 18052 12786 18104 12792
rect 18156 12804 18236 12832
rect 18156 12434 18184 12804
rect 18236 12786 18288 12792
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 17880 12406 18000 12434
rect 18064 12406 18184 12434
rect 17880 12374 17908 12406
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 18064 12102 18092 12406
rect 18236 12300 18288 12306
rect 18340 12288 18368 12718
rect 18288 12260 18368 12288
rect 18236 12242 18288 12248
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17880 11762 17908 12038
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 18064 11150 18092 12038
rect 18156 11898 18184 12174
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18340 11558 18368 12260
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18340 11150 18368 11494
rect 18524 11150 18552 18702
rect 18616 14822 18644 25366
rect 18788 21956 18840 21962
rect 18788 21898 18840 21904
rect 18694 19000 18750 19009
rect 18694 18935 18696 18944
rect 18748 18935 18750 18944
rect 18696 18906 18748 18912
rect 18708 18766 18736 18906
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 16697 18736 18566
rect 18694 16688 18750 16697
rect 18694 16623 18750 16632
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14618 18644 14758
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18616 12918 18644 13806
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10810 18368 10950
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18524 10674 18552 11086
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18144 10464 18196 10470
rect 18064 10424 18144 10452
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17788 9646 17908 9674
rect 17236 9438 17540 9466
rect 17236 9382 17264 9438
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16408 8786 16436 8978
rect 16316 8758 16436 8786
rect 16316 8022 16344 8758
rect 16868 8362 16896 9318
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17328 8362 17356 8910
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16316 6662 16344 7958
rect 16776 7206 16804 8026
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16316 5370 16344 5578
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16118 3632 16174 3641
rect 16118 3567 16174 3576
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16132 800 16160 3567
rect 16408 800 16436 7142
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16500 2774 16528 6054
rect 16672 5568 16724 5574
rect 16592 5516 16672 5522
rect 16592 5510 16724 5516
rect 16592 5494 16712 5510
rect 16592 5234 16620 5494
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16592 4185 16620 5170
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 16684 3534 16712 4422
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16776 3058 16804 7142
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16868 5166 16896 5578
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16868 4282 16896 4558
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16500 2746 16712 2774
rect 16684 800 16712 2746
rect 16960 800 16988 8298
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 7206 17264 7686
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 6866 17264 7142
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5302 17172 5714
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17144 2650 17172 4558
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17236 800 17264 3334
rect 17328 3058 17356 8298
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 6798 17632 7822
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17788 6458 17816 7958
rect 17880 7750 17908 9646
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17592 6180 17644 6186
rect 17592 6122 17644 6128
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17512 4622 17540 6054
rect 17604 5817 17632 6122
rect 17590 5808 17646 5817
rect 17696 5778 17724 6190
rect 17788 6118 17816 6190
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17590 5743 17646 5752
rect 17684 5772 17736 5778
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 4146 17540 4422
rect 17500 4140 17552 4146
rect 17604 4128 17632 5743
rect 17684 5714 17736 5720
rect 17682 5264 17738 5273
rect 17682 5199 17738 5208
rect 17696 5030 17724 5199
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17696 4690 17724 4966
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17684 4140 17736 4146
rect 17604 4100 17684 4128
rect 17500 4082 17552 4088
rect 17684 4082 17736 4088
rect 17500 4004 17552 4010
rect 17500 3946 17552 3952
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17512 800 17540 3946
rect 17590 2544 17646 2553
rect 17590 2479 17646 2488
rect 17604 2310 17632 2479
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17604 2038 17632 2246
rect 17592 2032 17644 2038
rect 17592 1974 17644 1980
rect 17788 800 17816 5034
rect 17880 4486 17908 6258
rect 17972 5914 18000 9930
rect 18064 6798 18092 10424
rect 18144 10406 18196 10412
rect 18248 9194 18276 10610
rect 18800 10470 18828 21898
rect 18892 21672 18920 28018
rect 19984 27872 20036 27878
rect 19984 27814 20036 27820
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19248 26784 19300 26790
rect 19248 26726 19300 26732
rect 19260 25838 19288 26726
rect 19340 26308 19392 26314
rect 19340 26250 19392 26256
rect 19352 25906 19380 26250
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 19064 25424 19116 25430
rect 19064 25366 19116 25372
rect 18892 21644 19012 21672
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18892 20942 18920 21490
rect 18880 20936 18932 20942
rect 18878 20904 18880 20913
rect 18932 20904 18934 20913
rect 18878 20839 18934 20848
rect 18892 20813 18920 20839
rect 18984 17377 19012 21644
rect 18970 17368 19026 17377
rect 18970 17303 19026 17312
rect 18984 16454 19012 17303
rect 19076 16590 19104 25366
rect 19260 25294 19288 25774
rect 19444 25702 19472 27338
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19708 26376 19760 26382
rect 19706 26344 19708 26353
rect 19760 26344 19762 26353
rect 19706 26279 19762 26288
rect 19720 26246 19748 26279
rect 19708 26240 19760 26246
rect 19708 26182 19760 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19156 24132 19208 24138
rect 19156 24074 19208 24080
rect 19168 23322 19196 24074
rect 19260 23662 19288 25230
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19352 24750 19380 25162
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19996 24818 20024 27814
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19444 24290 19472 24754
rect 19524 24676 19576 24682
rect 19524 24618 19576 24624
rect 19352 24262 19472 24290
rect 19352 24070 19380 24262
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19340 24064 19392 24070
rect 19338 24032 19340 24041
rect 19392 24032 19394 24041
rect 19338 23967 19394 23976
rect 19444 23866 19472 24142
rect 19536 24052 19564 24618
rect 19516 24024 19564 24052
rect 19984 24064 20036 24070
rect 19432 23860 19484 23866
rect 19516 23848 19544 24024
rect 19984 24006 20036 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19516 23820 19564 23848
rect 19432 23802 19484 23808
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19156 23316 19208 23322
rect 19156 23258 19208 23264
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19352 23225 19380 23258
rect 19338 23216 19394 23225
rect 19338 23151 19394 23160
rect 19536 22964 19564 23820
rect 19996 23798 20024 24006
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19444 22936 19564 22964
rect 19444 22234 19472 22936
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19444 21554 19472 21898
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 20088 21554 20116 28358
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 19444 21146 19472 21490
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19338 20496 19394 20505
rect 19338 20431 19394 20440
rect 19246 17232 19302 17241
rect 19246 17167 19302 17176
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 15910 19012 16390
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18984 15314 19012 15846
rect 19076 15502 19104 16526
rect 19260 16250 19288 17167
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 18984 15286 19104 15314
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18878 13424 18934 13433
rect 18878 13359 18880 13368
rect 18932 13359 18934 13368
rect 18880 13330 18932 13336
rect 18984 12986 19012 15098
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18984 12850 19012 12922
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18984 11898 19012 12106
rect 19076 12102 19104 15286
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18984 11150 19012 11698
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 19168 10606 19196 15438
rect 19260 12374 19288 16186
rect 19352 15502 19380 20431
rect 19444 18068 19472 21082
rect 20180 20942 20208 26930
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 20810
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 18698 20024 20538
rect 20272 19802 20300 28970
rect 20628 28484 20680 28490
rect 20628 28426 20680 28432
rect 20640 28218 20668 28426
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20444 27668 20496 27674
rect 20444 27610 20496 27616
rect 20456 27130 20484 27610
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20364 24070 20392 24754
rect 20352 24064 20404 24070
rect 20350 24032 20352 24041
rect 20404 24032 20406 24041
rect 20350 23967 20406 23976
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20180 19774 20300 19802
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20088 18766 20116 19110
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19524 18080 19576 18086
rect 19444 18040 19524 18068
rect 19524 18022 19576 18028
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19444 16726 19472 17546
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20088 17270 20116 18702
rect 20180 17678 20208 19774
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20272 19378 20300 19654
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20076 17264 20128 17270
rect 19982 17232 20038 17241
rect 20076 17206 20128 17212
rect 19982 17167 19984 17176
rect 20036 17167 20038 17176
rect 19984 17138 20036 17144
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19444 16250 19472 16662
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19352 14346 19380 15302
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19444 14278 19472 16186
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19628 15570 19656 15914
rect 20272 15706 20300 19314
rect 20364 17678 20392 23734
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20456 20602 20484 22578
rect 20548 22166 20576 25162
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20640 22438 20668 23054
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20640 22234 20668 22374
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 20732 22098 20760 29990
rect 20916 29646 20944 31282
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 21824 30184 21876 30190
rect 21824 30126 21876 30132
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21560 29646 21588 29786
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 21548 29640 21600 29646
rect 21548 29582 21600 29588
rect 20916 29306 20944 29582
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 21272 29300 21324 29306
rect 21272 29242 21324 29248
rect 21088 29232 21140 29238
rect 21088 29174 21140 29180
rect 20996 28960 21048 28966
rect 20996 28902 21048 28908
rect 20904 28076 20956 28082
rect 21008 28064 21036 28902
rect 21100 28626 21128 29174
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 21284 28082 21312 29242
rect 21560 28966 21588 29582
rect 21836 29238 21864 30126
rect 21928 29850 21956 30194
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 22112 29578 22140 31214
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22480 29646 22508 29990
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 21824 29232 21876 29238
rect 21824 29174 21876 29180
rect 21548 28960 21600 28966
rect 21548 28902 21600 28908
rect 21088 28076 21140 28082
rect 21008 28036 21088 28064
rect 20904 28018 20956 28024
rect 21088 28018 21140 28024
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 20916 27674 20944 28018
rect 21560 28014 21588 28902
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21548 28008 21600 28014
rect 21548 27950 21600 27956
rect 20904 27668 20956 27674
rect 20904 27610 20956 27616
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 21008 26518 21036 26998
rect 21836 26994 21864 28494
rect 22112 28218 22140 29514
rect 22664 29170 22692 29582
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22112 27538 22140 28154
rect 22204 28150 22232 28970
rect 22664 28762 22692 29106
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 22756 28626 22784 31350
rect 23032 30122 23060 31350
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 23308 30326 23336 31282
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23296 30320 23348 30326
rect 23296 30262 23348 30268
rect 23020 30116 23072 30122
rect 23020 30058 23072 30064
rect 22376 28620 22428 28626
rect 22376 28562 22428 28568
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 22388 28150 22416 28562
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 22836 28008 22888 28014
rect 22836 27950 22888 27956
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22008 27464 22060 27470
rect 22008 27406 22060 27412
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 20996 26512 21048 26518
rect 20996 26454 21048 26460
rect 20904 25424 20956 25430
rect 20904 25366 20956 25372
rect 20916 24682 20944 25366
rect 20904 24676 20956 24682
rect 20904 24618 20956 24624
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20916 23118 20944 24142
rect 21008 23798 21036 26454
rect 21088 24812 21140 24818
rect 21192 24800 21220 26930
rect 22020 25838 22048 27406
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22100 26308 22152 26314
rect 22100 26250 22152 26256
rect 22112 26042 22140 26250
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22664 25906 22692 26726
rect 22848 26489 22876 27950
rect 22834 26480 22890 26489
rect 22834 26415 22836 26424
rect 22888 26415 22890 26424
rect 22836 26386 22888 26392
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 22020 25378 22048 25774
rect 21140 24772 21220 24800
rect 21836 25350 22048 25378
rect 21088 24754 21140 24760
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 21100 23322 21128 24754
rect 21836 24274 21864 25350
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 21824 24268 21876 24274
rect 21824 24210 21876 24216
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21192 23526 21220 23666
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 21192 23254 21220 23462
rect 21180 23248 21232 23254
rect 21180 23190 21232 23196
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20534 21992 20590 22001
rect 20534 21927 20536 21936
rect 20588 21927 20590 21936
rect 20536 21898 20588 21904
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20548 21434 20576 21490
rect 20732 21434 20760 21830
rect 20548 21406 20760 21434
rect 20732 21162 20760 21406
rect 20824 21350 20852 22578
rect 20916 22030 20944 23054
rect 21192 23050 21220 23190
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21284 22778 21312 23054
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 20996 22160 21048 22166
rect 20996 22102 21048 22108
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20732 21134 20852 21162
rect 20916 21146 20944 21490
rect 20536 21072 20588 21078
rect 20536 21014 20588 21020
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20442 19544 20498 19553
rect 20442 19479 20498 19488
rect 20456 18306 20484 19479
rect 20548 18970 20576 21014
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20534 20760 20742
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20732 19922 20760 20470
rect 20824 20466 20852 21134
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 21008 20380 21036 22102
rect 21284 21894 21312 22714
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21284 20777 21312 21830
rect 21270 20768 21326 20777
rect 21270 20703 21326 20712
rect 20916 20352 21036 20380
rect 21088 20392 21140 20398
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20628 19780 20680 19786
rect 20628 19722 20680 19728
rect 20640 19242 20668 19722
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20732 18834 20760 19858
rect 20916 19378 20944 20352
rect 21088 20334 21140 20340
rect 21100 20058 21128 20334
rect 21376 20058 21404 22986
rect 21744 21978 21772 23598
rect 21928 23322 21956 25230
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22020 24614 22048 24754
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 22020 23168 22048 24550
rect 22284 24336 22336 24342
rect 22284 24278 22336 24284
rect 22296 23866 22324 24278
rect 22480 23905 22508 25842
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22572 24954 22600 25230
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22664 24206 22692 25230
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22466 23896 22522 23905
rect 22284 23860 22336 23866
rect 22466 23831 22522 23840
rect 22284 23802 22336 23808
rect 21928 23140 22048 23168
rect 21560 21950 21772 21978
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21560 21729 21588 21950
rect 21546 21720 21602 21729
rect 21546 21655 21602 21664
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20904 19372 20956 19378
rect 21008 19352 21036 19654
rect 20904 19314 20956 19320
rect 20996 19346 21048 19352
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20720 18352 20772 18358
rect 20456 18278 20576 18306
rect 20720 18294 20772 18300
rect 20548 17785 20576 18278
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20534 17776 20590 17785
rect 20534 17711 20590 17720
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20364 16153 20392 17206
rect 20548 16658 20576 17546
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20534 16552 20590 16561
rect 20534 16487 20590 16496
rect 20350 16144 20406 16153
rect 20350 16079 20406 16088
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 19708 15700 19760 15706
rect 19708 15642 19760 15648
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19720 15502 19748 15642
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 20074 15600 20130 15609
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19996 15337 20024 15574
rect 20180 15586 20208 15642
rect 20180 15558 20300 15586
rect 20074 15535 20130 15544
rect 19982 15328 20038 15337
rect 19574 15260 19882 15269
rect 19982 15263 20038 15272
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15201 20116 15535
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20074 15192 20130 15201
rect 20074 15127 20130 15136
rect 20180 14929 20208 15438
rect 20272 15366 20300 15558
rect 20364 15502 20392 15846
rect 20456 15570 20484 15982
rect 20548 15910 20576 16487
rect 20536 15904 20588 15910
rect 20534 15872 20536 15881
rect 20588 15872 20590 15881
rect 20534 15807 20590 15816
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20166 14920 20222 14929
rect 20166 14855 20222 14864
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19904 13954 19932 14010
rect 19996 13954 20024 14418
rect 20076 14272 20128 14278
rect 20074 14240 20076 14249
rect 20272 14260 20300 15302
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20128 14240 20300 14260
rect 20130 14232 20300 14240
rect 20074 14175 20130 14184
rect 20166 14104 20222 14113
rect 20166 14039 20222 14048
rect 19904 13926 20024 13954
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 11762 19288 12174
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19352 11218 19380 13262
rect 19628 13172 19656 13806
rect 19516 13144 19656 13172
rect 19516 12968 19544 13144
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19516 12940 19564 12968
rect 19432 12096 19484 12102
rect 19430 12064 19432 12073
rect 19536 12084 19564 12940
rect 20079 12232 20131 12238
rect 20079 12174 20131 12180
rect 19484 12064 19486 12073
rect 19430 11999 19486 12008
rect 19516 12056 19564 12084
rect 19516 11880 19544 12056
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19516 11852 19564 11880
rect 19536 11694 19564 11852
rect 19708 11824 19760 11830
rect 19706 11792 19708 11801
rect 19760 11792 19762 11801
rect 20088 11762 20116 12174
rect 19706 11727 19762 11736
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19812 11393 19840 11562
rect 19798 11384 19854 11393
rect 19996 11354 20024 11698
rect 20088 11558 20116 11698
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19798 11319 19854 11328
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 19352 10062 19380 11018
rect 19444 10266 19472 11222
rect 19982 11112 20038 11121
rect 19982 11047 20038 11056
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19536 10674 19564 10746
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 18328 9920 18380 9926
rect 19536 9908 19564 10474
rect 18328 9862 18380 9868
rect 19444 9880 19564 9908
rect 18340 9586 18368 9862
rect 19444 9722 19472 9880
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18156 9166 18276 9194
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 3738 17908 4422
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17972 3398 18000 4218
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17866 2816 17922 2825
rect 17866 2751 17922 2760
rect 17880 2514 17908 2751
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 18064 800 18092 5646
rect 18156 2774 18184 9166
rect 18616 8276 18644 9454
rect 19892 9376 19944 9382
rect 19890 9344 19892 9353
rect 19944 9344 19946 9353
rect 19890 9279 19946 9288
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18696 8288 18748 8294
rect 18616 8248 18696 8276
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7410 18276 7686
rect 18432 7546 18460 7754
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18616 7342 18644 8248
rect 18696 8230 18748 8236
rect 18984 7342 19012 8842
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 18616 6866 18644 7278
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18512 6792 18564 6798
rect 18236 6770 18288 6776
rect 18512 6734 18564 6740
rect 18236 6712 18288 6718
rect 18248 5914 18276 6712
rect 18524 6662 18552 6734
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18234 4448 18290 4457
rect 18234 4383 18290 4392
rect 18248 4214 18276 4383
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18156 2746 18276 2774
rect 18248 2582 18276 2746
rect 18236 2576 18288 2582
rect 18236 2518 18288 2524
rect 18248 2417 18276 2518
rect 18234 2408 18290 2417
rect 18234 2343 18290 2352
rect 18340 800 18368 5782
rect 18524 3670 18552 6598
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18512 3664 18564 3670
rect 18512 3606 18564 3612
rect 18616 800 18644 6054
rect 18708 5642 18736 6326
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18800 4264 18828 7142
rect 18984 4554 19012 7278
rect 19168 5846 19196 8434
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5370 19380 5646
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 18972 4548 19024 4554
rect 18972 4490 19024 4496
rect 18708 4236 18828 4264
rect 18708 2854 18736 4236
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18800 2106 18828 4082
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18892 800 18920 3878
rect 19168 800 19196 5102
rect 19260 4554 19288 5170
rect 19444 5114 19472 6054
rect 19996 5574 20024 11047
rect 20088 10674 20116 11494
rect 20180 10810 20208 14039
rect 20364 12424 20392 15098
rect 20548 14618 20576 15370
rect 20640 15026 20668 18226
rect 20732 17660 20760 18294
rect 20916 17882 20944 19314
rect 20996 19288 21048 19294
rect 21100 19156 21128 19994
rect 21008 19128 21128 19156
rect 21456 19168 21508 19174
rect 21008 18086 21036 19128
rect 21456 19110 21508 19116
rect 21468 18766 21496 19110
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20812 17808 20864 17814
rect 21008 17762 21036 18022
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 20864 17756 21036 17762
rect 20812 17750 21036 17756
rect 20824 17734 21036 17750
rect 20812 17672 20864 17678
rect 20732 17632 20812 17660
rect 20812 17614 20864 17620
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20732 16454 20760 16526
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20718 15736 20774 15745
rect 20718 15671 20774 15680
rect 20732 15162 20760 15671
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20824 15094 20852 17206
rect 20916 17202 20944 17734
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20916 16250 20944 17138
rect 21192 16998 21220 17206
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 20996 16448 21048 16454
rect 20994 16416 20996 16425
rect 21048 16416 21050 16425
rect 20994 16351 21050 16360
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20916 14482 20944 16050
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21362 16008 21418 16017
rect 21100 15366 21128 15982
rect 21362 15943 21418 15952
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21376 15094 21404 15943
rect 21468 15706 21496 17818
rect 21560 17134 21588 21655
rect 21836 20806 21864 21966
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21836 20466 21864 20742
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21928 18766 21956 23140
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22020 22710 22048 22986
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22020 22098 22048 22510
rect 22112 22506 22140 23054
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22020 19378 22048 20538
rect 22112 19854 22140 21966
rect 22204 21962 22232 22034
rect 22480 22030 22508 23831
rect 22756 22982 22784 26318
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22836 22094 22888 22098
rect 22572 22092 22888 22094
rect 22572 22066 22836 22092
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22296 21622 22324 21966
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22480 21418 22508 21966
rect 22572 21962 22600 22066
rect 22836 22034 22888 22040
rect 22652 22024 22704 22030
rect 22704 21984 22784 22012
rect 22652 21966 22704 21972
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22480 21146 22508 21354
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22100 19848 22152 19854
rect 22098 19816 22100 19825
rect 22152 19816 22154 19825
rect 22098 19751 22154 19760
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21652 17066 21680 17818
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21560 15881 21588 16594
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21546 15872 21602 15881
rect 21546 15807 21602 15816
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21364 15088 21416 15094
rect 21364 15030 21416 15036
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 20534 14240 20590 14249
rect 20534 14175 20590 14184
rect 20548 13938 20576 14175
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20548 12850 20576 13330
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20364 12396 20484 12424
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20272 11762 20300 12310
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20456 11642 20484 12396
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20272 11614 20484 11642
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20180 8514 20208 8910
rect 20272 8634 20300 11614
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20364 9466 20392 11290
rect 20456 11082 20484 11494
rect 20548 11150 20576 11494
rect 20640 11150 20668 11698
rect 20732 11354 20760 14282
rect 21008 14074 21036 14282
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21008 13938 21036 14010
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20916 13274 20944 13874
rect 21192 13530 21220 14758
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21100 13433 21128 13466
rect 21086 13424 21142 13433
rect 21284 13394 21312 13874
rect 21468 13462 21496 15506
rect 21560 13938 21588 15807
rect 21652 14482 21680 16458
rect 21744 16182 21772 18702
rect 22020 17954 22048 19314
rect 22112 19174 22140 19751
rect 22204 19718 22232 20810
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22204 19378 22232 19654
rect 22189 19372 22241 19378
rect 22189 19314 22241 19320
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21836 17926 22048 17954
rect 21836 16250 21864 17926
rect 22008 17672 22060 17678
rect 21914 17640 21970 17649
rect 22008 17614 22060 17620
rect 21914 17575 21970 17584
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 21732 15496 21784 15502
rect 21928 15450 21956 17575
rect 22020 17202 22048 17614
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 22020 15570 22048 17138
rect 22112 16096 22140 18158
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22204 16561 22232 17138
rect 22296 16590 22324 18566
rect 22388 17898 22416 20742
rect 22664 20505 22692 21422
rect 22756 20534 22784 21984
rect 22940 21554 22968 23258
rect 23032 23118 23060 30058
rect 23112 30048 23164 30054
rect 23112 29990 23164 29996
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 23018 22264 23074 22273
rect 23018 22199 23074 22208
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 22744 20528 22796 20534
rect 22650 20496 22706 20505
rect 22744 20470 22796 20476
rect 22650 20431 22706 20440
rect 22468 20324 22520 20330
rect 22468 20266 22520 20272
rect 22480 19990 22508 20266
rect 22468 19984 22520 19990
rect 22468 19926 22520 19932
rect 22560 19346 22612 19352
rect 22560 19288 22612 19294
rect 22572 19174 22600 19288
rect 22664 19242 22692 20431
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22468 18216 22520 18222
rect 22466 18184 22468 18193
rect 22520 18184 22522 18193
rect 22466 18119 22522 18128
rect 22572 18086 22600 18702
rect 22940 18630 22968 19246
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 23032 18290 23060 22199
rect 23124 21418 23152 29990
rect 23308 29646 23336 30262
rect 23768 29782 23796 31214
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 23756 29776 23808 29782
rect 23756 29718 23808 29724
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23952 29578 23980 29990
rect 24044 29646 24072 31282
rect 24504 30682 24532 31282
rect 26148 31136 26200 31142
rect 26148 31078 26200 31084
rect 24412 30654 24532 30682
rect 24412 30598 24440 30654
rect 24400 30592 24452 30598
rect 24400 30534 24452 30540
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 23940 29572 23992 29578
rect 23940 29514 23992 29520
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23308 29170 23336 29446
rect 24044 29306 24072 29582
rect 24032 29300 24084 29306
rect 24032 29242 24084 29248
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23216 28150 23244 28358
rect 23768 28150 23796 28358
rect 23204 28144 23256 28150
rect 23204 28086 23256 28092
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23216 25498 23244 26930
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23400 26518 23428 26726
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23584 26382 23612 27066
rect 23768 26450 23796 28086
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23768 25906 23796 26386
rect 23756 25900 23808 25906
rect 23756 25842 23808 25848
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 23204 25492 23256 25498
rect 23204 25434 23256 25440
rect 23308 24410 23336 25774
rect 23664 25356 23716 25362
rect 23664 25298 23716 25304
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23492 24818 23520 25162
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23584 24818 23612 25094
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23216 23254 23244 24142
rect 23308 23508 23336 24346
rect 23492 23866 23520 24754
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23308 23480 23428 23508
rect 23204 23248 23256 23254
rect 23204 23190 23256 23196
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23204 22568 23256 22574
rect 23204 22510 23256 22516
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23110 20904 23166 20913
rect 23110 20839 23166 20848
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22756 18086 22784 18158
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22388 17870 22600 17898
rect 22468 17808 22520 17814
rect 22468 17750 22520 17756
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16590 22416 16934
rect 22284 16584 22336 16590
rect 22190 16552 22246 16561
rect 22284 16526 22336 16532
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22190 16487 22246 16496
rect 22480 16114 22508 17750
rect 22192 16108 22244 16114
rect 22112 16068 22192 16096
rect 22468 16108 22520 16114
rect 22244 16068 22324 16096
rect 22192 16050 22244 16056
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 21732 15438 21784 15444
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 21744 13954 21772 15438
rect 21836 15422 21956 15450
rect 22100 15428 22152 15434
rect 21836 14822 21864 15422
rect 22100 15370 22152 15376
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21928 14074 21956 14894
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21548 13932 21600 13938
rect 21744 13926 21864 13954
rect 21548 13874 21600 13880
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21652 13530 21680 13670
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21086 13359 21142 13368
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 20916 13258 21036 13274
rect 20916 13252 21048 13258
rect 20916 13246 20996 13252
rect 20996 13194 21048 13200
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20916 12306 20944 12854
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20640 10962 20668 11086
rect 20548 10934 20668 10962
rect 20548 9466 20576 10934
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20640 10266 20668 10746
rect 21008 10674 21036 13194
rect 21652 12986 21680 13466
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 20996 10668 21048 10674
rect 20824 10628 20996 10656
rect 20824 10538 20852 10628
rect 20996 10610 21048 10616
rect 20812 10532 20864 10538
rect 20732 10492 20812 10520
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20364 9438 20484 9466
rect 20548 9438 20668 9466
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 8974 20392 9318
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20180 8486 20300 8514
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20180 7886 20208 8366
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20076 6248 20128 6254
rect 20074 6216 20076 6225
rect 20128 6216 20130 6225
rect 20074 6151 20130 6160
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 20088 5574 20116 5714
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 19352 5086 19472 5114
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19260 800 19288 4490
rect 19352 4078 19380 5086
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19352 3466 19380 3878
rect 19444 3602 19472 4966
rect 19628 4486 19656 5170
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19524 4004 19576 4010
rect 19524 3946 19576 3952
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19432 3392 19484 3398
rect 19536 3380 19564 3946
rect 19628 3738 19656 4082
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19812 3482 19840 4014
rect 19890 3768 19946 3777
rect 19890 3703 19892 3712
rect 19944 3703 19946 3712
rect 19892 3674 19944 3680
rect 19996 3602 20024 4966
rect 20088 4758 20116 5170
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19812 3454 20024 3482
rect 19432 3334 19484 3340
rect 19516 3352 19564 3380
rect 19444 2428 19472 3334
rect 19516 3176 19544 3352
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19516 3148 19564 3176
rect 19352 2400 19472 2428
rect 19352 1154 19380 2400
rect 19536 2360 19564 3148
rect 19996 2650 20024 3454
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19444 2332 19564 2360
rect 19340 1148 19392 1154
rect 19340 1090 19392 1096
rect 19444 800 19472 2332
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 19536 800 19564 1294
rect 19708 1148 19760 1154
rect 19708 1090 19760 1096
rect 19720 800 19748 1090
rect 19812 800 19840 2042
rect 20088 1578 20116 4558
rect 20180 4010 20208 7822
rect 20272 7002 20300 8486
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20272 6322 20300 6938
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20272 5642 20300 6122
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20272 4690 20300 5578
rect 20364 5114 20392 8774
rect 20456 5302 20484 9438
rect 20534 9344 20590 9353
rect 20534 9279 20590 9288
rect 20548 8974 20576 9279
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20548 6390 20576 7142
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20536 5160 20588 5166
rect 20364 5086 20484 5114
rect 20536 5102 20588 5108
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20272 3602 20300 4626
rect 20364 4622 20392 4966
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20180 3058 20208 3470
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19996 1550 20116 1578
rect 19996 800 20024 1550
rect 20180 1442 20208 2994
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20088 1414 20208 1442
rect 20088 800 20116 1414
rect 20272 800 20300 2926
rect 20364 1358 20392 4422
rect 20456 4078 20484 5086
rect 20548 4078 20576 5102
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20352 1352 20404 1358
rect 20352 1294 20404 1300
rect 20456 800 20484 2858
rect 20536 2576 20588 2582
rect 20640 2564 20668 9438
rect 20732 7954 20760 10492
rect 20812 10474 20864 10480
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20916 9042 20944 10474
rect 21100 10470 21128 11698
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21100 9586 21128 10406
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20824 8566 20852 8774
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20732 7342 20760 7890
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6322 20852 6598
rect 20916 6458 20944 8978
rect 21192 7546 21220 12922
rect 21744 12889 21772 13262
rect 21730 12880 21786 12889
rect 21730 12815 21786 12824
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21364 9988 21416 9994
rect 21364 9930 21416 9936
rect 21376 9110 21404 9930
rect 21468 9654 21496 9998
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 21364 9104 21416 9110
rect 21364 9046 21416 9052
rect 21376 8498 21404 9046
rect 21468 8634 21496 9590
rect 21744 9586 21772 12815
rect 21836 10266 21864 13926
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12458 21956 13330
rect 22020 12918 22048 14894
rect 22112 13841 22140 15370
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22204 14278 22232 15302
rect 22296 14906 22324 16068
rect 22468 16050 22520 16056
rect 22468 15972 22520 15978
rect 22468 15914 22520 15920
rect 22374 15736 22430 15745
rect 22374 15671 22376 15680
rect 22428 15671 22430 15680
rect 22376 15642 22428 15648
rect 22376 15360 22428 15366
rect 22374 15328 22376 15337
rect 22428 15328 22430 15337
rect 22374 15263 22430 15272
rect 22296 14878 22416 14906
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22098 13832 22154 13841
rect 22098 13767 22154 13776
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 22204 12782 22232 14214
rect 22296 12850 22324 14758
rect 22388 14618 22416 14878
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 21928 12434 22140 12458
rect 22480 12434 22508 15914
rect 22572 13530 22600 17870
rect 22756 16522 22784 18022
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 23032 16726 23060 17546
rect 23020 16720 23072 16726
rect 23020 16662 23072 16668
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22848 16250 22876 16526
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22848 15706 22876 16186
rect 23020 16108 23072 16114
rect 23020 16050 23072 16056
rect 23032 15978 23060 16050
rect 23020 15972 23072 15978
rect 23020 15914 23072 15920
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 23124 15502 23152 20839
rect 23216 18193 23244 22510
rect 23308 19854 23336 23054
rect 23400 22166 23428 23480
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23492 22438 23520 22986
rect 23584 22506 23612 24142
rect 23676 23730 23704 25298
rect 23860 24342 23888 28494
rect 24044 26994 24072 29242
rect 24308 28484 24360 28490
rect 24308 28426 24360 28432
rect 24320 27674 24348 28426
rect 24412 27946 24440 30534
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 24504 29034 24532 30194
rect 24964 29646 24992 30262
rect 26160 30258 26188 31078
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 68100 30728 68152 30734
rect 68098 30696 68100 30705
rect 68152 30696 68154 30705
rect 68098 30631 68154 30640
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 26148 30252 26200 30258
rect 26148 30194 26200 30200
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 28264 30252 28316 30258
rect 28264 30194 28316 30200
rect 27632 29646 27660 30194
rect 24952 29640 25004 29646
rect 24952 29582 25004 29588
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 24964 29238 24992 29582
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25596 29572 25648 29578
rect 25596 29514 25648 29520
rect 25136 29504 25188 29510
rect 25136 29446 25188 29452
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 24492 29028 24544 29034
rect 24492 28970 24544 28976
rect 24400 27940 24452 27946
rect 24400 27882 24452 27888
rect 24308 27668 24360 27674
rect 24308 27610 24360 27616
rect 24400 27056 24452 27062
rect 24400 26998 24452 27004
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 24412 26518 24440 26998
rect 24400 26512 24452 26518
rect 24214 26480 24270 26489
rect 24400 26454 24452 26460
rect 24214 26415 24270 26424
rect 24032 25220 24084 25226
rect 24032 25162 24084 25168
rect 23848 24336 23900 24342
rect 23848 24278 23900 24284
rect 23756 24132 23808 24138
rect 23756 24074 23808 24080
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 23400 22030 23428 22102
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23400 20874 23428 21830
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23400 18873 23428 20198
rect 23386 18864 23442 18873
rect 23386 18799 23442 18808
rect 23202 18184 23258 18193
rect 23202 18119 23258 18128
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 16794 23428 16934
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 23112 15496 23164 15502
rect 23400 15473 23428 16730
rect 23492 16114 23520 22374
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 23584 17882 23612 22170
rect 23676 20942 23704 22918
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23768 18290 23796 24074
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 20262 23888 21490
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23860 16046 23888 20198
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23952 19446 23980 19722
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23952 18766 23980 19382
rect 24044 19378 24072 25162
rect 24228 24818 24256 26415
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 24228 24274 24256 24618
rect 24216 24268 24268 24274
rect 24216 24210 24268 24216
rect 24228 23662 24256 24210
rect 24308 24064 24360 24070
rect 24308 24006 24360 24012
rect 24320 23730 24348 24006
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24216 23656 24268 23662
rect 24216 23598 24268 23604
rect 24320 20602 24348 23666
rect 24412 22642 24440 26454
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24504 22094 24532 28970
rect 24860 28484 24912 28490
rect 24860 28426 24912 28432
rect 24584 27872 24636 27878
rect 24584 27814 24636 27820
rect 24596 27402 24624 27814
rect 24872 27402 24900 28426
rect 25148 27606 25176 29446
rect 25240 28218 25268 29514
rect 25228 28212 25280 28218
rect 25228 28154 25280 28160
rect 25136 27600 25188 27606
rect 25136 27542 25188 27548
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 24412 22066 24532 22094
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24136 19854 24164 19994
rect 24412 19854 24440 22066
rect 24596 22030 24624 27338
rect 24872 26926 24900 27338
rect 25148 27062 25176 27542
rect 25608 27470 25636 29514
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25780 28960 25832 28966
rect 25780 28902 25832 28908
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25700 28082 25728 28358
rect 25792 28218 25820 28902
rect 25884 28490 25912 29446
rect 26240 29028 26292 29034
rect 26240 28970 26292 28976
rect 26252 28490 26280 28970
rect 27632 28762 27660 29582
rect 27804 29572 27856 29578
rect 27804 29514 27856 29520
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 25872 28484 25924 28490
rect 25872 28426 25924 28432
rect 26240 28484 26292 28490
rect 26240 28426 26292 28432
rect 25780 28212 25832 28218
rect 25780 28154 25832 28160
rect 25688 28076 25740 28082
rect 25688 28018 25740 28024
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25596 27464 25648 27470
rect 25596 27406 25648 27412
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25136 27056 25188 27062
rect 25136 26998 25188 27004
rect 25240 26994 25268 27270
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24768 26240 24820 26246
rect 24768 26182 24820 26188
rect 24780 24954 24808 26182
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24872 23866 24900 24142
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24872 23118 24900 23802
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 25056 23322 25084 23598
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24768 22976 24820 22982
rect 24768 22918 24820 22924
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24688 21962 24716 22442
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24688 21622 24716 21898
rect 24676 21616 24728 21622
rect 24676 21558 24728 21564
rect 24124 19848 24176 19854
rect 24124 19790 24176 19796
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24136 19378 24164 19790
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23952 18290 23980 18702
rect 24136 18290 24164 19314
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 24136 18154 24164 18226
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 24136 17746 24164 18090
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23112 15438 23164 15444
rect 23386 15464 23442 15473
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22664 14890 22692 15098
rect 22652 14884 22704 14890
rect 22652 14826 22704 14832
rect 22756 14498 22784 15370
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22664 14470 22784 14498
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22664 13308 22692 14470
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22756 13462 22784 14350
rect 22848 14074 22876 14962
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22664 13280 22876 13308
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 21928 12430 22232 12434
rect 22112 12406 22232 12430
rect 22204 12238 22232 12406
rect 22388 12406 22508 12434
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22296 11801 22324 12038
rect 22282 11792 22338 11801
rect 22282 11727 22338 11736
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21928 10062 21956 11630
rect 22388 11014 22416 12406
rect 22664 12306 22692 12582
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22388 10674 22416 10950
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21928 9722 21956 9998
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21456 7880 21508 7886
rect 21454 7848 21456 7857
rect 21508 7848 21510 7857
rect 21454 7783 21510 7792
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21284 6798 21312 7346
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 20904 6452 20956 6458
rect 21284 6440 21312 6734
rect 21652 6730 21680 9522
rect 21928 8974 21956 9658
rect 22572 9654 22600 9862
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 22020 7886 22048 9522
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22204 7410 22232 7822
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22756 7206 22784 12718
rect 22848 9042 22876 13280
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22940 8945 22968 15438
rect 23386 15399 23442 15408
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23492 15337 23520 15370
rect 23478 15328 23534 15337
rect 23478 15263 23534 15272
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23032 13530 23060 14962
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 13938 23428 14214
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 23400 13394 23428 13738
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23032 11694 23060 12174
rect 23124 12102 23152 12582
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23400 11898 23428 13330
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23020 11688 23072 11694
rect 23020 11630 23072 11636
rect 23492 11286 23520 15263
rect 23584 11830 23612 15846
rect 24136 15450 24164 17478
rect 24228 17338 24256 18294
rect 24780 18290 24808 22918
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24872 22273 24900 22374
rect 24858 22264 24914 22273
rect 24858 22199 24914 22208
rect 24964 22030 24992 22578
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24964 21554 24992 21966
rect 24952 21548 25004 21554
rect 24952 21490 25004 21496
rect 24964 20466 24992 21490
rect 25044 21344 25096 21350
rect 25044 21286 25096 21292
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24872 18970 24900 19110
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24596 16658 24624 17546
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24228 15570 24256 16390
rect 24412 16182 24440 16390
rect 24400 16176 24452 16182
rect 24400 16118 24452 16124
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24136 15422 24256 15450
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23952 14006 23980 14758
rect 24124 14340 24176 14346
rect 24124 14282 24176 14288
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13326 23704 13670
rect 23860 13326 23888 13874
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23952 13258 23980 13942
rect 24136 13938 24164 14282
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24136 13258 24164 13874
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 24124 13252 24176 13258
rect 24124 13194 24176 13200
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12918 24072 13126
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23492 10810 23520 11222
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 23124 9926 23152 10678
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23676 9654 23704 11086
rect 23768 10674 23796 12038
rect 23952 11762 23980 12650
rect 24044 12374 24072 12718
rect 24032 12368 24084 12374
rect 24032 12310 24084 12316
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23860 11286 23888 11494
rect 24044 11354 24072 12106
rect 24122 11384 24178 11393
rect 24032 11348 24084 11354
rect 24228 11354 24256 15422
rect 24398 15192 24454 15201
rect 24398 15127 24454 15136
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24320 13802 24348 15030
rect 24412 14414 24440 15127
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24504 12986 24532 14418
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24596 12238 24624 16594
rect 24688 14618 24716 17206
rect 24964 17134 24992 20402
rect 25056 19961 25084 21286
rect 25148 21078 25176 24890
rect 25240 24818 25268 25230
rect 25504 25152 25556 25158
rect 25504 25094 25556 25100
rect 25516 24818 25544 25094
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25240 23730 25268 24754
rect 25504 24676 25556 24682
rect 25504 24618 25556 24624
rect 25516 23730 25544 24618
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25503 23724 25555 23730
rect 25503 23666 25555 23672
rect 25502 23216 25558 23225
rect 25502 23151 25504 23160
rect 25556 23151 25558 23160
rect 25504 23122 25556 23128
rect 25228 21888 25280 21894
rect 25228 21830 25280 21836
rect 25136 21072 25188 21078
rect 25136 21014 25188 21020
rect 25042 19952 25098 19961
rect 25042 19887 25098 19896
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25148 18086 25176 18634
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25148 17746 25176 18022
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25148 17134 25176 17478
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 24964 16590 24992 17070
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 25148 16250 25176 17070
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 24766 14920 24822 14929
rect 24766 14855 24768 14864
rect 24820 14855 24822 14864
rect 24768 14826 24820 14832
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24780 14278 24808 14826
rect 25240 14385 25268 21830
rect 25608 21554 25636 27406
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25700 25294 25728 27270
rect 25792 26994 25820 27950
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25792 26586 25820 26930
rect 25780 26580 25832 26586
rect 25780 26522 25832 26528
rect 25778 26480 25834 26489
rect 25778 26415 25780 26424
rect 25832 26415 25834 26424
rect 25780 26386 25832 26392
rect 25792 26042 25820 26386
rect 25780 26036 25832 26042
rect 25780 25978 25832 25984
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25700 24342 25728 25230
rect 25780 24948 25832 24954
rect 25780 24890 25832 24896
rect 25792 24750 25820 24890
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 25688 24336 25740 24342
rect 25688 24278 25740 24284
rect 25780 23656 25832 23662
rect 25780 23598 25832 23604
rect 25688 23520 25740 23526
rect 25688 23462 25740 23468
rect 25700 22030 25728 23462
rect 25792 23186 25820 23598
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25884 22094 25912 28426
rect 26148 28008 26200 28014
rect 26148 27950 26200 27956
rect 26160 27606 26188 27950
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 26068 25362 26096 26318
rect 26160 26314 26188 27338
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26252 25906 26280 28426
rect 27344 28416 27396 28422
rect 27344 28358 27396 28364
rect 27356 28218 27384 28358
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 26424 28144 26476 28150
rect 26424 28086 26476 28092
rect 26332 27396 26384 27402
rect 26332 27338 26384 27344
rect 26344 27062 26372 27338
rect 26332 27056 26384 27062
rect 26332 26998 26384 27004
rect 26332 26920 26384 26926
rect 26436 26908 26464 28086
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 26384 26880 26464 26908
rect 26332 26862 26384 26868
rect 26608 26852 26660 26858
rect 26608 26794 26660 26800
rect 26424 26784 26476 26790
rect 26424 26726 26476 26732
rect 26436 26314 26464 26726
rect 26620 26586 26648 26794
rect 26608 26580 26660 26586
rect 26608 26522 26660 26528
rect 26712 26518 26740 27270
rect 27632 27062 27660 28698
rect 27816 28218 27844 29514
rect 28276 28762 28304 30194
rect 29276 30048 29328 30054
rect 29276 29990 29328 29996
rect 29288 29238 29316 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 68100 29640 68152 29646
rect 68100 29582 68152 29588
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 68112 29345 68140 29582
rect 68098 29336 68154 29345
rect 68098 29271 68154 29280
rect 29276 29232 29328 29238
rect 29276 29174 29328 29180
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 28724 28960 28776 28966
rect 28724 28902 28776 28908
rect 28264 28756 28316 28762
rect 28264 28698 28316 28704
rect 28736 28558 28764 28902
rect 28172 28552 28224 28558
rect 28172 28494 28224 28500
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28908 28552 28960 28558
rect 28908 28494 28960 28500
rect 28184 28218 28212 28494
rect 28920 28218 28948 28494
rect 29000 28484 29052 28490
rect 29000 28426 29052 28432
rect 29012 28218 29040 28426
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28908 28212 28960 28218
rect 28908 28154 28960 28160
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 27712 27600 27764 27606
rect 27712 27542 27764 27548
rect 27620 27056 27672 27062
rect 27620 26998 27672 27004
rect 27724 26586 27752 27542
rect 27988 27532 28040 27538
rect 27988 27474 28040 27480
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 27724 26450 27752 26522
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 27066 26344 27122 26353
rect 26424 26308 26476 26314
rect 27066 26279 27068 26288
rect 26424 26250 26476 26256
rect 27120 26279 27122 26288
rect 27068 26250 27120 26256
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26056 25356 26108 25362
rect 26056 25298 26108 25304
rect 26252 24886 26280 25366
rect 26332 25220 26384 25226
rect 26332 25162 26384 25168
rect 26240 24880 26292 24886
rect 26240 24822 26292 24828
rect 26344 24750 26372 25162
rect 26332 24744 26384 24750
rect 26332 24686 26384 24692
rect 25884 22066 26004 22094
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25424 21434 25452 21490
rect 25332 21406 25452 21434
rect 25504 21412 25556 21418
rect 25332 20466 25360 21406
rect 25504 21354 25556 21360
rect 25412 20936 25464 20942
rect 25412 20878 25464 20884
rect 25424 20602 25452 20878
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25424 18426 25452 18702
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25516 17954 25544 21354
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25608 20058 25636 20402
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25424 17926 25544 17954
rect 25424 16425 25452 17926
rect 25504 17536 25556 17542
rect 25504 17478 25556 17484
rect 25410 16416 25466 16425
rect 25410 16351 25466 16360
rect 25226 14376 25282 14385
rect 25226 14311 25282 14320
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 25424 14006 25452 16351
rect 25516 14113 25544 17478
rect 25502 14104 25558 14113
rect 25502 14039 25558 14048
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24688 12714 24716 13194
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24964 12918 24992 13126
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 25056 12850 25084 13262
rect 25424 12850 25452 13942
rect 25504 13456 25556 13462
rect 25504 13398 25556 13404
rect 25044 12844 25096 12850
rect 25424 12844 25484 12850
rect 25424 12804 25432 12844
rect 25044 12786 25096 12792
rect 25432 12786 25484 12792
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24688 12442 24716 12650
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24582 11928 24638 11937
rect 24582 11863 24584 11872
rect 24636 11863 24638 11872
rect 24584 11834 24636 11840
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24122 11319 24178 11328
rect 24216 11348 24268 11354
rect 24032 11290 24084 11296
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 23860 10674 23888 11222
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 23952 11014 23980 11154
rect 24136 11082 24164 11319
rect 24216 11290 24268 11296
rect 24228 11150 24256 11290
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 23768 9586 23796 10610
rect 23952 10130 23980 10950
rect 23940 10124 23992 10130
rect 23940 10066 23992 10072
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 22926 8936 22982 8945
rect 22926 8871 22982 8880
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 23860 7002 23888 8502
rect 23952 8498 23980 10066
rect 24044 10062 24072 11018
rect 24688 10810 24716 11698
rect 24780 11150 24808 12174
rect 24964 11830 24992 12718
rect 25056 12306 25084 12786
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 25516 11898 25544 13398
rect 25608 12209 25636 19450
rect 25700 19378 25728 19858
rect 25976 19854 26004 22066
rect 26332 21072 26384 21078
rect 26332 21014 26384 21020
rect 26344 20398 26372 21014
rect 26332 20392 26384 20398
rect 26332 20334 26384 20340
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25700 18630 25728 19314
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25700 17678 25728 18566
rect 25780 18216 25832 18222
rect 25778 18184 25780 18193
rect 25832 18184 25834 18193
rect 25778 18119 25834 18128
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25780 17604 25832 17610
rect 25780 17546 25832 17552
rect 25792 17066 25820 17546
rect 25884 17338 25912 18022
rect 25964 17740 26016 17746
rect 25964 17682 26016 17688
rect 25976 17338 26004 17682
rect 26068 17678 26096 20198
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26160 19378 26188 19722
rect 26344 19378 26372 20334
rect 26436 20330 26464 26250
rect 27724 24818 27752 26386
rect 27804 26036 27856 26042
rect 27804 25978 27856 25984
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 27172 24410 27200 24754
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 27356 24070 27384 24754
rect 27528 24608 27580 24614
rect 27528 24550 27580 24556
rect 27540 24206 27568 24550
rect 27816 24274 27844 25978
rect 28000 25906 28028 27474
rect 28092 27470 28120 28018
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 28092 25974 28120 27406
rect 29104 27062 29132 29106
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 29196 27130 29224 28018
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 28172 27056 28224 27062
rect 28172 26998 28224 27004
rect 29092 27056 29144 27062
rect 29092 26998 29144 27004
rect 28080 25968 28132 25974
rect 28080 25910 28132 25916
rect 28184 25906 28212 26998
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 28172 25900 28224 25906
rect 28172 25842 28224 25848
rect 28184 25362 28212 25842
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 27804 24268 27856 24274
rect 27804 24210 27856 24216
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 26976 23792 27028 23798
rect 26976 23734 27028 23740
rect 26988 23186 27016 23734
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27172 23526 27200 23598
rect 27068 23520 27120 23526
rect 27068 23462 27120 23468
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 27080 23118 27108 23462
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 27356 22234 27384 24006
rect 27816 23798 27844 24210
rect 28368 24206 28396 24754
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 28184 23905 28212 24074
rect 28170 23896 28226 23905
rect 28170 23831 28172 23840
rect 28224 23831 28226 23840
rect 28172 23802 28224 23808
rect 27804 23792 27856 23798
rect 27804 23734 27856 23740
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 27632 21962 27660 22170
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 27436 21888 27488 21894
rect 27436 21830 27488 21836
rect 26988 21729 27016 21830
rect 26974 21720 27030 21729
rect 26974 21655 27030 21664
rect 27448 21622 27476 21830
rect 27436 21616 27488 21622
rect 27436 21558 27488 21564
rect 26514 20496 26570 20505
rect 26514 20431 26516 20440
rect 26568 20431 26570 20440
rect 26516 20402 26568 20408
rect 26424 20324 26476 20330
rect 26424 20266 26476 20272
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 26528 19553 26556 19654
rect 26514 19544 26570 19553
rect 26514 19479 26570 19488
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26160 18698 26188 19314
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26148 18148 26200 18154
rect 26148 18090 26200 18096
rect 26160 17678 26188 18090
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 25780 17060 25832 17066
rect 25780 17002 25832 17008
rect 25884 16232 25912 17274
rect 25792 16204 25912 16232
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25700 12986 25728 13194
rect 25792 12986 25820 16204
rect 25976 16130 26004 17274
rect 26252 17134 26280 17750
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 25884 16114 26004 16130
rect 25872 16108 26004 16114
rect 25924 16102 26004 16108
rect 25872 16050 25924 16056
rect 26436 15910 26464 16526
rect 26424 15904 26476 15910
rect 26424 15846 26476 15852
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26344 14346 26372 15438
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 26436 14006 26464 14758
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 26148 12708 26200 12714
rect 26148 12650 26200 12656
rect 26160 12238 26188 12650
rect 26620 12442 26648 19110
rect 26712 18766 26740 19314
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26700 18760 26752 18766
rect 26700 18702 26752 18708
rect 26712 17678 26740 18702
rect 26896 18698 26924 19246
rect 27448 18834 27476 21558
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27436 18828 27488 18834
rect 27436 18770 27488 18776
rect 27632 18766 27660 20878
rect 27816 20058 27844 23462
rect 28920 23322 28948 24210
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 29288 22094 29316 29174
rect 30840 29164 30892 29170
rect 30840 29106 30892 29112
rect 32496 29164 32548 29170
rect 32496 29106 32548 29112
rect 33508 29164 33560 29170
rect 33508 29106 33560 29112
rect 29920 29028 29972 29034
rect 29920 28970 29972 28976
rect 29368 28008 29420 28014
rect 29368 27950 29420 27956
rect 29380 27130 29408 27950
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 29932 26994 29960 28970
rect 30656 28688 30708 28694
rect 30656 28630 30708 28636
rect 30380 28552 30432 28558
rect 30564 28552 30616 28558
rect 30432 28512 30564 28540
rect 30380 28494 30432 28500
rect 30564 28494 30616 28500
rect 30472 28416 30524 28422
rect 30470 28384 30472 28393
rect 30524 28384 30526 28393
rect 30470 28319 30526 28328
rect 30378 28248 30434 28257
rect 30378 28183 30434 28192
rect 30392 28150 30420 28183
rect 30380 28144 30432 28150
rect 30380 28086 30432 28092
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30288 27464 30340 27470
rect 30288 27406 30340 27412
rect 30300 27130 30328 27406
rect 30288 27124 30340 27130
rect 30288 27066 30340 27072
rect 29920 26988 29972 26994
rect 29972 26948 30052 26976
rect 29920 26930 29972 26936
rect 29644 26920 29696 26926
rect 29644 26862 29696 26868
rect 29552 26240 29604 26246
rect 29552 26182 29604 26188
rect 29564 25974 29592 26182
rect 29552 25968 29604 25974
rect 29552 25910 29604 25916
rect 29552 25288 29604 25294
rect 29552 25230 29604 25236
rect 29460 24268 29512 24274
rect 29564 24256 29592 25230
rect 29512 24228 29592 24256
rect 29460 24210 29512 24216
rect 29564 23730 29592 24228
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29564 22778 29592 23054
rect 29552 22772 29604 22778
rect 29552 22714 29604 22720
rect 29288 22066 29408 22094
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 28000 20466 28028 21490
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 28184 19854 28212 21966
rect 28276 21690 28304 21966
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28460 20874 28488 21966
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28460 19922 28488 20810
rect 29288 20806 29316 21490
rect 29276 20800 29328 20806
rect 29276 20742 29328 20748
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28540 20256 28592 20262
rect 28540 20198 28592 20204
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28552 19854 28580 20198
rect 29012 20058 29040 20402
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 28172 19848 28224 19854
rect 28170 19816 28172 19825
rect 28540 19848 28592 19854
rect 28224 19816 28226 19825
rect 28540 19790 28592 19796
rect 28170 19751 28226 19760
rect 28816 19372 28868 19378
rect 28816 19314 28868 19320
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 26884 18692 26936 18698
rect 26884 18634 26936 18640
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27356 18290 27384 18566
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 26700 17672 26752 17678
rect 26700 17614 26752 17620
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26712 15502 26740 17614
rect 26804 17066 26832 17614
rect 26792 17060 26844 17066
rect 26792 17002 26844 17008
rect 26988 16114 27016 18226
rect 27160 17536 27212 17542
rect 27160 17478 27212 17484
rect 27172 16114 27200 17478
rect 27632 17270 27660 18702
rect 27804 18692 27856 18698
rect 27804 18634 27856 18640
rect 27816 18426 27844 18634
rect 27804 18420 27856 18426
rect 27804 18362 27856 18368
rect 28552 18290 28580 18702
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 27356 16114 27384 16934
rect 27632 16794 27660 17206
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27632 16674 27660 16730
rect 27540 16658 27660 16674
rect 27528 16652 27660 16658
rect 27580 16646 27660 16652
rect 27528 16594 27580 16600
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 26700 15496 26752 15502
rect 26988 15484 27016 16050
rect 27356 15706 27384 16050
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27068 15496 27120 15502
rect 26988 15456 27068 15484
rect 26700 15438 26752 15444
rect 27068 15438 27120 15444
rect 26700 15020 26752 15026
rect 26700 14962 26752 14968
rect 26712 14618 26740 14962
rect 26792 14952 26844 14958
rect 26792 14894 26844 14900
rect 26804 14618 26832 14894
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26804 13394 26832 14554
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 27172 12850 27200 13670
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26988 12306 27016 12786
rect 26976 12300 27028 12306
rect 26976 12242 27028 12248
rect 26148 12232 26200 12238
rect 25594 12200 25650 12209
rect 26148 12174 26200 12180
rect 25594 12135 25650 12144
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 26528 11830 26556 12038
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 26516 11824 26568 11830
rect 26516 11766 26568 11772
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24228 8498 24256 10406
rect 24688 10130 24716 10610
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24872 9178 24900 11630
rect 24964 10674 24992 11766
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25056 11529 25084 11698
rect 25042 11520 25098 11529
rect 25042 11455 25098 11464
rect 25700 11354 25728 11698
rect 25780 11688 25832 11694
rect 25976 11665 26004 11698
rect 26620 11694 26648 12038
rect 26988 11762 27016 12242
rect 27264 11898 27292 12786
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 26608 11688 26660 11694
rect 25780 11630 25832 11636
rect 25962 11656 26018 11665
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 23952 7478 23980 8434
rect 24504 8362 24532 8842
rect 24688 8566 24716 8910
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24780 8378 24808 8434
rect 24492 8356 24544 8362
rect 24780 8350 24900 8378
rect 24492 8298 24544 8304
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 23940 7472 23992 7478
rect 23940 7414 23992 7420
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23952 6798 23980 7414
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21364 6452 21416 6458
rect 21284 6412 21364 6440
rect 20904 6394 20956 6400
rect 21364 6394 21416 6400
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20916 5778 20944 6394
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 21008 6225 21036 6258
rect 20994 6216 21050 6225
rect 20994 6151 21050 6160
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 21652 5710 21680 6666
rect 23492 6322 23520 6734
rect 24688 6730 24716 7686
rect 24872 7410 24900 8350
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24780 6730 24808 7142
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 23020 5568 23072 5574
rect 23020 5510 23072 5516
rect 20824 4214 20852 5510
rect 23032 5370 23060 5510
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23492 5234 23520 6258
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23676 5234 23704 5850
rect 24228 5846 24256 6190
rect 24504 5914 24532 6258
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24216 5840 24268 5846
rect 24216 5782 24268 5788
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4214 20944 4966
rect 21192 4826 21220 5170
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21652 4282 21680 4626
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 23492 4214 23520 5170
rect 23676 4826 23704 5170
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 24228 4690 24256 5782
rect 24584 5704 24636 5710
rect 24780 5692 24808 6666
rect 24964 6458 24992 8910
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 25056 7750 25084 8230
rect 25148 7886 25176 8366
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25240 7818 25268 9998
rect 25332 7886 25360 11086
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25516 9110 25544 9454
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25516 8430 25544 9046
rect 25700 8838 25728 9998
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25700 8498 25728 8774
rect 25792 8634 25820 11630
rect 26608 11630 26660 11636
rect 25962 11591 26018 11600
rect 27356 10962 27384 15642
rect 27540 14958 27568 16594
rect 27724 16182 27752 18158
rect 28000 17542 28028 18226
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27816 16250 27844 17138
rect 28000 16794 28028 17478
rect 28552 17354 28580 18226
rect 28828 17882 28856 19314
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 29090 17776 29146 17785
rect 29090 17711 29146 17720
rect 29104 17678 29132 17711
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 29288 17610 29316 20742
rect 29380 17746 29408 22066
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29368 17740 29420 17746
rect 29368 17682 29420 17688
rect 29276 17604 29328 17610
rect 29276 17546 29328 17552
rect 28460 17326 28580 17354
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 27804 16244 27856 16250
rect 27804 16186 27856 16192
rect 27712 16176 27764 16182
rect 27712 16118 27764 16124
rect 27724 15434 27752 16118
rect 27712 15428 27764 15434
rect 27712 15370 27764 15376
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27540 14634 27568 14894
rect 27724 14890 27752 15370
rect 27712 14884 27764 14890
rect 27712 14826 27764 14832
rect 27448 14618 27568 14634
rect 27436 14612 27568 14618
rect 27488 14606 27568 14612
rect 27436 14554 27488 14560
rect 28000 14278 28028 16730
rect 28080 16516 28132 16522
rect 28080 16458 28132 16464
rect 28092 16250 28120 16458
rect 28460 16454 28488 17326
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29196 16522 29224 16934
rect 29472 16697 29500 17750
rect 29550 17640 29606 17649
rect 29550 17575 29606 17584
rect 29564 17542 29592 17575
rect 29552 17536 29604 17542
rect 29552 17478 29604 17484
rect 29552 16992 29604 16998
rect 29552 16934 29604 16940
rect 29458 16688 29514 16697
rect 29458 16623 29514 16632
rect 29564 16590 29592 16934
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29184 16516 29236 16522
rect 29184 16458 29236 16464
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28080 16244 28132 16250
rect 28080 16186 28132 16192
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28078 16144 28134 16153
rect 28078 16079 28134 16088
rect 28092 14414 28120 16079
rect 28184 15502 28212 16186
rect 28460 15978 28488 16390
rect 28448 15972 28500 15978
rect 28448 15914 28500 15920
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28184 14618 28212 15438
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 28276 15094 28304 15302
rect 28552 15162 28580 16390
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 28644 15366 28672 16118
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 28632 15360 28684 15366
rect 28630 15328 28632 15337
rect 28684 15328 28686 15337
rect 28630 15263 28686 15272
rect 28540 15156 28592 15162
rect 28540 15098 28592 15104
rect 28264 15088 28316 15094
rect 28264 15030 28316 15036
rect 28736 15026 28764 16050
rect 29092 15972 29144 15978
rect 29092 15914 29144 15920
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28736 14618 28764 14962
rect 28172 14612 28224 14618
rect 28172 14554 28224 14560
rect 28724 14612 28776 14618
rect 28724 14554 28776 14560
rect 28908 14544 28960 14550
rect 28908 14486 28960 14492
rect 28448 14476 28500 14482
rect 28448 14418 28500 14424
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27526 13424 27582 13433
rect 27526 13359 27582 13368
rect 27540 12782 27568 13359
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 27632 12986 27660 13194
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27434 12608 27490 12617
rect 27434 12543 27490 12552
rect 27448 11898 27476 12543
rect 27528 12436 27580 12442
rect 27528 12378 27580 12384
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27540 11762 27568 12378
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27632 11150 27660 11494
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27356 10934 27660 10962
rect 27528 10804 27580 10810
rect 27528 10746 27580 10752
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26712 10470 26740 10678
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26252 8974 26280 9998
rect 26608 9104 26660 9110
rect 26608 9046 26660 9052
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 26424 8560 26476 8566
rect 26424 8502 26476 8508
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 25504 8424 25556 8430
rect 25504 8366 25556 8372
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26068 7886 26096 8026
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 25228 7812 25280 7818
rect 25228 7754 25280 7760
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25056 6730 25084 7686
rect 25700 6798 25728 7686
rect 26252 7546 26280 7822
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 25688 6792 25740 6798
rect 25688 6734 25740 6740
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 24636 5664 24808 5692
rect 24584 5646 24636 5652
rect 24780 5370 24808 5664
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 25148 5234 25176 5646
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 24216 4684 24268 4690
rect 24216 4626 24268 4632
rect 25228 4548 25280 4554
rect 25228 4490 25280 4496
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20904 4208 20956 4214
rect 20904 4150 20956 4156
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 20824 4010 20852 4150
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20916 3913 20944 4150
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 20996 3936 21048 3942
rect 20902 3904 20958 3913
rect 20996 3878 21048 3884
rect 20902 3839 20958 3848
rect 20916 3194 20944 3839
rect 21008 3534 21036 3878
rect 21192 3738 21220 4082
rect 24688 3942 24716 4082
rect 25240 4078 25268 4490
rect 25424 4146 25452 6258
rect 25596 5772 25648 5778
rect 25596 5714 25648 5720
rect 25608 5370 25636 5714
rect 25700 5710 25728 6394
rect 26344 6322 26372 7414
rect 26436 7410 26464 8502
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26436 7002 26464 7346
rect 26424 6996 26476 7002
rect 26424 6938 26476 6944
rect 26332 6316 26384 6322
rect 26332 6258 26384 6264
rect 26344 5914 26372 6258
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25872 5636 25924 5642
rect 25872 5578 25924 5584
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25608 4146 25636 5306
rect 25884 5302 25912 5578
rect 25872 5296 25924 5302
rect 25872 5238 25924 5244
rect 25884 4554 25912 5238
rect 26528 4622 26556 8434
rect 26620 5302 26648 9046
rect 26712 5914 26740 10406
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27252 9988 27304 9994
rect 27252 9930 27304 9936
rect 27264 9450 27292 9930
rect 27252 9444 27304 9450
rect 27252 9386 27304 9392
rect 27356 9178 27384 10066
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 27540 9110 27568 10746
rect 27632 10538 27660 10934
rect 27620 10532 27672 10538
rect 27620 10474 27672 10480
rect 27528 9104 27580 9110
rect 27528 9046 27580 9052
rect 27632 9042 27660 10474
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27712 9512 27764 9518
rect 27712 9454 27764 9460
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27264 8498 27292 8842
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27252 8492 27304 8498
rect 27252 8434 27304 8440
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 26896 6458 26924 8026
rect 27264 7342 27292 8434
rect 27632 7478 27660 8774
rect 27724 8498 27752 9454
rect 27816 9178 27844 9522
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27724 7954 27752 8434
rect 27712 7948 27764 7954
rect 27712 7890 27764 7896
rect 27816 7886 27844 8978
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27620 7472 27672 7478
rect 27620 7414 27672 7420
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 27632 6662 27660 7414
rect 27816 7206 27844 7822
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 26884 6452 26936 6458
rect 26884 6394 26936 6400
rect 27908 5914 27936 13670
rect 28000 9586 28028 14214
rect 28092 13734 28120 14350
rect 28276 14249 28304 14350
rect 28262 14240 28318 14249
rect 28262 14175 28318 14184
rect 28460 13870 28488 14418
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 28644 13530 28672 13874
rect 28632 13524 28684 13530
rect 28684 13484 28764 13512
rect 28632 13466 28684 13472
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 28448 12436 28500 12442
rect 28448 12378 28500 12384
rect 28460 12186 28488 12378
rect 28644 12356 28672 12786
rect 28736 12434 28764 13484
rect 28920 12442 28948 14486
rect 28998 12744 29054 12753
rect 28998 12679 29054 12688
rect 28908 12436 28960 12442
rect 28736 12406 28856 12434
rect 28644 12328 28764 12356
rect 28368 12158 28488 12186
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28540 12164 28592 12170
rect 28368 10418 28396 12158
rect 28540 12106 28592 12112
rect 28552 11830 28580 12106
rect 28540 11824 28592 11830
rect 28540 11766 28592 11772
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28460 10606 28488 11698
rect 28552 11354 28580 11766
rect 28644 11762 28672 12174
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28540 11348 28592 11354
rect 28540 11290 28592 11296
rect 28448 10600 28500 10606
rect 28448 10542 28500 10548
rect 28368 10390 28488 10418
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 28092 8378 28120 9454
rect 28264 9376 28316 9382
rect 28264 9318 28316 9324
rect 28276 9042 28304 9318
rect 28368 9178 28396 9998
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28264 9036 28316 9042
rect 28264 8978 28316 8984
rect 28172 8424 28224 8430
rect 28092 8372 28172 8378
rect 28092 8366 28224 8372
rect 28460 8378 28488 10390
rect 28644 9994 28672 11698
rect 28632 9988 28684 9994
rect 28632 9930 28684 9936
rect 28644 9654 28672 9930
rect 28632 9648 28684 9654
rect 28632 9590 28684 9596
rect 28092 8350 28212 8366
rect 28460 8350 28580 8378
rect 27988 7880 28040 7886
rect 27988 7822 28040 7828
rect 28000 7546 28028 7822
rect 28092 7818 28120 8350
rect 28552 8090 28580 8350
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 27988 7540 28040 7546
rect 27988 7482 28040 7488
rect 28368 6798 28396 7686
rect 28552 7206 28580 8026
rect 28448 7200 28500 7206
rect 28448 7142 28500 7148
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28356 6792 28408 6798
rect 28356 6734 28408 6740
rect 28460 6361 28488 7142
rect 28632 6792 28684 6798
rect 28632 6734 28684 6740
rect 28446 6352 28502 6361
rect 27988 6316 28040 6322
rect 28446 6287 28502 6296
rect 27988 6258 28040 6264
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 27344 5908 27396 5914
rect 27344 5850 27396 5856
rect 27896 5908 27948 5914
rect 27896 5850 27948 5856
rect 26976 5636 27028 5642
rect 26976 5578 27028 5584
rect 26608 5296 26660 5302
rect 26608 5238 26660 5244
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 25872 4548 25924 4554
rect 25872 4490 25924 4496
rect 25688 4480 25740 4486
rect 25688 4422 25740 4428
rect 25700 4146 25728 4422
rect 26620 4282 26648 5238
rect 26988 5234 27016 5578
rect 27252 5568 27304 5574
rect 27252 5510 27304 5516
rect 27264 5370 27292 5510
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27356 5234 27384 5850
rect 27908 5778 27936 5850
rect 27896 5772 27948 5778
rect 27896 5714 27948 5720
rect 27896 5636 27948 5642
rect 27896 5578 27948 5584
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 26608 4276 26660 4282
rect 26608 4218 26660 4224
rect 26988 4146 27016 5170
rect 27356 5030 27384 5170
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27632 4214 27660 4966
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20588 2536 20668 2564
rect 20536 2518 20588 2524
rect 20732 800 20760 2790
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21008 800 21036 2382
rect 21284 800 21312 2926
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21560 800 21588 2790
rect 21744 2650 21772 2994
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21836 800 21864 3470
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21928 2514 21956 2586
rect 22100 2576 22152 2582
rect 22100 2518 22152 2524
rect 21916 2508 21968 2514
rect 21916 2450 21968 2456
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22020 2378 22048 2450
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 22112 800 22140 2518
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22388 800 22416 2382
rect 22664 800 22692 3470
rect 22928 2848 22980 2854
rect 22928 2790 22980 2796
rect 22940 800 22968 2790
rect 23204 2576 23256 2582
rect 23204 2518 23256 2524
rect 23216 800 23244 2518
rect 23492 800 23520 3470
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 23768 800 23796 2790
rect 24044 800 24072 2790
rect 24320 800 24348 3470
rect 24584 2372 24636 2378
rect 24584 2314 24636 2320
rect 24596 800 24624 2314
rect 24688 2038 24716 3878
rect 27908 3534 27936 5578
rect 28000 5370 28028 6258
rect 28644 6186 28672 6734
rect 28632 6180 28684 6186
rect 28632 6122 28684 6128
rect 28644 5846 28672 6122
rect 28356 5840 28408 5846
rect 28356 5782 28408 5788
rect 28632 5840 28684 5846
rect 28632 5782 28684 5788
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 27988 5364 28040 5370
rect 28184 5352 28212 5646
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 27988 5306 28040 5312
rect 28092 5324 28212 5352
rect 28092 5234 28120 5324
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28184 4554 28212 5170
rect 28172 4548 28224 4554
rect 28172 4490 28224 4496
rect 28276 3602 28304 5510
rect 28368 4146 28396 5782
rect 28736 5098 28764 12328
rect 28828 12322 28856 12406
rect 28908 12378 28960 12384
rect 28828 12306 28948 12322
rect 28828 12300 28960 12306
rect 28828 12294 28908 12300
rect 28908 12242 28960 12248
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28828 11762 28856 12174
rect 29012 11762 29040 12679
rect 29104 12646 29132 15914
rect 29552 15632 29604 15638
rect 29552 15574 29604 15580
rect 29564 15162 29592 15574
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 29656 13394 29684 26862
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 29748 23730 29776 26250
rect 29736 23724 29788 23730
rect 29736 23666 29788 23672
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29840 18970 29868 19314
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 29828 17876 29880 17882
rect 29828 17818 29880 17824
rect 29840 17678 29868 17818
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29828 17672 29880 17678
rect 29828 17614 29880 17620
rect 29748 17218 29776 17614
rect 29932 17610 29960 23054
rect 29920 17604 29972 17610
rect 29920 17546 29972 17552
rect 29748 17202 29868 17218
rect 29748 17196 29880 17202
rect 29748 17190 29828 17196
rect 29828 17138 29880 17144
rect 29840 16658 29868 17138
rect 29932 17134 29960 17546
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29828 16652 29880 16658
rect 29828 16594 29880 16600
rect 29932 16590 29960 17070
rect 30024 16590 30052 26948
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 30300 24138 30328 24754
rect 30288 24132 30340 24138
rect 30288 24074 30340 24080
rect 30300 23322 30328 24074
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30116 22710 30144 22918
rect 30104 22704 30156 22710
rect 30104 22646 30156 22652
rect 30116 22030 30144 22646
rect 30392 22094 30420 27950
rect 30576 27538 30604 28494
rect 30668 28218 30696 28630
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 30760 28393 30788 28494
rect 30746 28384 30802 28393
rect 30746 28319 30802 28328
rect 30852 28257 30880 29106
rect 32128 28960 32180 28966
rect 32128 28902 32180 28908
rect 30838 28248 30894 28257
rect 30656 28212 30708 28218
rect 30838 28183 30894 28192
rect 30656 28154 30708 28160
rect 32140 28150 32168 28902
rect 32508 28762 32536 29106
rect 32496 28756 32548 28762
rect 32496 28698 32548 28704
rect 32128 28144 32180 28150
rect 32128 28086 32180 28092
rect 33520 28082 33548 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 33508 28076 33560 28082
rect 33508 28018 33560 28024
rect 30564 27532 30616 27538
rect 30564 27474 30616 27480
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30760 26450 30788 27406
rect 30852 27062 30880 28018
rect 31024 27872 31076 27878
rect 31024 27814 31076 27820
rect 32128 27872 32180 27878
rect 32128 27814 32180 27820
rect 30840 27056 30892 27062
rect 30892 27016 30972 27044
rect 30840 26998 30892 27004
rect 30748 26444 30800 26450
rect 30748 26386 30800 26392
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 30668 25906 30696 26318
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 30760 25362 30788 26386
rect 30840 26376 30892 26382
rect 30840 26318 30892 26324
rect 30852 26042 30880 26318
rect 30840 26036 30892 26042
rect 30840 25978 30892 25984
rect 30944 25906 30972 27016
rect 31036 26790 31064 27814
rect 32140 27062 32168 27814
rect 32508 27606 32536 28018
rect 32496 27600 32548 27606
rect 32496 27542 32548 27548
rect 32128 27056 32180 27062
rect 32128 26998 32180 27004
rect 31024 26784 31076 26790
rect 31024 26726 31076 26732
rect 31036 26382 31064 26726
rect 33520 26450 33548 28018
rect 67638 27976 67694 27985
rect 67638 27911 67640 27920
rect 67692 27911 67694 27920
rect 67640 27882 67692 27888
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 67640 26784 67692 26790
rect 67640 26726 67692 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 67652 26625 67680 26726
rect 67638 26616 67694 26625
rect 67638 26551 67694 26560
rect 33508 26444 33560 26450
rect 33508 26386 33560 26392
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 30748 25356 30800 25362
rect 30748 25298 30800 25304
rect 30944 24954 30972 25842
rect 31220 25498 31248 26250
rect 31852 26240 31904 26246
rect 31852 26182 31904 26188
rect 31864 25906 31892 26182
rect 33520 26042 33548 26386
rect 34060 26376 34112 26382
rect 34060 26318 34112 26324
rect 33508 26036 33560 26042
rect 33508 25978 33560 25984
rect 31852 25900 31904 25906
rect 31852 25842 31904 25848
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32680 25900 32732 25906
rect 32680 25842 32732 25848
rect 32864 25900 32916 25906
rect 32864 25842 32916 25848
rect 31576 25696 31628 25702
rect 31576 25638 31628 25644
rect 31208 25492 31260 25498
rect 31208 25434 31260 25440
rect 31588 25226 31616 25638
rect 31576 25220 31628 25226
rect 31576 25162 31628 25168
rect 31760 25220 31812 25226
rect 31760 25162 31812 25168
rect 30932 24948 30984 24954
rect 30932 24890 30984 24896
rect 30564 24336 30616 24342
rect 30564 24278 30616 24284
rect 30576 24070 30604 24278
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 30472 23588 30524 23594
rect 30472 23530 30524 23536
rect 30484 22778 30512 23530
rect 30656 23044 30708 23050
rect 30656 22986 30708 22992
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30208 22066 30420 22094
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 30116 18290 30144 19314
rect 30104 18284 30156 18290
rect 30104 18226 30156 18232
rect 29920 16584 29972 16590
rect 29826 16552 29882 16561
rect 29920 16526 29972 16532
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 29826 16487 29828 16496
rect 29880 16487 29882 16496
rect 29828 16458 29880 16464
rect 29932 16114 29960 16526
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29840 13462 29868 15438
rect 29920 15360 29972 15366
rect 29920 15302 29972 15308
rect 29828 13456 29880 13462
rect 29828 13398 29880 13404
rect 29644 13388 29696 13394
rect 29644 13330 29696 13336
rect 29840 13326 29868 13398
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29828 13184 29880 13190
rect 29828 13126 29880 13132
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 28816 11756 28868 11762
rect 29000 11756 29052 11762
rect 28868 11716 28948 11744
rect 28816 11698 28868 11704
rect 28920 10130 28948 11716
rect 29000 11698 29052 11704
rect 29012 11354 29040 11698
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 29012 10266 29040 10542
rect 29000 10260 29052 10266
rect 29000 10202 29052 10208
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 28724 5092 28776 5098
rect 28724 5034 28776 5040
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 28356 4140 28408 4146
rect 28356 4082 28408 4088
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 28552 3534 28580 4422
rect 28736 4146 28764 5034
rect 29012 4622 29040 9862
rect 29104 8498 29132 12582
rect 29656 12238 29684 12718
rect 29840 12442 29868 13126
rect 29828 12436 29880 12442
rect 29828 12378 29880 12384
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29932 11354 29960 15302
rect 30116 15194 30144 18226
rect 30208 17202 30236 22066
rect 30668 21690 30696 22986
rect 31116 22432 31168 22438
rect 31116 22374 31168 22380
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 31128 21554 31156 22374
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31220 21622 31248 21898
rect 31208 21616 31260 21622
rect 31208 21558 31260 21564
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 31220 21078 31248 21558
rect 30656 21072 30708 21078
rect 30656 21014 30708 21020
rect 31208 21072 31260 21078
rect 31208 21014 31260 21020
rect 30288 21004 30340 21010
rect 30288 20946 30340 20952
rect 30300 20806 30328 20946
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30668 19446 30696 21014
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31128 19786 31156 20878
rect 31116 19780 31168 19786
rect 31116 19722 31168 19728
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 30748 19712 30800 19718
rect 30748 19654 30800 19660
rect 30656 19440 30708 19446
rect 30656 19382 30708 19388
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30300 18290 30328 19110
rect 30668 18902 30696 19382
rect 30760 19378 30788 19654
rect 30748 19372 30800 19378
rect 30748 19314 30800 19320
rect 31128 18902 31156 19722
rect 31220 19514 31248 19722
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 30656 18896 30708 18902
rect 30656 18838 30708 18844
rect 31116 18896 31168 18902
rect 31116 18838 31168 18844
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30392 18154 30420 18770
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30748 18692 30800 18698
rect 30748 18634 30800 18640
rect 30760 18426 30788 18634
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30196 16448 30248 16454
rect 30196 16390 30248 16396
rect 30208 15570 30236 16390
rect 30300 15978 30328 18022
rect 30852 17785 30880 18702
rect 30838 17776 30894 17785
rect 30838 17711 30894 17720
rect 30840 17536 30892 17542
rect 30840 17478 30892 17484
rect 30852 17270 30880 17478
rect 30840 17264 30892 17270
rect 30840 17206 30892 17212
rect 30380 16720 30432 16726
rect 30380 16662 30432 16668
rect 30654 16688 30710 16697
rect 30288 15972 30340 15978
rect 30288 15914 30340 15920
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30392 15484 30420 16662
rect 30654 16623 30710 16632
rect 30472 15496 30524 15502
rect 30392 15456 30472 15484
rect 30116 15166 30328 15194
rect 30300 13870 30328 15166
rect 30392 15162 30420 15456
rect 30472 15438 30524 15444
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30484 14482 30512 15302
rect 30472 14476 30524 14482
rect 30392 14436 30472 14464
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 30288 13456 30340 13462
rect 30288 13398 30340 13404
rect 30010 13288 30066 13297
rect 30010 13223 30012 13232
rect 30064 13223 30066 13232
rect 30012 13194 30064 13200
rect 30300 12850 30328 13398
rect 30392 13258 30420 14436
rect 30472 14418 30524 14424
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30472 13320 30524 13326
rect 30472 13262 30524 13268
rect 30380 13252 30432 13258
rect 30380 13194 30432 13200
rect 30392 12918 30420 13194
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30380 12640 30432 12646
rect 30380 12582 30432 12588
rect 30286 12472 30342 12481
rect 30286 12407 30288 12416
rect 30340 12407 30342 12416
rect 30288 12378 30340 12384
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 29644 11280 29696 11286
rect 29642 11248 29644 11257
rect 29696 11248 29698 11257
rect 29642 11183 29698 11192
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29564 10577 29592 10610
rect 29550 10568 29606 10577
rect 29550 10503 29606 10512
rect 29932 10266 29960 11086
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 30024 10713 30052 10746
rect 30010 10704 30066 10713
rect 30010 10639 30066 10648
rect 30392 10470 30420 12582
rect 30380 10464 30432 10470
rect 30380 10406 30432 10412
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29368 9988 29420 9994
rect 29368 9930 29420 9936
rect 29380 8634 29408 9930
rect 29368 8628 29420 8634
rect 29368 8570 29420 8576
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 29104 8090 29132 8434
rect 29092 8084 29144 8090
rect 29092 8026 29144 8032
rect 29104 7546 29132 8026
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 29472 5914 29500 9998
rect 29736 9988 29788 9994
rect 29736 9930 29788 9936
rect 29748 9654 29776 9930
rect 29736 9648 29788 9654
rect 29736 9590 29788 9596
rect 29552 9104 29604 9110
rect 29604 9052 29684 9058
rect 29552 9046 29684 9052
rect 29564 9030 29684 9046
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29564 6798 29592 8910
rect 29656 8634 29684 9030
rect 29840 8838 29868 9998
rect 29828 8832 29880 8838
rect 29828 8774 29880 8780
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 30484 8022 30512 13262
rect 30576 10198 30604 14214
rect 30668 11898 30696 16623
rect 30852 16182 30880 17206
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30944 16114 30972 16526
rect 31312 16114 31340 24006
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31392 22092 31444 22098
rect 31392 22034 31444 22040
rect 31404 21894 31432 22034
rect 31392 21888 31444 21894
rect 31392 21830 31444 21836
rect 31404 21554 31432 21830
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31404 21010 31432 21490
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 31404 20534 31432 20946
rect 31392 20528 31444 20534
rect 31392 20470 31444 20476
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30760 15745 30788 15846
rect 30746 15736 30802 15745
rect 30746 15671 30802 15680
rect 30944 15026 30972 16050
rect 31208 16040 31260 16046
rect 31208 15982 31260 15988
rect 31220 15026 31248 15982
rect 31496 15026 31524 23666
rect 30748 15020 30800 15026
rect 30748 14962 30800 14968
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31484 15020 31536 15026
rect 31484 14962 31536 14968
rect 30760 13938 30788 14962
rect 30932 14884 30984 14890
rect 30932 14826 30984 14832
rect 30840 14816 30892 14822
rect 30840 14758 30892 14764
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 30760 13326 30788 13874
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 30656 11892 30708 11898
rect 30656 11834 30708 11840
rect 30668 11694 30696 11834
rect 30852 11830 30880 14758
rect 30840 11824 30892 11830
rect 30840 11766 30892 11772
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30668 10810 30696 11630
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30668 10470 30696 10746
rect 30656 10464 30708 10470
rect 30656 10406 30708 10412
rect 30564 10192 30616 10198
rect 30564 10134 30616 10140
rect 30944 8514 30972 14826
rect 31220 14414 31248 14962
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31404 13938 31432 14350
rect 31588 13938 31616 25162
rect 31772 24682 31800 25162
rect 31760 24676 31812 24682
rect 31760 24618 31812 24624
rect 31668 24132 31720 24138
rect 31668 24074 31720 24080
rect 31680 23730 31708 24074
rect 31772 23866 31800 24618
rect 31760 23860 31812 23866
rect 31760 23802 31812 23808
rect 31668 23724 31720 23730
rect 31668 23666 31720 23672
rect 31668 22636 31720 22642
rect 31668 22578 31720 22584
rect 31680 21622 31708 22578
rect 31760 22024 31812 22030
rect 31760 21966 31812 21972
rect 31668 21616 31720 21622
rect 31668 21558 31720 21564
rect 31680 20942 31708 21558
rect 31668 20936 31720 20942
rect 31668 20878 31720 20884
rect 31772 20466 31800 21966
rect 31760 20460 31812 20466
rect 31760 20402 31812 20408
rect 31864 14498 31892 25842
rect 32508 24818 32536 25842
rect 32692 25498 32720 25842
rect 32680 25492 32732 25498
rect 32680 25434 32732 25440
rect 32680 25220 32732 25226
rect 32680 25162 32732 25168
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32508 24698 32536 24754
rect 32416 24670 32536 24698
rect 31944 24200 31996 24206
rect 31944 24142 31996 24148
rect 31956 23186 31984 24142
rect 32220 24064 32272 24070
rect 32220 24006 32272 24012
rect 32128 23656 32180 23662
rect 32128 23598 32180 23604
rect 31944 23180 31996 23186
rect 31944 23122 31996 23128
rect 32140 23050 32168 23598
rect 32232 23594 32260 24006
rect 32416 23730 32444 24670
rect 32496 23860 32548 23866
rect 32496 23802 32548 23808
rect 32508 23746 32536 23802
rect 32404 23724 32456 23730
rect 32324 23684 32404 23712
rect 32220 23588 32272 23594
rect 32220 23530 32272 23536
rect 32324 23474 32352 23684
rect 32508 23718 32628 23746
rect 32404 23666 32456 23672
rect 32600 23526 32628 23718
rect 32232 23446 32352 23474
rect 32404 23520 32456 23526
rect 32404 23462 32456 23468
rect 32588 23520 32640 23526
rect 32588 23462 32640 23468
rect 32232 23118 32260 23446
rect 32416 23118 32444 23462
rect 32220 23112 32272 23118
rect 32220 23054 32272 23060
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32588 23112 32640 23118
rect 32588 23054 32640 23060
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 32600 22778 32628 23054
rect 32588 22772 32640 22778
rect 32588 22714 32640 22720
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 32048 22030 32076 22374
rect 32404 22092 32456 22098
rect 32692 22094 32720 25162
rect 32876 24954 32904 25842
rect 32956 25832 33008 25838
rect 32956 25774 33008 25780
rect 32864 24948 32916 24954
rect 32864 24890 32916 24896
rect 32968 24854 32996 25774
rect 33140 25696 33192 25702
rect 33140 25638 33192 25644
rect 33152 25294 33180 25638
rect 33140 25288 33192 25294
rect 33140 25230 33192 25236
rect 32876 24826 32996 24854
rect 32876 24750 32904 24826
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33416 24812 33468 24818
rect 33416 24754 33468 24760
rect 32864 24744 32916 24750
rect 32864 24686 32916 24692
rect 32772 24132 32824 24138
rect 32772 24074 32824 24080
rect 32784 23526 32812 24074
rect 32876 23798 32904 24686
rect 32956 24608 33008 24614
rect 32956 24550 33008 24556
rect 32968 24138 32996 24550
rect 33152 24410 33180 24754
rect 33140 24404 33192 24410
rect 33140 24346 33192 24352
rect 33428 24342 33456 24754
rect 33416 24336 33468 24342
rect 33416 24278 33468 24284
rect 32956 24132 33008 24138
rect 32956 24074 33008 24080
rect 32864 23792 32916 23798
rect 32864 23734 32916 23740
rect 32968 23610 32996 24074
rect 33692 23860 33744 23866
rect 33692 23802 33744 23808
rect 33784 23860 33836 23866
rect 33784 23802 33836 23808
rect 32876 23582 32996 23610
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 32784 23118 32812 23462
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 32692 22066 32812 22094
rect 32404 22034 32456 22040
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 31944 20868 31996 20874
rect 31944 20810 31996 20816
rect 31956 20602 31984 20810
rect 32232 20806 32260 21966
rect 32416 21894 32444 22034
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 31944 20596 31996 20602
rect 31944 20538 31996 20544
rect 31944 20256 31996 20262
rect 31944 20198 31996 20204
rect 31956 18834 31984 20198
rect 32232 20058 32260 20742
rect 32404 20460 32456 20466
rect 32404 20402 32456 20408
rect 32220 20052 32272 20058
rect 32220 19994 32272 20000
rect 32416 19854 32444 20402
rect 32404 19848 32456 19854
rect 32404 19790 32456 19796
rect 31944 18828 31996 18834
rect 31944 18770 31996 18776
rect 32416 18766 32444 19790
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32404 18760 32456 18766
rect 32404 18702 32456 18708
rect 32232 17746 32260 18702
rect 32600 18426 32628 21626
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 32312 17808 32364 17814
rect 32312 17750 32364 17756
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32324 17338 32352 17750
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32416 17338 32444 17478
rect 32312 17332 32364 17338
rect 32312 17274 32364 17280
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 32048 17066 32076 17138
rect 32036 17060 32088 17066
rect 32036 17002 32088 17008
rect 32232 16658 32260 17138
rect 32312 17128 32364 17134
rect 32364 17088 32444 17116
rect 32312 17070 32364 17076
rect 32310 16688 32366 16697
rect 32220 16652 32272 16658
rect 32310 16623 32366 16632
rect 32220 16594 32272 16600
rect 32324 16590 32352 16623
rect 32312 16584 32364 16590
rect 32312 16526 32364 16532
rect 32312 15904 32364 15910
rect 32312 15846 32364 15852
rect 32324 15502 32352 15846
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 32324 15094 32352 15438
rect 32312 15088 32364 15094
rect 32312 15030 32364 15036
rect 31864 14470 31984 14498
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 31392 13932 31444 13938
rect 31392 13874 31444 13880
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31024 13728 31076 13734
rect 31024 13670 31076 13676
rect 31036 12102 31064 13670
rect 31864 13462 31892 14350
rect 31852 13456 31904 13462
rect 31852 13398 31904 13404
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31864 12866 31892 12922
rect 31772 12838 31892 12866
rect 31772 12714 31800 12838
rect 31956 12782 31984 14470
rect 32312 13456 32364 13462
rect 32312 13398 32364 13404
rect 32324 12850 32352 13398
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 31944 12776 31996 12782
rect 31944 12718 31996 12724
rect 31760 12708 31812 12714
rect 31760 12650 31812 12656
rect 31392 12640 31444 12646
rect 31392 12582 31444 12588
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31024 12096 31076 12102
rect 31024 12038 31076 12044
rect 31128 11354 31156 12174
rect 31300 11756 31352 11762
rect 31300 11698 31352 11704
rect 31312 11354 31340 11698
rect 31404 11626 31432 12582
rect 32416 12374 32444 17088
rect 32600 15881 32628 18362
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 32586 15872 32642 15881
rect 32586 15807 32642 15816
rect 32600 13462 32628 15807
rect 32692 14822 32720 16050
rect 32784 15434 32812 22066
rect 32876 17354 32904 23582
rect 33416 23520 33468 23526
rect 33416 23462 33468 23468
rect 33428 23050 33456 23462
rect 33704 23322 33732 23802
rect 33692 23316 33744 23322
rect 33692 23258 33744 23264
rect 33796 23254 33824 23802
rect 33784 23248 33836 23254
rect 33784 23190 33836 23196
rect 33416 23044 33468 23050
rect 33416 22986 33468 22992
rect 32956 22432 33008 22438
rect 32956 22374 33008 22380
rect 32968 22094 32996 22374
rect 32968 22066 33364 22094
rect 32968 21418 32996 22066
rect 33336 22030 33364 22066
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 33152 21690 33180 21966
rect 33140 21684 33192 21690
rect 33140 21626 33192 21632
rect 32956 21412 33008 21418
rect 32956 21354 33008 21360
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 32968 20262 32996 20878
rect 33232 20800 33284 20806
rect 33232 20742 33284 20748
rect 33244 20466 33272 20742
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 32956 20256 33008 20262
rect 32956 20198 33008 20204
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 32876 17326 32996 17354
rect 32864 17196 32916 17202
rect 32864 17138 32916 17144
rect 32876 16794 32904 17138
rect 32864 16788 32916 16794
rect 32864 16730 32916 16736
rect 32772 15428 32824 15434
rect 32772 15370 32824 15376
rect 32968 15178 32996 17326
rect 33232 16516 33284 16522
rect 33232 16458 33284 16464
rect 33244 16402 33272 16458
rect 32784 15150 32996 15178
rect 33152 16374 33272 16402
rect 32680 14816 32732 14822
rect 32680 14758 32732 14764
rect 32588 13456 32640 13462
rect 32588 13398 32640 13404
rect 32404 12368 32456 12374
rect 32404 12310 32456 12316
rect 31392 11620 31444 11626
rect 31392 11562 31444 11568
rect 31390 11384 31446 11393
rect 31116 11348 31168 11354
rect 31116 11290 31168 11296
rect 31300 11348 31352 11354
rect 31390 11319 31446 11328
rect 31300 11290 31352 11296
rect 31024 11280 31076 11286
rect 31024 11222 31076 11228
rect 30760 8486 30972 8514
rect 30472 8016 30524 8022
rect 30472 7958 30524 7964
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30300 7018 30328 7142
rect 30300 6990 30420 7018
rect 29552 6792 29604 6798
rect 29552 6734 29604 6740
rect 30392 6322 30420 6990
rect 30760 6798 30788 8486
rect 30932 8424 30984 8430
rect 30932 8366 30984 8372
rect 30944 6798 30972 8366
rect 31036 8090 31064 11222
rect 31404 11150 31432 11319
rect 31666 11248 31722 11257
rect 31666 11183 31722 11192
rect 32128 11212 32180 11218
rect 31680 11150 31708 11183
rect 32128 11154 32180 11160
rect 31208 11144 31260 11150
rect 31208 11086 31260 11092
rect 31392 11144 31444 11150
rect 31392 11086 31444 11092
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31220 10674 31248 11086
rect 31576 11076 31628 11082
rect 31576 11018 31628 11024
rect 31392 11008 31444 11014
rect 31392 10950 31444 10956
rect 31404 10742 31432 10950
rect 31392 10736 31444 10742
rect 31392 10678 31444 10684
rect 31208 10668 31260 10674
rect 31208 10610 31260 10616
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 31312 10198 31340 10610
rect 31300 10192 31352 10198
rect 31300 10134 31352 10140
rect 31404 10044 31432 10678
rect 31588 10538 31616 11018
rect 32140 10810 32168 11154
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 32220 10668 32272 10674
rect 32220 10610 32272 10616
rect 31576 10532 31628 10538
rect 31576 10474 31628 10480
rect 31588 10062 31616 10474
rect 31312 10016 31432 10044
rect 31576 10056 31628 10062
rect 31312 9518 31340 10016
rect 31576 9998 31628 10004
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 31312 9042 31340 9454
rect 31300 9036 31352 9042
rect 31300 8978 31352 8984
rect 31588 8974 31616 9998
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 31024 7948 31076 7954
rect 31024 7890 31076 7896
rect 31036 7478 31064 7890
rect 31024 7472 31076 7478
rect 31076 7432 31156 7460
rect 31024 7414 31076 7420
rect 31024 7200 31076 7206
rect 31024 7142 31076 7148
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30932 6792 30984 6798
rect 30932 6734 30984 6740
rect 30564 6724 30616 6730
rect 30564 6666 30616 6672
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29472 5302 29500 5850
rect 29460 5296 29512 5302
rect 29460 5238 29512 5244
rect 30484 5098 30512 6598
rect 30576 6458 30604 6666
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 30760 5914 30788 6734
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 30748 5908 30800 5914
rect 30748 5850 30800 5856
rect 30472 5092 30524 5098
rect 30472 5034 30524 5040
rect 30760 4826 30788 5850
rect 30748 4820 30800 4826
rect 30748 4762 30800 4768
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29012 4282 29040 4558
rect 30852 4554 30880 6258
rect 30944 5778 30972 6734
rect 31036 6322 31064 7142
rect 31128 7002 31156 7432
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31116 6996 31168 7002
rect 31116 6938 31168 6944
rect 31404 6730 31432 7346
rect 31392 6724 31444 6730
rect 31392 6666 31444 6672
rect 31024 6316 31076 6322
rect 31024 6258 31076 6264
rect 30932 5772 30984 5778
rect 30932 5714 30984 5720
rect 30944 5302 30972 5714
rect 31300 5568 31352 5574
rect 31300 5510 31352 5516
rect 30932 5296 30984 5302
rect 30932 5238 30984 5244
rect 31312 5234 31340 5510
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 30840 4548 30892 4554
rect 30840 4490 30892 4496
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 31496 4214 31524 8842
rect 31576 8560 31628 8566
rect 31576 8502 31628 8508
rect 31588 6730 31616 8502
rect 31760 8492 31812 8498
rect 31760 8434 31812 8440
rect 31668 7880 31720 7886
rect 31772 7868 31800 8434
rect 31720 7840 31800 7868
rect 31668 7822 31720 7828
rect 31852 7812 31904 7818
rect 31852 7754 31904 7760
rect 31864 7274 31892 7754
rect 31956 7478 31984 8910
rect 31944 7472 31996 7478
rect 31944 7414 31996 7420
rect 31852 7268 31904 7274
rect 31852 7210 31904 7216
rect 31576 6724 31628 6730
rect 31576 6666 31628 6672
rect 32232 6662 32260 10610
rect 32312 10056 32364 10062
rect 32312 9998 32364 10004
rect 32324 8974 32352 9998
rect 32416 9722 32444 12310
rect 32692 12306 32720 14758
rect 32784 12714 32812 15150
rect 32956 15020 33008 15026
rect 32956 14962 33008 14968
rect 32968 14006 32996 14962
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 33060 14074 33088 14554
rect 33152 14550 33180 16374
rect 33336 15337 33364 17614
rect 33322 15328 33378 15337
rect 33322 15263 33378 15272
rect 33140 14544 33192 14550
rect 33140 14486 33192 14492
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 33048 14068 33100 14074
rect 33048 14010 33100 14016
rect 32956 14000 33008 14006
rect 32956 13942 33008 13948
rect 33048 13932 33100 13938
rect 33152 13920 33180 14350
rect 33324 14340 33376 14346
rect 33324 14282 33376 14288
rect 33336 13938 33364 14282
rect 33428 14278 33456 22986
rect 33508 22636 33560 22642
rect 33508 22578 33560 22584
rect 33520 21690 33548 22578
rect 33968 21888 34020 21894
rect 33968 21830 34020 21836
rect 33508 21684 33560 21690
rect 33508 21626 33560 21632
rect 33980 21622 34008 21830
rect 33968 21616 34020 21622
rect 33968 21558 34020 21564
rect 34072 21146 34100 26318
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 34428 26036 34480 26042
rect 34428 25978 34480 25984
rect 34440 25362 34468 25978
rect 34704 25900 34756 25906
rect 34704 25842 34756 25848
rect 34428 25356 34480 25362
rect 34428 25298 34480 25304
rect 34440 24818 34468 25298
rect 34716 25158 34744 25842
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 68100 25288 68152 25294
rect 68098 25256 68100 25265
rect 68152 25256 68154 25265
rect 68098 25191 68154 25200
rect 34704 25152 34756 25158
rect 34704 25094 34756 25100
rect 34428 24812 34480 24818
rect 34428 24754 34480 24760
rect 34440 24206 34468 24754
rect 34428 24200 34480 24206
rect 34428 24142 34480 24148
rect 34440 23798 34468 24142
rect 34428 23792 34480 23798
rect 34428 23734 34480 23740
rect 34336 22024 34388 22030
rect 34336 21966 34388 21972
rect 34520 22024 34572 22030
rect 34520 21966 34572 21972
rect 34348 21554 34376 21966
rect 34336 21548 34388 21554
rect 34336 21490 34388 21496
rect 34532 21350 34560 21966
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 34060 21140 34112 21146
rect 34060 21082 34112 21088
rect 34428 21004 34480 21010
rect 34428 20946 34480 20952
rect 33968 19168 34020 19174
rect 33968 19110 34020 19116
rect 33980 18698 34008 19110
rect 34244 18760 34296 18766
rect 34244 18702 34296 18708
rect 33968 18692 34020 18698
rect 33968 18634 34020 18640
rect 33980 17882 34008 18634
rect 34060 18624 34112 18630
rect 34060 18566 34112 18572
rect 34072 18154 34100 18566
rect 34256 18426 34284 18702
rect 34244 18420 34296 18426
rect 34244 18362 34296 18368
rect 34440 18358 34468 20946
rect 34532 20466 34560 21286
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34532 19446 34560 20402
rect 34520 19440 34572 19446
rect 34520 19382 34572 19388
rect 34428 18352 34480 18358
rect 34428 18294 34480 18300
rect 34060 18148 34112 18154
rect 34060 18090 34112 18096
rect 33968 17876 34020 17882
rect 33968 17818 34020 17824
rect 33876 17672 33928 17678
rect 33876 17614 33928 17620
rect 33888 17338 33916 17614
rect 33876 17332 33928 17338
rect 33876 17274 33928 17280
rect 33968 16448 34020 16454
rect 33968 16390 34020 16396
rect 33980 16250 34008 16390
rect 33968 16244 34020 16250
rect 33968 16186 34020 16192
rect 33782 15328 33838 15337
rect 33782 15263 33838 15272
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 33100 13892 33180 13920
rect 33324 13932 33376 13938
rect 33048 13874 33100 13880
rect 33324 13874 33376 13880
rect 33600 13932 33652 13938
rect 33600 13874 33652 13880
rect 32864 13796 32916 13802
rect 32864 13738 32916 13744
rect 32876 13530 32904 13738
rect 32864 13524 32916 13530
rect 32864 13466 32916 13472
rect 33060 13326 33088 13874
rect 33048 13320 33100 13326
rect 33100 13280 33180 13308
rect 33048 13262 33100 13268
rect 33048 13184 33100 13190
rect 33048 13126 33100 13132
rect 33060 12714 33088 13126
rect 32772 12708 32824 12714
rect 32772 12650 32824 12656
rect 33048 12708 33100 12714
rect 33048 12650 33100 12656
rect 32956 12368 33008 12374
rect 32956 12310 33008 12316
rect 32680 12300 32732 12306
rect 32680 12242 32732 12248
rect 32968 12102 32996 12310
rect 32956 12096 33008 12102
rect 32956 12038 33008 12044
rect 33060 11830 33088 12650
rect 33152 12374 33180 13280
rect 33336 13258 33364 13874
rect 33416 13456 33468 13462
rect 33416 13398 33468 13404
rect 33324 13252 33376 13258
rect 33324 13194 33376 13200
rect 33140 12368 33192 12374
rect 33140 12310 33192 12316
rect 33152 11898 33180 12310
rect 33140 11892 33192 11898
rect 33140 11834 33192 11840
rect 33048 11824 33100 11830
rect 33048 11766 33100 11772
rect 32680 11144 32732 11150
rect 32680 11086 32732 11092
rect 32496 11076 32548 11082
rect 32496 11018 32548 11024
rect 32508 10742 32536 11018
rect 32496 10736 32548 10742
rect 32496 10678 32548 10684
rect 32692 9722 32720 11086
rect 33152 10130 33180 11834
rect 33336 10674 33364 13194
rect 33428 12238 33456 13398
rect 33612 12442 33640 13874
rect 33600 12436 33652 12442
rect 33796 12434 33824 15263
rect 33600 12378 33652 12384
rect 33704 12406 33824 12434
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33612 11830 33640 12378
rect 33600 11824 33652 11830
rect 33600 11766 33652 11772
rect 33416 11756 33468 11762
rect 33416 11698 33468 11704
rect 33428 11150 33456 11698
rect 33416 11144 33468 11150
rect 33416 11086 33468 11092
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 33140 10124 33192 10130
rect 33140 10066 33192 10072
rect 32404 9716 32456 9722
rect 32404 9658 32456 9664
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 33336 9586 33364 10610
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 32588 9512 32640 9518
rect 32588 9454 32640 9460
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 32494 8936 32550 8945
rect 32324 8498 32352 8910
rect 32494 8871 32550 8880
rect 32508 8838 32536 8871
rect 32600 8838 32628 9454
rect 33704 9178 33732 12406
rect 34072 9586 34100 18090
rect 34440 17814 34468 18294
rect 34624 17882 34652 20878
rect 34716 20466 34744 25094
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 68100 24200 68152 24206
rect 68100 24142 68152 24148
rect 36728 24064 36780 24070
rect 36728 24006 36780 24012
rect 36740 23866 36768 24006
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 68112 23905 68140 24142
rect 68098 23896 68154 23905
rect 36728 23860 36780 23866
rect 68098 23831 68154 23840
rect 36728 23802 36780 23808
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 37372 22636 37424 22642
rect 37372 22578 37424 22584
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 37384 22094 37412 22578
rect 37384 22066 37504 22094
rect 37476 22030 37504 22066
rect 37464 22024 37516 22030
rect 37464 21966 37516 21972
rect 34888 21888 34940 21894
rect 34888 21830 34940 21836
rect 34900 21690 34928 21830
rect 34888 21684 34940 21690
rect 34888 21626 34940 21632
rect 37476 21554 37504 21966
rect 37568 21690 37596 22578
rect 67638 22536 67694 22545
rect 67638 22471 67640 22480
rect 67692 22471 67694 22480
rect 67640 22442 67692 22448
rect 38660 22432 38712 22438
rect 38660 22374 38712 22380
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 35992 21548 36044 21554
rect 35992 21490 36044 21496
rect 36176 21548 36228 21554
rect 36176 21490 36228 21496
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 37464 21548 37516 21554
rect 37464 21490 37516 21496
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 36004 20942 36032 21490
rect 36188 21146 36216 21490
rect 36176 21140 36228 21146
rect 36176 21082 36228 21088
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 36280 20874 36308 21490
rect 37188 20936 37240 20942
rect 37188 20878 37240 20884
rect 37372 20936 37424 20942
rect 37372 20878 37424 20884
rect 36268 20868 36320 20874
rect 36268 20810 36320 20816
rect 36084 20800 36136 20806
rect 36084 20742 36136 20748
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34716 20058 34744 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34704 20052 34756 20058
rect 34704 19994 34756 20000
rect 34612 17876 34664 17882
rect 34612 17818 34664 17824
rect 34428 17808 34480 17814
rect 34428 17750 34480 17756
rect 34336 17672 34388 17678
rect 34336 17614 34388 17620
rect 34348 17202 34376 17614
rect 34336 17196 34388 17202
rect 34336 17138 34388 17144
rect 34152 16992 34204 16998
rect 34152 16934 34204 16940
rect 34164 16590 34192 16934
rect 34152 16584 34204 16590
rect 34152 16526 34204 16532
rect 34164 15502 34192 16526
rect 34612 16108 34664 16114
rect 34612 16050 34664 16056
rect 34624 15706 34652 16050
rect 34612 15700 34664 15706
rect 34612 15642 34664 15648
rect 34716 15570 34744 19994
rect 35532 19984 35584 19990
rect 35532 19926 35584 19932
rect 35544 19446 35572 19926
rect 36096 19854 36124 20742
rect 36174 20632 36230 20641
rect 36174 20567 36230 20576
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 35532 19440 35584 19446
rect 35532 19382 35584 19388
rect 34888 19372 34940 19378
rect 34888 19314 34940 19320
rect 34900 19258 34928 19314
rect 34808 19230 34928 19258
rect 34808 18970 34836 19230
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34796 18964 34848 18970
rect 34796 18906 34848 18912
rect 35072 18964 35124 18970
rect 35072 18906 35124 18912
rect 35084 18766 35112 18906
rect 35069 18760 35121 18766
rect 35069 18702 35121 18708
rect 35084 18290 35112 18702
rect 35072 18284 35124 18290
rect 35072 18226 35124 18232
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34808 17542 34836 18158
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 34808 17202 34836 17478
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15564 34756 15570
rect 34704 15506 34756 15512
rect 34152 15496 34204 15502
rect 34152 15438 34204 15444
rect 34612 15360 34664 15366
rect 34612 15302 34664 15308
rect 34624 14890 34652 15302
rect 34716 15094 34744 15506
rect 34704 15088 34756 15094
rect 34704 15030 34756 15036
rect 35348 15088 35400 15094
rect 35348 15030 35400 15036
rect 34612 14884 34664 14890
rect 34612 14826 34664 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 34624 14006 34652 14282
rect 34796 14272 34848 14278
rect 34796 14214 34848 14220
rect 34612 14000 34664 14006
rect 34612 13942 34664 13948
rect 34808 13938 34836 14214
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 35072 13932 35124 13938
rect 35072 13874 35124 13880
rect 35084 13818 35112 13874
rect 34808 13790 35112 13818
rect 34244 13728 34296 13734
rect 34244 13670 34296 13676
rect 34256 12918 34284 13670
rect 34808 13462 34836 13790
rect 35176 13734 35204 14282
rect 35164 13728 35216 13734
rect 35164 13670 35216 13676
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 13456 34848 13462
rect 34796 13398 34848 13404
rect 34888 13456 34940 13462
rect 34888 13398 34940 13404
rect 34704 13252 34756 13258
rect 34704 13194 34756 13200
rect 34244 12912 34296 12918
rect 34244 12854 34296 12860
rect 34256 12782 34284 12854
rect 34336 12844 34388 12850
rect 34336 12786 34388 12792
rect 34244 12776 34296 12782
rect 34244 12718 34296 12724
rect 34348 12434 34376 12786
rect 34256 12406 34376 12434
rect 34256 12238 34284 12406
rect 34520 12368 34572 12374
rect 34520 12310 34572 12316
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 34256 11762 34284 12174
rect 34336 12164 34388 12170
rect 34336 12106 34388 12112
rect 34348 11898 34376 12106
rect 34336 11892 34388 11898
rect 34336 11834 34388 11840
rect 34532 11830 34560 12310
rect 34612 12096 34664 12102
rect 34612 12038 34664 12044
rect 34520 11824 34572 11830
rect 34520 11766 34572 11772
rect 34244 11756 34296 11762
rect 34244 11698 34296 11704
rect 34152 11552 34204 11558
rect 34152 11494 34204 11500
rect 34164 10674 34192 11494
rect 34152 10668 34204 10674
rect 34152 10610 34204 10616
rect 34060 9580 34112 9586
rect 34060 9522 34112 9528
rect 33692 9172 33744 9178
rect 33692 9114 33744 9120
rect 33704 8974 33732 9114
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 33968 8968 34020 8974
rect 33968 8910 34020 8916
rect 32772 8900 32824 8906
rect 32772 8842 32824 8848
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 32588 8832 32640 8838
rect 32588 8774 32640 8780
rect 32600 8650 32628 8774
rect 32508 8622 32628 8650
rect 32508 8498 32536 8622
rect 32784 8566 32812 8842
rect 32772 8560 32824 8566
rect 32772 8502 32824 8508
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32508 7818 32536 8434
rect 33704 8090 33732 8910
rect 33980 8634 34008 8910
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 33968 8356 34020 8362
rect 33968 8298 34020 8304
rect 33692 8084 33744 8090
rect 33692 8026 33744 8032
rect 32772 7948 32824 7954
rect 32772 7890 32824 7896
rect 32496 7812 32548 7818
rect 32496 7754 32548 7760
rect 32404 7472 32456 7478
rect 32404 7414 32456 7420
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 31852 6656 31904 6662
rect 31852 6598 31904 6604
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 31668 6112 31720 6118
rect 31668 6054 31720 6060
rect 31680 5574 31708 6054
rect 31864 5710 31892 6598
rect 32324 6458 32352 7142
rect 32416 7002 32444 7414
rect 32404 6996 32456 7002
rect 32404 6938 32456 6944
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32784 6390 32812 7890
rect 33232 7744 33284 7750
rect 33232 7686 33284 7692
rect 32956 6724 33008 6730
rect 32956 6666 33008 6672
rect 32968 6458 32996 6666
rect 32956 6452 33008 6458
rect 32956 6394 33008 6400
rect 33244 6390 33272 7686
rect 33508 7200 33560 7206
rect 33508 7142 33560 7148
rect 32772 6384 32824 6390
rect 32678 6352 32734 6361
rect 32772 6326 32824 6332
rect 33232 6384 33284 6390
rect 33232 6326 33284 6332
rect 32678 6287 32680 6296
rect 32732 6287 32734 6296
rect 32680 6258 32732 6264
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 31668 5568 31720 5574
rect 31668 5510 31720 5516
rect 32692 5302 32720 6258
rect 32784 6118 32812 6326
rect 33140 6180 33192 6186
rect 33140 6122 33192 6128
rect 32772 6112 32824 6118
rect 32772 6054 32824 6060
rect 33152 5710 33180 6122
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 32680 5296 32732 5302
rect 32680 5238 32732 5244
rect 31576 5228 31628 5234
rect 31576 5170 31628 5176
rect 31588 4622 31616 5170
rect 33244 4826 33272 6326
rect 33520 6322 33548 7142
rect 33508 6316 33560 6322
rect 33508 6258 33560 6264
rect 33520 5302 33548 6258
rect 33980 5302 34008 8298
rect 34072 6186 34100 9522
rect 34164 8498 34192 10610
rect 34256 8974 34284 11698
rect 34428 11620 34480 11626
rect 34428 11562 34480 11568
rect 34440 11393 34468 11562
rect 34426 11384 34482 11393
rect 34426 11319 34482 11328
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34336 10736 34388 10742
rect 34336 10678 34388 10684
rect 34244 8968 34296 8974
rect 34244 8910 34296 8916
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34164 7410 34192 8434
rect 34152 7404 34204 7410
rect 34152 7346 34204 7352
rect 34060 6180 34112 6186
rect 34060 6122 34112 6128
rect 34256 5710 34284 8910
rect 34348 8634 34376 10678
rect 34440 10470 34468 11086
rect 34624 10742 34652 12038
rect 34716 11150 34744 13194
rect 34900 12628 34928 13398
rect 34808 12600 34928 12628
rect 34808 12434 34836 12600
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12442 35388 15030
rect 35440 14340 35492 14346
rect 35440 14282 35492 14288
rect 35452 14074 35480 14282
rect 35440 14068 35492 14074
rect 35440 14010 35492 14016
rect 35544 13938 35572 19382
rect 36096 18834 36124 19790
rect 36188 19786 36216 20567
rect 37096 19848 37148 19854
rect 37096 19790 37148 19796
rect 36176 19780 36228 19786
rect 36176 19722 36228 19728
rect 36084 18828 36136 18834
rect 36084 18770 36136 18776
rect 36096 18358 36124 18770
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 36096 17882 36124 18294
rect 36084 17876 36136 17882
rect 36084 17818 36136 17824
rect 36188 17762 36216 19722
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36556 19378 36584 19654
rect 37108 19378 37136 19790
rect 37200 19718 37228 20878
rect 37384 20058 37412 20878
rect 37372 20052 37424 20058
rect 37372 19994 37424 20000
rect 37476 19922 37504 21490
rect 37752 21146 37780 21490
rect 37740 21140 37792 21146
rect 37740 21082 37792 21088
rect 37556 20936 37608 20942
rect 37556 20878 37608 20884
rect 37568 20262 37596 20878
rect 37648 20868 37700 20874
rect 37648 20810 37700 20816
rect 37556 20256 37608 20262
rect 37556 20198 37608 20204
rect 37464 19916 37516 19922
rect 37464 19858 37516 19864
rect 37372 19848 37424 19854
rect 37372 19790 37424 19796
rect 37188 19712 37240 19718
rect 37188 19654 37240 19660
rect 37280 19508 37332 19514
rect 37280 19450 37332 19456
rect 36544 19372 36596 19378
rect 36544 19314 36596 19320
rect 37096 19372 37148 19378
rect 37096 19314 37148 19320
rect 36268 19236 36320 19242
rect 36268 19178 36320 19184
rect 36452 19236 36504 19242
rect 36452 19178 36504 19184
rect 36280 18970 36308 19178
rect 36268 18964 36320 18970
rect 36268 18906 36320 18912
rect 36268 18624 36320 18630
rect 36268 18566 36320 18572
rect 36280 18290 36308 18566
rect 36464 18426 36492 19178
rect 37292 18766 37320 19450
rect 37384 19378 37412 19790
rect 37372 19372 37424 19378
rect 37372 19314 37424 19320
rect 37280 18760 37332 18766
rect 37280 18702 37332 18708
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 36452 18420 36504 18426
rect 36452 18362 36504 18368
rect 36268 18284 36320 18290
rect 36268 18226 36320 18232
rect 36096 17734 36216 17762
rect 35992 17604 36044 17610
rect 35992 17546 36044 17552
rect 35808 17536 35860 17542
rect 35808 17478 35860 17484
rect 35716 17264 35768 17270
rect 35716 17206 35768 17212
rect 35728 16046 35756 17206
rect 35820 16726 35848 17478
rect 35808 16720 35860 16726
rect 35808 16662 35860 16668
rect 35900 16652 35952 16658
rect 35900 16594 35952 16600
rect 35716 16040 35768 16046
rect 35716 15982 35768 15988
rect 35728 15434 35756 15982
rect 35716 15428 35768 15434
rect 35716 15370 35768 15376
rect 35912 14822 35940 16594
rect 36004 16114 36032 17546
rect 35992 16108 36044 16114
rect 35992 16050 36044 16056
rect 36004 15638 36032 16050
rect 35992 15632 36044 15638
rect 35992 15574 36044 15580
rect 35900 14816 35952 14822
rect 35900 14758 35952 14764
rect 35808 14408 35860 14414
rect 35808 14350 35860 14356
rect 35532 13932 35584 13938
rect 35532 13874 35584 13880
rect 35532 13728 35584 13734
rect 35532 13670 35584 13676
rect 35544 13258 35572 13670
rect 35820 13530 35848 14350
rect 35900 13864 35952 13870
rect 35900 13806 35952 13812
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35716 13320 35768 13326
rect 35716 13262 35768 13268
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35440 12844 35492 12850
rect 35440 12786 35492 12792
rect 35348 12436 35400 12442
rect 34808 12406 35112 12434
rect 35084 11762 35112 12406
rect 35348 12378 35400 12384
rect 35072 11756 35124 11762
rect 35072 11698 35124 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 34612 10736 34664 10742
rect 34612 10678 34664 10684
rect 34428 10464 34480 10470
rect 34428 10406 34480 10412
rect 34440 9994 34468 10406
rect 34428 9988 34480 9994
rect 34428 9930 34480 9936
rect 34336 8628 34388 8634
rect 34336 8570 34388 8576
rect 34440 7886 34468 9930
rect 34624 8838 34652 10678
rect 34716 10674 34744 11086
rect 34704 10668 34756 10674
rect 34704 10610 34756 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34888 9988 34940 9994
rect 34888 9930 34940 9936
rect 34796 9920 34848 9926
rect 34796 9862 34848 9868
rect 34808 9654 34836 9862
rect 34796 9648 34848 9654
rect 34796 9590 34848 9596
rect 34704 9580 34756 9586
rect 34704 9522 34756 9528
rect 34716 9178 34744 9522
rect 34900 9466 34928 9930
rect 34808 9438 34928 9466
rect 34808 9382 34836 9438
rect 34796 9376 34848 9382
rect 34796 9318 34848 9324
rect 34704 9172 34756 9178
rect 34704 9114 34756 9120
rect 34808 9042 34836 9318
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 9036 34848 9042
rect 34796 8978 34848 8984
rect 34612 8832 34664 8838
rect 34612 8774 34664 8780
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34532 7478 34560 8026
rect 34520 7472 34572 7478
rect 34520 7414 34572 7420
rect 34624 7410 34652 8774
rect 35268 8566 35296 8774
rect 35256 8560 35308 8566
rect 35256 8502 35308 8508
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34612 7404 34664 7410
rect 34612 7346 34664 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34244 5704 34296 5710
rect 34244 5646 34296 5652
rect 34072 5302 34100 5646
rect 33508 5296 33560 5302
rect 33508 5238 33560 5244
rect 33968 5296 34020 5302
rect 33968 5238 34020 5244
rect 34060 5296 34112 5302
rect 34060 5238 34112 5244
rect 33232 4820 33284 4826
rect 33232 4762 33284 4768
rect 31576 4616 31628 4622
rect 31576 4558 31628 4564
rect 31484 4208 31536 4214
rect 31484 4150 31536 4156
rect 31588 4146 31616 4558
rect 33980 4282 34008 5238
rect 34256 5234 34284 5646
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34244 5228 34296 5234
rect 34244 5170 34296 5176
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 34072 4486 34100 5102
rect 34060 4480 34112 4486
rect 34060 4422 34112 4428
rect 33968 4276 34020 4282
rect 33968 4218 34020 4224
rect 34532 4146 34560 5510
rect 34624 5302 34652 6054
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35360 5642 35388 12378
rect 35452 11898 35480 12786
rect 35728 12374 35756 13262
rect 35716 12368 35768 12374
rect 35716 12310 35768 12316
rect 35912 12238 35940 13806
rect 36096 13297 36124 17734
rect 36176 16992 36228 16998
rect 36176 16934 36228 16940
rect 36188 16590 36216 16934
rect 36176 16584 36228 16590
rect 36280 16561 36308 18226
rect 36728 17604 36780 17610
rect 36728 17546 36780 17552
rect 36740 17202 36768 17546
rect 36544 17196 36596 17202
rect 36544 17138 36596 17144
rect 36728 17196 36780 17202
rect 36728 17138 36780 17144
rect 36556 16794 36584 17138
rect 36544 16788 36596 16794
rect 36544 16730 36596 16736
rect 36176 16526 36228 16532
rect 36266 16552 36322 16561
rect 36266 16487 36322 16496
rect 36544 16516 36596 16522
rect 36544 16458 36596 16464
rect 36556 16250 36584 16458
rect 36544 16244 36596 16250
rect 36544 16186 36596 16192
rect 36176 15360 36228 15366
rect 36176 15302 36228 15308
rect 36188 15162 36216 15302
rect 36176 15156 36228 15162
rect 36176 15098 36228 15104
rect 37096 14408 37148 14414
rect 37096 14350 37148 14356
rect 36452 14272 36504 14278
rect 36452 14214 36504 14220
rect 36464 14006 36492 14214
rect 36452 14000 36504 14006
rect 36452 13942 36504 13948
rect 36176 13932 36228 13938
rect 36176 13874 36228 13880
rect 36360 13932 36412 13938
rect 36360 13874 36412 13880
rect 36188 13462 36216 13874
rect 36176 13456 36228 13462
rect 36176 13398 36228 13404
rect 36372 13394 36400 13874
rect 36360 13388 36412 13394
rect 36360 13330 36412 13336
rect 36082 13288 36138 13297
rect 36082 13223 36138 13232
rect 35900 12232 35952 12238
rect 35900 12174 35952 12180
rect 35440 11892 35492 11898
rect 35440 11834 35492 11840
rect 35716 11824 35768 11830
rect 35716 11766 35768 11772
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 35452 11354 35480 11630
rect 35440 11348 35492 11354
rect 35440 11290 35492 11296
rect 35728 11014 35756 11766
rect 36360 11756 36412 11762
rect 36360 11698 36412 11704
rect 35716 11008 35768 11014
rect 35716 10950 35768 10956
rect 35728 10266 35756 10950
rect 36372 10742 36400 11698
rect 36464 11694 36492 13942
rect 37108 12850 37136 14350
rect 37096 12844 37148 12850
rect 37096 12786 37148 12792
rect 37108 12238 37136 12786
rect 37096 12232 37148 12238
rect 37096 12174 37148 12180
rect 37108 11830 37136 12174
rect 37096 11824 37148 11830
rect 37096 11766 37148 11772
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36360 10736 36412 10742
rect 36360 10678 36412 10684
rect 36372 10470 36400 10678
rect 36464 10606 36492 11630
rect 36820 11552 36872 11558
rect 36820 11494 36872 11500
rect 36832 11082 36860 11494
rect 37108 11150 37136 11766
rect 37292 11762 37320 18566
rect 37384 12714 37412 19314
rect 37476 18766 37504 19858
rect 37556 19372 37608 19378
rect 37556 19314 37608 19320
rect 37568 19174 37596 19314
rect 37556 19168 37608 19174
rect 37556 19110 37608 19116
rect 37464 18760 37516 18766
rect 37464 18702 37516 18708
rect 37476 18290 37504 18702
rect 37568 18630 37596 19110
rect 37660 18970 37688 20810
rect 38672 20806 38700 22374
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 39304 21616 39356 21622
rect 39304 21558 39356 21564
rect 38844 21344 38896 21350
rect 38844 21286 38896 21292
rect 38660 20800 38712 20806
rect 38660 20742 38712 20748
rect 38856 20641 38884 21286
rect 38842 20632 38898 20641
rect 38842 20567 38898 20576
rect 38108 19780 38160 19786
rect 38108 19722 38160 19728
rect 38120 19514 38148 19722
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 38108 19508 38160 19514
rect 38108 19450 38160 19456
rect 38856 19378 38884 19654
rect 38476 19372 38528 19378
rect 38476 19314 38528 19320
rect 38844 19372 38896 19378
rect 38844 19314 38896 19320
rect 38488 18970 38516 19314
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 38476 18964 38528 18970
rect 38476 18906 38528 18912
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 38016 18284 38068 18290
rect 38016 18226 38068 18232
rect 38028 17882 38056 18226
rect 38752 18080 38804 18086
rect 38752 18022 38804 18028
rect 38016 17876 38068 17882
rect 38016 17818 38068 17824
rect 38660 17672 38712 17678
rect 38660 17614 38712 17620
rect 37740 17604 37792 17610
rect 37740 17546 37792 17552
rect 37752 17270 37780 17546
rect 38672 17338 38700 17614
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 37740 17264 37792 17270
rect 38764 17218 38792 18022
rect 38856 17678 38884 19314
rect 38844 17672 38896 17678
rect 38844 17614 38896 17620
rect 37740 17206 37792 17212
rect 38672 17202 38792 17218
rect 38476 17196 38528 17202
rect 38476 17138 38528 17144
rect 38660 17196 38792 17202
rect 38712 17190 38792 17196
rect 38660 17138 38712 17144
rect 37648 16584 37700 16590
rect 37648 16526 37700 16532
rect 37464 16448 37516 16454
rect 37464 16390 37516 16396
rect 37476 16114 37504 16390
rect 37660 16182 37688 16526
rect 38488 16182 38516 17138
rect 37648 16176 37700 16182
rect 37648 16118 37700 16124
rect 38476 16176 38528 16182
rect 38476 16118 38528 16124
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37476 12986 37504 16050
rect 37556 15360 37608 15366
rect 37556 15302 37608 15308
rect 37568 15094 37596 15302
rect 37556 15088 37608 15094
rect 37556 15030 37608 15036
rect 37660 15026 37688 16118
rect 38672 15706 38700 17138
rect 39120 16584 39172 16590
rect 39120 16526 39172 16532
rect 38660 15700 38712 15706
rect 38660 15642 38712 15648
rect 39132 15570 39160 16526
rect 39120 15564 39172 15570
rect 39120 15506 39172 15512
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 38844 14408 38896 14414
rect 38842 14376 38844 14385
rect 39028 14408 39080 14414
rect 38896 14376 38898 14385
rect 39132 14396 39160 15506
rect 39316 15162 39344 21558
rect 67640 21344 67692 21350
rect 67640 21286 67692 21292
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 67652 21185 67680 21286
rect 67638 21176 67694 21185
rect 67638 21111 67694 21120
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 40408 20256 40460 20262
rect 40408 20198 40460 20204
rect 39304 15156 39356 15162
rect 39304 15098 39356 15104
rect 40224 15156 40276 15162
rect 40224 15098 40276 15104
rect 39080 14368 39160 14396
rect 39028 14350 39080 14356
rect 38842 14311 38898 14320
rect 39132 13394 39160 14368
rect 39316 14074 39344 15098
rect 39948 14612 40000 14618
rect 39948 14554 40000 14560
rect 39396 14408 39448 14414
rect 39396 14350 39448 14356
rect 39304 14068 39356 14074
rect 39304 14010 39356 14016
rect 39120 13388 39172 13394
rect 39120 13330 39172 13336
rect 37464 12980 37516 12986
rect 37464 12922 37516 12928
rect 37372 12708 37424 12714
rect 37372 12650 37424 12656
rect 38844 12708 38896 12714
rect 38844 12650 38896 12656
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37476 12442 37504 12582
rect 37464 12436 37516 12442
rect 38856 12434 38884 12650
rect 39132 12442 39160 13330
rect 39316 13326 39344 14010
rect 39408 13938 39436 14350
rect 39764 14340 39816 14346
rect 39764 14282 39816 14288
rect 39776 14074 39804 14282
rect 39764 14068 39816 14074
rect 39764 14010 39816 14016
rect 39960 14006 39988 14554
rect 40236 14414 40264 15098
rect 40224 14408 40276 14414
rect 40224 14350 40276 14356
rect 40316 14272 40368 14278
rect 40316 14214 40368 14220
rect 39948 14000 40000 14006
rect 39948 13942 40000 13948
rect 39396 13932 39448 13938
rect 39396 13874 39448 13880
rect 39764 13932 39816 13938
rect 39764 13874 39816 13880
rect 39304 13320 39356 13326
rect 39304 13262 39356 13268
rect 39120 12436 39172 12442
rect 38856 12406 39068 12434
rect 37464 12378 37516 12384
rect 37476 12238 37504 12378
rect 39040 12238 39068 12406
rect 39120 12378 39172 12384
rect 37464 12232 37516 12238
rect 37464 12174 37516 12180
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 39040 11898 39068 12174
rect 39028 11892 39080 11898
rect 39028 11834 39080 11840
rect 37280 11756 37332 11762
rect 37280 11698 37332 11704
rect 38936 11348 38988 11354
rect 38936 11290 38988 11296
rect 37556 11280 37608 11286
rect 37554 11248 37556 11257
rect 37608 11248 37610 11257
rect 37554 11183 37610 11192
rect 37096 11144 37148 11150
rect 37096 11086 37148 11092
rect 36728 11076 36780 11082
rect 36728 11018 36780 11024
rect 36820 11076 36872 11082
rect 36820 11018 36872 11024
rect 36452 10600 36504 10606
rect 36452 10542 36504 10548
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 35716 10260 35768 10266
rect 35716 10202 35768 10208
rect 35624 9988 35676 9994
rect 35624 9930 35676 9936
rect 35636 9518 35664 9930
rect 36740 9518 36768 11018
rect 37568 10742 37596 11183
rect 38844 11144 38896 11150
rect 38844 11086 38896 11092
rect 38660 10804 38712 10810
rect 38660 10746 38712 10752
rect 37556 10736 37608 10742
rect 37556 10678 37608 10684
rect 38292 10192 38344 10198
rect 38292 10134 38344 10140
rect 37556 10056 37608 10062
rect 37556 9998 37608 10004
rect 37568 9722 37596 9998
rect 37556 9716 37608 9722
rect 37556 9658 37608 9664
rect 35624 9512 35676 9518
rect 35624 9454 35676 9460
rect 36728 9512 36780 9518
rect 36728 9454 36780 9460
rect 35532 8492 35584 8498
rect 35532 8434 35584 8440
rect 35544 8090 35572 8434
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35544 6866 35572 8026
rect 35636 7954 35664 9454
rect 36360 9376 36412 9382
rect 36360 9318 36412 9324
rect 36372 8566 36400 9318
rect 36740 9042 36768 9454
rect 36728 9036 36780 9042
rect 36728 8978 36780 8984
rect 36360 8560 36412 8566
rect 36360 8502 36412 8508
rect 36268 8288 36320 8294
rect 36268 8230 36320 8236
rect 35624 7948 35676 7954
rect 35624 7890 35676 7896
rect 36280 7886 36308 8230
rect 36372 8022 36400 8502
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37292 8090 37320 8434
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 36360 8016 36412 8022
rect 36360 7958 36412 7964
rect 35900 7880 35952 7886
rect 35900 7822 35952 7828
rect 36268 7880 36320 7886
rect 36268 7822 36320 7828
rect 35912 7410 35940 7822
rect 36176 7744 36228 7750
rect 36176 7686 36228 7692
rect 35900 7404 35952 7410
rect 36084 7404 36136 7410
rect 35900 7346 35952 7352
rect 36004 7364 36084 7392
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35532 6860 35584 6866
rect 35532 6802 35584 6808
rect 35636 6322 35664 7142
rect 36004 6866 36032 7364
rect 36084 7346 36136 7352
rect 36084 7268 36136 7274
rect 36188 7256 36216 7686
rect 36372 7546 36400 7958
rect 36268 7540 36320 7546
rect 36268 7482 36320 7488
rect 36360 7540 36412 7546
rect 36360 7482 36412 7488
rect 36136 7228 36216 7256
rect 36084 7210 36136 7216
rect 36280 6934 36308 7482
rect 36544 7200 36596 7206
rect 36544 7142 36596 7148
rect 36268 6928 36320 6934
rect 36268 6870 36320 6876
rect 35992 6860 36044 6866
rect 35992 6802 36044 6808
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 35532 6112 35584 6118
rect 35532 6054 35584 6060
rect 35072 5636 35124 5642
rect 35072 5578 35124 5584
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 35084 5370 35112 5578
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 35072 5364 35124 5370
rect 35072 5306 35124 5312
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34808 4826 34836 5306
rect 35348 5024 35400 5030
rect 35348 4966 35400 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34796 4820 34848 4826
rect 34796 4762 34848 4768
rect 35164 4616 35216 4622
rect 35164 4558 35216 4564
rect 35176 4146 35204 4558
rect 35360 4554 35388 4966
rect 35544 4622 35572 6054
rect 35636 5778 35664 6258
rect 35624 5772 35676 5778
rect 35624 5714 35676 5720
rect 35636 5302 35664 5714
rect 35624 5296 35676 5302
rect 35624 5238 35676 5244
rect 35636 5166 35664 5238
rect 36004 5234 36032 6258
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 36280 5216 36308 6870
rect 36556 6730 36584 7142
rect 36544 6724 36596 6730
rect 36544 6666 36596 6672
rect 37280 6724 37332 6730
rect 37280 6666 37332 6672
rect 37188 6248 37240 6254
rect 37188 6190 37240 6196
rect 37200 5370 37228 6190
rect 37292 5642 37320 6666
rect 37280 5636 37332 5642
rect 37280 5578 37332 5584
rect 37188 5364 37240 5370
rect 37188 5306 37240 5312
rect 36360 5228 36412 5234
rect 36280 5188 36360 5216
rect 35624 5160 35676 5166
rect 35624 5102 35676 5108
rect 35532 4616 35584 4622
rect 35532 4558 35584 4564
rect 35348 4548 35400 4554
rect 35348 4490 35400 4496
rect 36280 4282 36308 5188
rect 36360 5170 36412 5176
rect 36820 5228 36872 5234
rect 36820 5170 36872 5176
rect 36636 5024 36688 5030
rect 36636 4966 36688 4972
rect 36648 4690 36676 4966
rect 36636 4684 36688 4690
rect 36636 4626 36688 4632
rect 36832 4486 36860 5170
rect 37292 4622 37320 5578
rect 38304 5302 38332 10134
rect 38384 7200 38436 7206
rect 38384 7142 38436 7148
rect 38396 5710 38424 7142
rect 38672 6798 38700 10746
rect 38856 9586 38884 11086
rect 38948 10674 38976 11290
rect 38936 10668 38988 10674
rect 38936 10610 38988 10616
rect 38948 9994 38976 10610
rect 38936 9988 38988 9994
rect 38936 9930 38988 9936
rect 38844 9580 38896 9586
rect 38844 9522 38896 9528
rect 38856 8498 38884 9522
rect 38844 8492 38896 8498
rect 38844 8434 38896 8440
rect 39040 7410 39068 11834
rect 39132 11762 39160 12378
rect 39776 11830 39804 13874
rect 40132 13456 40184 13462
rect 40132 13398 40184 13404
rect 39948 13252 40000 13258
rect 39948 13194 40000 13200
rect 39764 11824 39816 11830
rect 39764 11766 39816 11772
rect 39120 11756 39172 11762
rect 39120 11698 39172 11704
rect 39132 11218 39160 11698
rect 39120 11212 39172 11218
rect 39120 11154 39172 11160
rect 39960 10674 39988 13194
rect 40144 11234 40172 13398
rect 40328 12102 40356 14214
rect 40420 12238 40448 20198
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 68100 19848 68152 19854
rect 68098 19816 68100 19825
rect 68152 19816 68154 19825
rect 68098 19751 68154 19760
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 68100 18760 68152 18766
rect 68100 18702 68152 18708
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 68112 18465 68140 18702
rect 68098 18456 68154 18465
rect 68098 18391 68154 18400
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 67638 17096 67694 17105
rect 67638 17031 67640 17040
rect 67692 17031 67694 17040
rect 67640 17002 67692 17008
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 67640 15904 67692 15910
rect 67640 15846 67692 15852
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 67652 15745 67680 15846
rect 67638 15736 67694 15745
rect 67638 15671 67694 15680
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 68100 14408 68152 14414
rect 40498 14376 40554 14385
rect 40498 14311 40500 14320
rect 40552 14311 40554 14320
rect 68098 14376 68100 14385
rect 68152 14376 68154 14385
rect 68098 14311 68154 14320
rect 40500 14282 40552 14288
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 40500 13320 40552 13326
rect 40500 13262 40552 13268
rect 68100 13320 68152 13326
rect 68100 13262 68152 13268
rect 40512 12850 40540 13262
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 68112 13025 68140 13262
rect 68098 13016 68154 13025
rect 68098 12951 68154 12960
rect 40500 12844 40552 12850
rect 40500 12786 40552 12792
rect 40408 12232 40460 12238
rect 40408 12174 40460 12180
rect 40224 12096 40276 12102
rect 40224 12038 40276 12044
rect 40316 12096 40368 12102
rect 40316 12038 40368 12044
rect 40236 11898 40264 12038
rect 40224 11892 40276 11898
rect 40224 11834 40276 11840
rect 40144 11206 40264 11234
rect 40420 11218 40448 12174
rect 40132 11144 40184 11150
rect 40132 11086 40184 11092
rect 40144 10742 40172 11086
rect 40236 11014 40264 11206
rect 40408 11212 40460 11218
rect 40408 11154 40460 11160
rect 40512 11150 40540 12786
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 40684 12164 40736 12170
rect 40684 12106 40736 12112
rect 40696 11830 40724 12106
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 40684 11824 40736 11830
rect 40684 11766 40736 11772
rect 67638 11656 67694 11665
rect 67638 11591 67640 11600
rect 67692 11591 67694 11600
rect 67640 11562 67692 11568
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 40316 11144 40368 11150
rect 40316 11086 40368 11092
rect 40500 11144 40552 11150
rect 40500 11086 40552 11092
rect 40224 11008 40276 11014
rect 40224 10950 40276 10956
rect 40132 10736 40184 10742
rect 40132 10678 40184 10684
rect 39948 10668 40000 10674
rect 39948 10610 40000 10616
rect 39764 10464 39816 10470
rect 39764 10406 39816 10412
rect 39776 10062 39804 10406
rect 40236 10198 40264 10950
rect 40328 10810 40356 11086
rect 40316 10804 40368 10810
rect 40316 10746 40368 10752
rect 40224 10192 40276 10198
rect 40224 10134 40276 10140
rect 40512 10062 40540 11086
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 67640 10464 67692 10470
rect 67640 10406 67692 10412
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 67652 10305 67680 10406
rect 67638 10296 67694 10305
rect 67638 10231 67694 10240
rect 39764 10056 39816 10062
rect 39764 9998 39816 10004
rect 40500 10056 40552 10062
rect 40500 9998 40552 10004
rect 39776 9722 39804 9998
rect 39856 9920 39908 9926
rect 39856 9862 39908 9868
rect 39764 9716 39816 9722
rect 39764 9658 39816 9664
rect 39868 9654 39896 9862
rect 39856 9648 39908 9654
rect 39856 9590 39908 9596
rect 40512 8022 40540 9998
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 68100 8968 68152 8974
rect 68098 8936 68100 8945
rect 68152 8936 68154 8945
rect 68098 8871 68154 8880
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 40500 8016 40552 8022
rect 40500 7958 40552 7964
rect 68100 7880 68152 7886
rect 68100 7822 68152 7828
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 68112 7585 68140 7822
rect 68098 7576 68154 7585
rect 68098 7511 68154 7520
rect 38844 7404 38896 7410
rect 38844 7346 38896 7352
rect 39028 7404 39080 7410
rect 39028 7346 39080 7352
rect 38856 7002 38884 7346
rect 38844 6996 38896 7002
rect 38844 6938 38896 6944
rect 38660 6792 38712 6798
rect 38660 6734 38712 6740
rect 38672 5914 38700 6734
rect 38752 6724 38804 6730
rect 38752 6666 38804 6672
rect 38660 5908 38712 5914
rect 38660 5850 38712 5856
rect 38384 5704 38436 5710
rect 38384 5646 38436 5652
rect 38292 5296 38344 5302
rect 38292 5238 38344 5244
rect 38304 4826 38332 5238
rect 38764 5234 38792 6666
rect 39040 6322 39068 7346
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 39028 6316 39080 6322
rect 39028 6258 39080 6264
rect 67638 6216 67694 6225
rect 67638 6151 67640 6160
rect 67692 6151 67694 6160
rect 67640 6122 67692 6128
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 38752 5228 38804 5234
rect 38752 5170 38804 5176
rect 58808 5160 58860 5166
rect 58808 5102 58860 5108
rect 58716 5024 58768 5030
rect 58716 4966 58768 4972
rect 38292 4820 38344 4826
rect 38292 4762 38344 4768
rect 57244 4752 57296 4758
rect 57244 4694 57296 4700
rect 58256 4752 58308 4758
rect 58256 4694 58308 4700
rect 37280 4616 37332 4622
rect 37280 4558 37332 4564
rect 57152 4616 57204 4622
rect 57152 4558 57204 4564
rect 36820 4480 36872 4486
rect 36820 4422 36872 4428
rect 36268 4276 36320 4282
rect 36268 4218 36320 4224
rect 36832 4214 36860 4422
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 36820 4208 36872 4214
rect 36820 4150 36872 4156
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 34520 4140 34572 4146
rect 34520 4082 34572 4088
rect 35164 4140 35216 4146
rect 35164 4082 35216 4088
rect 28736 3534 28764 4082
rect 29012 3738 29040 4082
rect 56140 3936 56192 3942
rect 56140 3878 56192 3884
rect 56324 3936 56376 3942
rect 56324 3878 56376 3884
rect 56968 3936 57020 3942
rect 56968 3878 57020 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 41144 3664 41196 3670
rect 41144 3606 41196 3612
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 29828 3528 29880 3534
rect 29828 3470 29880 3476
rect 30656 3528 30708 3534
rect 30656 3470 30708 3476
rect 31484 3528 31536 3534
rect 31484 3470 31536 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24676 2032 24728 2038
rect 24676 1974 24728 1980
rect 24872 800 24900 2790
rect 25148 800 25176 3470
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25424 800 25452 2382
rect 25700 800 25728 2790
rect 25976 800 26004 3470
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26252 800 26280 2790
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26528 800 26556 2450
rect 26804 800 26832 3470
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 27080 800 27108 2790
rect 27344 2576 27396 2582
rect 27344 2518 27396 2524
rect 27356 800 27384 2518
rect 27632 800 27660 3470
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 28724 2848 28776 2854
rect 28724 2790 28776 2796
rect 29276 2848 29328 2854
rect 29276 2790 29328 2796
rect 27896 2372 27948 2378
rect 27896 2314 27948 2320
rect 27908 800 27936 2314
rect 28184 800 28212 2790
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 28460 800 28488 2382
rect 28736 800 28764 2790
rect 29000 2576 29052 2582
rect 29000 2518 29052 2524
rect 29012 800 29040 2518
rect 29288 800 29316 2790
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29564 800 29592 2382
rect 29840 800 29868 3470
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30116 800 30144 2790
rect 30392 800 30420 2790
rect 30668 800 30696 3470
rect 31208 2848 31260 2854
rect 31208 2790 31260 2796
rect 30932 2576 30984 2582
rect 30932 2518 30984 2524
rect 30944 800 30972 2518
rect 31220 800 31248 2790
rect 31496 800 31524 3470
rect 32036 2848 32088 2854
rect 32036 2790 32088 2796
rect 31760 2372 31812 2378
rect 31760 2314 31812 2320
rect 31772 800 31800 2314
rect 32048 800 32076 2790
rect 32324 800 32352 3470
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32588 2440 32640 2446
rect 32588 2382 32640 2388
rect 32600 800 32628 2382
rect 32876 800 32904 2790
rect 33152 800 33180 3470
rect 37280 2984 37332 2990
rect 37280 2926 37332 2932
rect 33692 2848 33744 2854
rect 33692 2790 33744 2796
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33428 800 33456 2382
rect 33704 800 33732 2790
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 33980 800 34008 2382
rect 34256 800 34284 2790
rect 34532 800 34560 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35072 2440 35124 2446
rect 35072 2382 35124 2388
rect 34808 800 34836 2382
rect 35084 800 35112 2382
rect 35360 800 35388 2790
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35636 800 35664 2382
rect 35912 800 35940 2382
rect 36188 800 36216 2790
rect 36452 2440 36504 2446
rect 36452 2382 36504 2388
rect 36464 800 36492 2382
rect 36740 800 36768 2790
rect 37004 2508 37056 2514
rect 37004 2450 37056 2456
rect 37016 800 37044 2450
rect 37292 800 37320 2926
rect 38384 2916 38436 2922
rect 38384 2858 38436 2864
rect 37832 2848 37884 2854
rect 37832 2790 37884 2796
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 37568 800 37596 2382
rect 37844 800 37872 2790
rect 38108 2508 38160 2514
rect 38108 2450 38160 2456
rect 38120 800 38148 2450
rect 38396 800 38424 2858
rect 38936 2848 38988 2854
rect 38936 2790 38988 2796
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38672 800 38700 2382
rect 38948 800 38976 2790
rect 39224 800 39252 3470
rect 39764 2916 39816 2922
rect 39764 2858 39816 2864
rect 39488 2372 39540 2378
rect 39488 2314 39540 2320
rect 39500 800 39528 2314
rect 39776 800 39804 2858
rect 40052 800 40080 3470
rect 40316 2848 40368 2854
rect 40316 2790 40368 2796
rect 40328 800 40356 2790
rect 40592 2576 40644 2582
rect 40592 2518 40644 2524
rect 40604 800 40632 2518
rect 40880 800 40908 3470
rect 41156 800 41184 3606
rect 55772 3596 55824 3602
rect 55772 3538 55824 3544
rect 42524 3528 42576 3534
rect 42524 3470 42576 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 45008 3528 45060 3534
rect 45008 3470 45060 3476
rect 45284 3528 45336 3534
rect 45284 3470 45336 3476
rect 46112 3528 46164 3534
rect 46112 3470 46164 3476
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 47768 3528 47820 3534
rect 47768 3470 47820 3476
rect 48872 3528 48924 3534
rect 48872 3470 48924 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50804 3528 50856 3534
rect 50804 3470 50856 3476
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 52736 3528 52788 3534
rect 52736 3470 52788 3476
rect 53012 3528 53064 3534
rect 53012 3470 53064 3476
rect 54668 3528 54720 3534
rect 54668 3470 54720 3476
rect 55496 3528 55548 3534
rect 55496 3470 55548 3476
rect 42248 2916 42300 2922
rect 42248 2858 42300 2864
rect 41696 2848 41748 2854
rect 41696 2790 41748 2796
rect 41420 2508 41472 2514
rect 41420 2450 41472 2456
rect 41432 800 41460 2450
rect 41708 800 41736 2790
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 41984 800 42012 2382
rect 42260 800 42288 2858
rect 42536 800 42564 3470
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42812 800 42840 2790
rect 43088 800 43116 3470
rect 44732 2984 44784 2990
rect 44732 2926 44784 2932
rect 43628 2916 43680 2922
rect 43628 2858 43680 2864
rect 43352 2508 43404 2514
rect 43352 2450 43404 2456
rect 43364 800 43392 2450
rect 43640 800 43668 2858
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 43904 2372 43956 2378
rect 43904 2314 43956 2320
rect 43916 800 43944 2314
rect 44192 800 44220 2790
rect 44456 2576 44508 2582
rect 44456 2518 44508 2524
rect 44468 800 44496 2518
rect 44744 800 44772 2926
rect 45020 800 45048 3470
rect 45296 800 45324 3470
rect 45560 2848 45612 2854
rect 45560 2790 45612 2796
rect 45572 800 45600 2790
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 45848 800 45876 2382
rect 46124 800 46152 3470
rect 46664 2848 46716 2854
rect 46664 2790 46716 2796
rect 46388 2508 46440 2514
rect 46388 2450 46440 2456
rect 46400 800 46428 2450
rect 46676 800 46704 2790
rect 46952 800 46980 3470
rect 47492 2916 47544 2922
rect 47492 2858 47544 2864
rect 47216 2372 47268 2378
rect 47216 2314 47268 2320
rect 47228 800 47256 2314
rect 47504 800 47532 2858
rect 47780 800 47808 3470
rect 48596 2984 48648 2990
rect 48596 2926 48648 2932
rect 48044 2848 48096 2854
rect 48044 2790 48096 2796
rect 48056 800 48084 2790
rect 48320 2576 48372 2582
rect 48320 2518 48372 2524
rect 48332 800 48360 2518
rect 48608 800 48636 2926
rect 48884 800 48912 3470
rect 49424 2916 49476 2922
rect 49424 2858 49476 2864
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 49160 800 49188 2450
rect 49436 800 49464 2858
rect 49976 2848 50028 2854
rect 49976 2790 50028 2796
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 49712 800 49740 2382
rect 49988 800 50016 2790
rect 50172 1850 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50620 2916 50672 2922
rect 50620 2858 50672 2864
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50172 1822 50292 1850
rect 50264 800 50292 1822
rect 50632 1442 50660 2858
rect 50540 1414 50660 1442
rect 50540 800 50568 1414
rect 50816 800 50844 3470
rect 51080 2508 51132 2514
rect 51080 2450 51132 2456
rect 51092 800 51120 2450
rect 51368 800 51396 3470
rect 52460 2984 52512 2990
rect 52460 2926 52512 2932
rect 51908 2848 51960 2854
rect 51908 2790 51960 2796
rect 51632 2440 51684 2446
rect 51632 2382 51684 2388
rect 51644 800 51672 2382
rect 51920 800 51948 2790
rect 52184 2576 52236 2582
rect 52184 2518 52236 2524
rect 52196 800 52224 2518
rect 52472 800 52500 2926
rect 52748 800 52776 3470
rect 53024 800 53052 3470
rect 53564 2984 53616 2990
rect 53564 2926 53616 2932
rect 53288 2916 53340 2922
rect 53288 2858 53340 2864
rect 53300 800 53328 2858
rect 53576 800 53604 2926
rect 54392 2916 54444 2922
rect 54392 2858 54444 2864
rect 53840 2848 53892 2854
rect 53840 2790 53892 2796
rect 53852 800 53880 2790
rect 54116 2372 54168 2378
rect 54116 2314 54168 2320
rect 54128 800 54156 2314
rect 54404 800 54432 2858
rect 54680 800 54708 3470
rect 55220 2984 55272 2990
rect 55220 2926 55272 2932
rect 55232 2650 55260 2926
rect 55404 2848 55456 2854
rect 55404 2790 55456 2796
rect 55220 2644 55272 2650
rect 55220 2586 55272 2592
rect 54944 2508 54996 2514
rect 54944 2450 54996 2456
rect 54956 800 54984 2450
rect 55416 1442 55444 2790
rect 55232 1414 55444 1442
rect 55232 800 55260 1414
rect 55508 800 55536 3470
rect 55680 2916 55732 2922
rect 55680 2858 55732 2864
rect 55692 800 55720 2858
rect 55784 800 55812 3538
rect 55956 3188 56008 3194
rect 55956 3130 56008 3136
rect 55864 2576 55916 2582
rect 55864 2518 55916 2524
rect 55876 800 55904 2518
rect 55968 800 55996 3130
rect 56048 2848 56100 2854
rect 56048 2790 56100 2796
rect 56060 800 56088 2790
rect 56152 800 56180 3878
rect 56232 3528 56284 3534
rect 56232 3470 56284 3476
rect 56244 800 56272 3470
rect 56336 800 56364 3878
rect 56508 3664 56560 3670
rect 56508 3606 56560 3612
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 56428 800 56456 2382
rect 56520 800 56548 3606
rect 56784 3596 56836 3602
rect 56784 3538 56836 3544
rect 56692 2984 56744 2990
rect 56692 2926 56744 2932
rect 56704 1442 56732 2926
rect 56612 1414 56732 1442
rect 56612 800 56640 1414
rect 56796 1306 56824 3538
rect 56876 2304 56928 2310
rect 56876 2246 56928 2252
rect 56704 1278 56824 1306
rect 56704 800 56732 1278
rect 56784 1216 56836 1222
rect 56784 1158 56836 1164
rect 56796 800 56824 1158
rect 56888 800 56916 2246
rect 56980 800 57008 3878
rect 57060 2916 57112 2922
rect 57060 2858 57112 2864
rect 57072 1222 57100 2858
rect 57060 1216 57112 1222
rect 57060 1158 57112 1164
rect 57060 1080 57112 1086
rect 57060 1022 57112 1028
rect 57072 800 57100 1022
rect 57164 800 57192 4558
rect 57256 800 57284 4694
rect 57612 4616 57664 4622
rect 57612 4558 57664 4564
rect 57520 4004 57572 4010
rect 57520 3946 57572 3952
rect 57336 3528 57388 3534
rect 57336 3470 57388 3476
rect 57348 800 57376 3470
rect 57428 2644 57480 2650
rect 57428 2586 57480 2592
rect 57440 800 57468 2586
rect 57532 800 57560 3946
rect 57624 800 57652 4558
rect 57980 4140 58032 4146
rect 57980 4082 58032 4088
rect 57796 3732 57848 3738
rect 57796 3674 57848 3680
rect 57704 3120 57756 3126
rect 57704 3062 57756 3068
rect 57716 800 57744 3062
rect 57808 800 57836 3674
rect 57886 3224 57942 3233
rect 57886 3159 57942 3168
rect 57900 800 57928 3159
rect 57992 800 58020 4082
rect 58072 3936 58124 3942
rect 58072 3878 58124 3884
rect 58084 3738 58112 3878
rect 58072 3732 58124 3738
rect 58072 3674 58124 3680
rect 58072 3188 58124 3194
rect 58072 3130 58124 3136
rect 58084 2582 58112 3130
rect 58164 3052 58216 3058
rect 58164 2994 58216 3000
rect 58072 2576 58124 2582
rect 58072 2518 58124 2524
rect 58072 2100 58124 2106
rect 58072 2042 58124 2048
rect 58084 800 58112 2042
rect 58176 800 58204 2994
rect 58268 800 58296 4694
rect 58624 4004 58676 4010
rect 58624 3946 58676 3952
rect 58348 3664 58400 3670
rect 58348 3606 58400 3612
rect 58360 800 58388 3606
rect 58440 2984 58492 2990
rect 58440 2926 58492 2932
rect 58452 800 58480 2926
rect 58532 1964 58584 1970
rect 58532 1906 58584 1912
rect 58544 800 58572 1906
rect 58636 800 58664 3946
rect 58728 800 58756 4966
rect 58820 800 58848 5102
rect 59268 5092 59320 5098
rect 59268 5034 59320 5040
rect 58900 4684 58952 4690
rect 58900 4626 58952 4632
rect 58912 800 58940 4626
rect 59176 4072 59228 4078
rect 59176 4014 59228 4020
rect 58992 3596 59044 3602
rect 58992 3538 59044 3544
rect 59004 800 59032 3538
rect 59084 2032 59136 2038
rect 59084 1974 59136 1980
rect 59096 800 59124 1974
rect 59188 800 59216 4014
rect 59280 800 59308 5034
rect 67640 5024 67692 5030
rect 67640 4966 67692 4972
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 67652 4865 67680 4966
rect 67638 4856 67694 4865
rect 67638 4791 67694 4800
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 60464 3528 60516 3534
rect 68100 3528 68152 3534
rect 60464 3470 60516 3476
rect 68098 3496 68100 3505
rect 68152 3496 68154 3505
rect 60476 3233 60504 3470
rect 68098 3431 68154 3440
rect 60462 3224 60518 3233
rect 60462 3159 60518 3168
rect 60464 3120 60516 3126
rect 60464 3062 60516 3068
rect 59360 2916 59412 2922
rect 59360 2858 59412 2864
rect 59372 800 59400 2858
rect 60476 2854 60504 3062
rect 59452 2848 59504 2854
rect 59452 2790 59504 2796
rect 60464 2848 60516 2854
rect 60464 2790 60516 2796
rect 59464 1086 59492 2790
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 63684 2508 63736 2514
rect 63684 2450 63736 2456
rect 61752 2440 61804 2446
rect 61752 2382 61804 2388
rect 63040 2440 63092 2446
rect 63040 2382 63092 2388
rect 61764 2106 61792 2382
rect 61752 2100 61804 2106
rect 61752 2042 61804 2048
rect 63052 1970 63080 2382
rect 63696 2038 63724 2450
rect 66996 2440 67048 2446
rect 66996 2382 67048 2388
rect 67548 2440 67600 2446
rect 67548 2382 67600 2388
rect 67008 2145 67036 2382
rect 66994 2136 67050 2145
rect 66994 2071 67050 2080
rect 63684 2032 63736 2038
rect 63684 1974 63736 1980
rect 63040 1964 63092 1970
rect 63040 1906 63092 1912
rect 59452 1080 59504 1086
rect 59452 1022 59504 1028
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54758 0 54814 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55034 0 55090 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55310 0 55366 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55862 0 55918 800
rect 55954 0 56010 800
rect 56046 0 56102 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56598 0 56654 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56874 0 56930 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57150 0 57206 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57610 0 57666 800
rect 57702 0 57758 800
rect 57794 0 57850 800
rect 57886 0 57942 800
rect 57978 0 58034 800
rect 58070 0 58126 800
rect 58162 0 58218 800
rect 58254 0 58310 800
rect 58346 0 58402 800
rect 58438 0 58494 800
rect 58530 0 58586 800
rect 58622 0 58678 800
rect 58714 0 58770 800
rect 58806 0 58862 800
rect 58898 0 58954 800
rect 58990 0 59046 800
rect 59082 0 59138 800
rect 59174 0 59230 800
rect 59266 0 59322 800
rect 59358 0 59414 800
rect 67560 785 67588 2382
rect 67546 776 67602 785
rect 67546 711 67602 720
<< via2 >>
rect 67546 59200 67602 59256
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 66994 57840 67050 57896
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 68098 56480 68154 56536
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 67638 55140 67694 55176
rect 67638 55120 67640 55140
rect 67640 55120 67692 55140
rect 67692 55120 67694 55140
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 67546 53760 67602 53816
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 68098 52436 68100 52456
rect 68100 52436 68152 52456
rect 68152 52436 68154 52456
rect 68098 52400 68154 52436
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 68098 51040 68154 51096
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 67638 49716 67640 49736
rect 67640 49716 67692 49736
rect 67692 49716 67694 49736
rect 67638 49680 67694 49716
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 67638 48320 67694 48376
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 68098 46996 68100 47016
rect 68100 46996 68152 47016
rect 68152 46996 68154 47016
rect 68098 46960 68154 46996
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 68098 45600 68154 45656
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 67638 44260 67694 44296
rect 67638 44240 67640 44260
rect 67640 44240 67692 44260
rect 67692 44240 67694 44260
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 67638 42880 67694 42936
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 68098 41556 68100 41576
rect 68100 41556 68152 41576
rect 68152 41556 68154 41576
rect 68098 41520 68154 41556
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 68098 40160 68154 40216
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 67638 38820 67694 38856
rect 67638 38800 67640 38820
rect 67640 38800 67692 38820
rect 67692 38800 67694 38820
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 67638 37440 67694 37496
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 68098 36116 68100 36136
rect 68100 36116 68152 36136
rect 68152 36116 68154 36136
rect 68098 36080 68154 36116
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 68098 34720 68154 34776
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 67638 33380 67694 33416
rect 67638 33360 67640 33380
rect 67640 33360 67692 33380
rect 67692 33360 67694 33380
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 67638 32000 67694 32056
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 9770 30676 9772 30696
rect 9772 30676 9824 30696
rect 9824 30676 9826 30696
rect 9770 30640 9826 30676
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 2594 18808 2650 18864
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 2502 17312 2558 17368
rect 2134 3984 2190 4040
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 3790 16224 3846 16280
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 2962 3476 2964 3496
rect 2964 3476 3016 3496
rect 3016 3476 3018 3496
rect 2962 3440 3018 3476
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3422 4256 3478 4312
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3882 3440 3938 3496
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5538 19760 5594 19816
rect 5446 18672 5502 18728
rect 7194 21800 7250 21856
rect 6642 19388 6644 19408
rect 6644 19388 6696 19408
rect 6696 19388 6698 19408
rect 6642 19352 6698 19388
rect 5906 17176 5962 17232
rect 7378 16360 7434 16416
rect 7654 15700 7710 15736
rect 7654 15680 7656 15700
rect 7656 15680 7708 15700
rect 7708 15680 7710 15700
rect 5630 10648 5686 10704
rect 4710 4664 4766 4720
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4618 3032 4674 3088
rect 1950 1808 2006 1864
rect 3054 2080 3110 2136
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5814 3984 5870 4040
rect 4066 1944 4122 2000
rect 6274 3032 6330 3088
rect 11978 30676 11980 30696
rect 11980 30676 12032 30696
rect 12032 30676 12034 30696
rect 11978 30640 12034 30676
rect 12162 29300 12218 29336
rect 12162 29280 12164 29300
rect 12164 29280 12216 29300
rect 12216 29280 12218 29300
rect 10322 27784 10378 27840
rect 10782 27668 10838 27704
rect 10782 27648 10784 27668
rect 10784 27648 10836 27668
rect 10836 27648 10838 27668
rect 9678 21936 9734 21992
rect 9402 21800 9458 21856
rect 9310 21528 9366 21584
rect 9310 21392 9366 21448
rect 9586 21392 9642 21448
rect 10598 21528 10654 21584
rect 8942 19352 8998 19408
rect 10598 19760 10654 19816
rect 9770 16244 9826 16280
rect 9770 16224 9772 16244
rect 9772 16224 9824 16244
rect 9824 16224 9826 16244
rect 8390 15952 8446 16008
rect 7654 8336 7710 8392
rect 9494 15580 9496 15600
rect 9496 15580 9548 15600
rect 9548 15580 9550 15600
rect 9494 15544 9550 15580
rect 9586 11600 9642 11656
rect 6734 3732 6790 3768
rect 6734 3712 6736 3732
rect 6736 3712 6788 3732
rect 6788 3712 6790 3732
rect 8298 7520 8354 7576
rect 7562 3576 7618 3632
rect 6826 3168 6882 3224
rect 8298 5788 8300 5808
rect 8300 5788 8352 5808
rect 8352 5788 8354 5808
rect 8298 5752 8354 5788
rect 8942 4392 8998 4448
rect 8850 4276 8906 4312
rect 8850 4256 8852 4276
rect 8852 4256 8904 4276
rect 8904 4256 8906 4276
rect 8942 3712 8998 3768
rect 8850 3304 8906 3360
rect 5262 2352 5318 2408
rect 5170 2216 5226 2272
rect 2410 1672 2466 1728
rect 9310 5208 9366 5264
rect 10874 13776 10930 13832
rect 10598 11500 10600 11520
rect 10600 11500 10652 11520
rect 10652 11500 10654 11520
rect 10598 11464 10654 11500
rect 12162 27648 12218 27704
rect 12530 27784 12586 27840
rect 12806 27648 12862 27704
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 11058 11092 11060 11112
rect 11060 11092 11112 11112
rect 11112 11092 11114 11112
rect 11058 11056 11114 11092
rect 9678 4256 9734 4312
rect 9126 3440 9182 3496
rect 10138 3984 10194 4040
rect 10046 3576 10102 3632
rect 9034 1536 9090 1592
rect 10506 4800 10562 4856
rect 10414 4528 10470 4584
rect 10506 4156 10508 4176
rect 10508 4156 10560 4176
rect 10560 4156 10562 4176
rect 10506 4120 10562 4156
rect 10690 6740 10692 6760
rect 10692 6740 10744 6760
rect 10744 6740 10746 6760
rect 10690 6704 10746 6740
rect 10598 3848 10654 3904
rect 10506 3032 10562 3088
rect 10414 2760 10470 2816
rect 10690 3712 10746 3768
rect 11058 7520 11114 7576
rect 10966 6840 11022 6896
rect 10874 3440 10930 3496
rect 10598 2932 10600 2952
rect 10600 2932 10652 2952
rect 10652 2932 10654 2952
rect 10598 2896 10654 2932
rect 10874 2760 10930 2816
rect 12070 10532 12126 10568
rect 12070 10512 12072 10532
rect 12072 10512 12124 10532
rect 12124 10512 12126 10532
rect 11610 4664 11666 4720
rect 11242 2644 11298 2680
rect 11242 2624 11244 2644
rect 11244 2624 11296 2644
rect 11296 2624 11298 2644
rect 11978 4700 11980 4720
rect 11980 4700 12032 4720
rect 12032 4700 12034 4720
rect 11978 4664 12034 4700
rect 11794 3984 11850 4040
rect 12530 23468 12532 23488
rect 12532 23468 12584 23488
rect 12584 23468 12586 23488
rect 12530 23432 12586 23468
rect 12622 18808 12678 18864
rect 12622 17176 12678 17232
rect 12990 14320 13046 14376
rect 12346 12708 12402 12744
rect 12346 12688 12348 12708
rect 12348 12688 12400 12708
rect 12400 12688 12402 12708
rect 12806 13676 12808 13696
rect 12808 13676 12860 13696
rect 12860 13676 12862 13696
rect 12806 13640 12862 13676
rect 12898 13368 12954 13424
rect 13450 19508 13506 19544
rect 13450 19488 13452 19508
rect 13452 19488 13504 19508
rect 13504 19488 13506 19508
rect 13450 15428 13506 15464
rect 13450 15408 13452 15428
rect 13452 15408 13504 15428
rect 13504 15408 13506 15428
rect 13082 12416 13138 12472
rect 13174 12280 13230 12336
rect 13726 19780 13782 19816
rect 13726 19760 13728 19780
rect 13728 19760 13780 19780
rect 13780 19760 13782 19780
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 12530 6704 12586 6760
rect 12346 4800 12402 4856
rect 12714 3848 12770 3904
rect 12622 1672 12678 1728
rect 13174 4664 13230 4720
rect 13082 3576 13138 3632
rect 13266 3884 13268 3904
rect 13268 3884 13320 3904
rect 13320 3884 13322 3904
rect 13266 3848 13322 3884
rect 13266 2896 13322 2952
rect 13174 2080 13230 2136
rect 13082 1944 13138 2000
rect 13450 2916 13506 2952
rect 13450 2896 13452 2916
rect 13452 2896 13504 2916
rect 13504 2896 13506 2916
rect 13450 2760 13506 2816
rect 13818 4392 13874 4448
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 14278 15136 14334 15192
rect 14370 13640 14426 13696
rect 14646 13640 14702 13696
rect 14462 12552 14518 12608
rect 15382 12824 15438 12880
rect 14370 10668 14426 10704
rect 14370 10648 14372 10668
rect 14372 10648 14424 10668
rect 14424 10648 14426 10668
rect 14002 4392 14058 4448
rect 13910 3848 13966 3904
rect 13726 3576 13782 3632
rect 13818 2760 13874 2816
rect 14922 6840 14978 6896
rect 16302 19896 16358 19952
rect 15842 13932 15898 13968
rect 15842 13912 15844 13932
rect 15844 13912 15896 13932
rect 15896 13912 15898 13932
rect 14922 4528 14978 4584
rect 14370 3168 14426 3224
rect 14646 3340 14648 3360
rect 14648 3340 14700 3360
rect 14700 3340 14702 3360
rect 14646 3304 14702 3340
rect 14554 2932 14556 2952
rect 14556 2932 14608 2952
rect 14608 2932 14610 2952
rect 14554 2896 14610 2932
rect 15106 4256 15162 4312
rect 15014 2644 15070 2680
rect 15014 2624 15016 2644
rect 15016 2624 15068 2644
rect 15068 2624 15070 2644
rect 15566 2216 15622 2272
rect 16578 21564 16580 21584
rect 16580 21564 16632 21584
rect 16632 21564 16634 21584
rect 16578 21528 16634 21564
rect 18510 20748 18512 20768
rect 18512 20748 18564 20768
rect 18564 20748 18566 20768
rect 18510 20712 18566 20748
rect 18234 19488 18290 19544
rect 17130 12980 17186 13016
rect 17130 12960 17132 12980
rect 17132 12960 17184 12980
rect 17184 12960 17186 12980
rect 17590 13912 17646 13968
rect 16578 12144 16634 12200
rect 16486 11212 16542 11248
rect 16486 11192 16488 11212
rect 16488 11192 16540 11212
rect 16540 11192 16542 11212
rect 17314 10920 17370 10976
rect 17222 10648 17278 10704
rect 17866 12960 17922 13016
rect 18694 18964 18750 19000
rect 18694 18944 18696 18964
rect 18696 18944 18748 18964
rect 18748 18944 18750 18964
rect 18694 16632 18750 16688
rect 16118 3576 16174 3632
rect 16578 4120 16634 4176
rect 17590 5752 17646 5808
rect 17682 5208 17738 5264
rect 17590 2488 17646 2544
rect 18878 20884 18880 20904
rect 18880 20884 18932 20904
rect 18932 20884 18934 20904
rect 18878 20848 18934 20884
rect 18970 17312 19026 17368
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19706 26324 19708 26344
rect 19708 26324 19760 26344
rect 19760 26324 19762 26344
rect 19706 26288 19762 26324
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19338 24012 19340 24032
rect 19340 24012 19392 24032
rect 19392 24012 19394 24032
rect 19338 23976 19394 24012
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19338 23160 19394 23216
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19338 20440 19394 20496
rect 19246 17176 19302 17232
rect 18878 13388 18934 13424
rect 18878 13368 18880 13388
rect 18880 13368 18932 13388
rect 18932 13368 18934 13388
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20350 24012 20352 24032
rect 20352 24012 20404 24032
rect 20404 24012 20406 24032
rect 20350 23976 20406 24012
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19982 17196 20038 17232
rect 19982 17176 19984 17196
rect 19984 17176 20036 17196
rect 20036 17176 20038 17196
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 22834 26444 22890 26480
rect 22834 26424 22836 26444
rect 22836 26424 22888 26444
rect 22888 26424 22890 26444
rect 20534 21956 20590 21992
rect 20534 21936 20536 21956
rect 20536 21936 20588 21956
rect 20588 21936 20590 21956
rect 20442 19488 20498 19544
rect 21270 20712 21326 20768
rect 22466 23840 22522 23896
rect 21546 21664 21602 21720
rect 20534 17720 20590 17776
rect 20534 16496 20590 16552
rect 20350 16088 20406 16144
rect 20074 15544 20130 15600
rect 19982 15272 20038 15328
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20074 15136 20130 15192
rect 20534 15852 20536 15872
rect 20536 15852 20588 15872
rect 20588 15852 20590 15872
rect 20534 15816 20590 15852
rect 20166 14864 20222 14920
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 20074 14220 20076 14240
rect 20076 14220 20128 14240
rect 20128 14220 20130 14240
rect 20074 14184 20130 14220
rect 20166 14048 20222 14104
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19430 12044 19432 12064
rect 19432 12044 19484 12064
rect 19484 12044 19486 12064
rect 19430 12008 19486 12044
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19706 11772 19708 11792
rect 19708 11772 19760 11792
rect 19760 11772 19762 11792
rect 19706 11736 19762 11772
rect 19798 11328 19854 11384
rect 19982 11056 20038 11112
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 17866 2760 17922 2816
rect 19890 9324 19892 9344
rect 19892 9324 19944 9344
rect 19944 9324 19946 9344
rect 19890 9288 19946 9324
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 18234 4392 18290 4448
rect 18234 2352 18290 2408
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20718 15680 20774 15736
rect 20994 16396 20996 16416
rect 20996 16396 21048 16416
rect 21048 16396 21050 16416
rect 20994 16360 21050 16396
rect 21362 15952 21418 16008
rect 22098 19796 22100 19816
rect 22100 19796 22152 19816
rect 22152 19796 22154 19816
rect 22098 19760 22154 19796
rect 21546 15816 21602 15872
rect 20534 14184 20590 14240
rect 21086 13368 21142 13424
rect 21914 17584 21970 17640
rect 23018 22208 23074 22264
rect 22650 20440 22706 20496
rect 22466 18164 22468 18184
rect 22468 18164 22520 18184
rect 22520 18164 22522 18184
rect 22466 18128 22522 18164
rect 23110 20848 23166 20904
rect 22190 16496 22246 16552
rect 20074 6196 20076 6216
rect 20076 6196 20128 6216
rect 20128 6196 20130 6216
rect 20074 6160 20130 6196
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19890 3732 19946 3768
rect 19890 3712 19892 3732
rect 19892 3712 19944 3732
rect 19944 3712 19946 3732
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20534 9288 20590 9344
rect 21730 12824 21786 12880
rect 22374 15700 22430 15736
rect 22374 15680 22376 15700
rect 22376 15680 22428 15700
rect 22428 15680 22430 15700
rect 22374 15308 22376 15328
rect 22376 15308 22428 15328
rect 22428 15308 22430 15328
rect 22374 15272 22430 15308
rect 22098 13776 22154 13832
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 68098 30676 68100 30696
rect 68100 30676 68152 30696
rect 68152 30676 68154 30696
rect 68098 30640 68154 30676
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 24214 26424 24270 26480
rect 23386 18808 23442 18864
rect 23202 18128 23258 18184
rect 22282 11736 22338 11792
rect 21454 7828 21456 7848
rect 21456 7828 21508 7848
rect 21508 7828 21510 7848
rect 21454 7792 21510 7828
rect 23386 15408 23442 15464
rect 23478 15272 23534 15328
rect 24858 22208 24914 22264
rect 24122 11328 24178 11384
rect 24398 15136 24454 15192
rect 25502 23180 25558 23216
rect 25502 23160 25504 23180
rect 25504 23160 25556 23180
rect 25556 23160 25558 23180
rect 25042 19896 25098 19952
rect 24766 14884 24822 14920
rect 24766 14864 24768 14884
rect 24768 14864 24820 14884
rect 24820 14864 24822 14884
rect 25778 26444 25834 26480
rect 25778 26424 25780 26444
rect 25780 26424 25832 26444
rect 25832 26424 25834 26444
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 68098 29280 68154 29336
rect 27066 26308 27122 26344
rect 27066 26288 27068 26308
rect 27068 26288 27120 26308
rect 27120 26288 27122 26308
rect 25410 16360 25466 16416
rect 25226 14320 25282 14376
rect 25502 14048 25558 14104
rect 24582 11892 24638 11928
rect 24582 11872 24584 11892
rect 24584 11872 24636 11892
rect 24636 11872 24638 11892
rect 22926 8880 22982 8936
rect 25778 18164 25780 18184
rect 25780 18164 25832 18184
rect 25832 18164 25834 18184
rect 25778 18128 25834 18164
rect 28170 23860 28226 23896
rect 28170 23840 28172 23860
rect 28172 23840 28224 23860
rect 28224 23840 28226 23860
rect 26974 21664 27030 21720
rect 26514 20460 26570 20496
rect 26514 20440 26516 20460
rect 26516 20440 26568 20460
rect 26568 20440 26570 20460
rect 26514 19488 26570 19544
rect 30470 28364 30472 28384
rect 30472 28364 30524 28384
rect 30524 28364 30526 28384
rect 30470 28328 30526 28364
rect 30378 28192 30434 28248
rect 28170 19796 28172 19816
rect 28172 19796 28224 19816
rect 28224 19796 28226 19816
rect 28170 19760 28226 19796
rect 25594 12144 25650 12200
rect 25042 11464 25098 11520
rect 20994 6160 21050 6216
rect 25962 11600 26018 11656
rect 29090 17720 29146 17776
rect 29550 17584 29606 17640
rect 29458 16632 29514 16688
rect 28078 16088 28134 16144
rect 28630 15308 28632 15328
rect 28632 15308 28684 15328
rect 28684 15308 28686 15328
rect 28630 15272 28686 15308
rect 27526 13368 27582 13424
rect 27434 12552 27490 12608
rect 20902 3848 20958 3904
rect 28262 14184 28318 14240
rect 28998 12688 29054 12744
rect 28446 6296 28502 6352
rect 30746 28328 30802 28384
rect 30838 28192 30894 28248
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 67638 27940 67694 27976
rect 67638 27920 67640 27940
rect 67640 27920 67692 27940
rect 67692 27920 67694 27940
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 67638 26560 67694 26616
rect 29826 16516 29882 16552
rect 29826 16496 29828 16516
rect 29828 16496 29880 16516
rect 29880 16496 29882 16516
rect 30838 17720 30894 17776
rect 30654 16632 30710 16688
rect 30010 13252 30066 13288
rect 30010 13232 30012 13252
rect 30012 13232 30064 13252
rect 30064 13232 30066 13252
rect 30286 12436 30342 12472
rect 30286 12416 30288 12436
rect 30288 12416 30340 12436
rect 30340 12416 30342 12436
rect 29642 11228 29644 11248
rect 29644 11228 29696 11248
rect 29696 11228 29698 11248
rect 29642 11192 29698 11228
rect 29550 10512 29606 10568
rect 30010 10648 30066 10704
rect 30746 15680 30802 15736
rect 32310 16632 32366 16688
rect 32586 15816 32642 15872
rect 31390 11328 31446 11384
rect 31666 11192 31722 11248
rect 33322 15272 33378 15328
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 68098 25236 68100 25256
rect 68100 25236 68152 25256
rect 68152 25236 68154 25256
rect 68098 25200 68154 25236
rect 33782 15272 33838 15328
rect 32494 8880 32550 8936
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 68098 23840 68154 23896
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 67638 22500 67694 22536
rect 67638 22480 67640 22500
rect 67640 22480 67692 22500
rect 67692 22480 67694 22500
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 36174 20576 36230 20632
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 32678 6316 32734 6352
rect 32678 6296 32680 6316
rect 32680 6296 32732 6316
rect 32732 6296 32734 6316
rect 34426 11328 34482 11384
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 36266 16496 36322 16552
rect 36082 13232 36138 13288
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 38842 20576 38898 20632
rect 38842 14356 38844 14376
rect 38844 14356 38896 14376
rect 38896 14356 38898 14376
rect 38842 14320 38898 14356
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 67638 21120 67694 21176
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 37554 11228 37556 11248
rect 37556 11228 37608 11248
rect 37608 11228 37610 11248
rect 37554 11192 37610 11228
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 68098 19796 68100 19816
rect 68100 19796 68152 19816
rect 68152 19796 68154 19816
rect 68098 19760 68154 19796
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 68098 18400 68154 18456
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 67638 17060 67694 17096
rect 67638 17040 67640 17060
rect 67640 17040 67692 17060
rect 67692 17040 67694 17060
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 67638 15680 67694 15736
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 40498 14340 40554 14376
rect 40498 14320 40500 14340
rect 40500 14320 40552 14340
rect 40552 14320 40554 14340
rect 68098 14356 68100 14376
rect 68100 14356 68152 14376
rect 68152 14356 68154 14376
rect 68098 14320 68154 14356
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 68098 12960 68154 13016
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 67638 11620 67694 11656
rect 67638 11600 67640 11620
rect 67640 11600 67692 11620
rect 67692 11600 67694 11620
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 67638 10240 67694 10296
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 68098 8916 68100 8936
rect 68100 8916 68152 8936
rect 68152 8916 68154 8936
rect 68098 8880 68154 8916
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 68098 7520 68154 7576
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 67638 6180 67694 6216
rect 67638 6160 67640 6180
rect 67640 6160 67692 6180
rect 67692 6160 67694 6180
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 57886 3168 57942 3224
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 67638 4800 67694 4856
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 68098 3476 68100 3496
rect 68100 3476 68152 3496
rect 68152 3476 68154 3496
rect 68098 3440 68154 3476
rect 60462 3168 60518 3224
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 66994 2080 67050 2136
rect 67546 720 67602 776
<< metal3 >>
rect 67541 59258 67607 59261
rect 69200 59258 70000 59288
rect 67541 59256 70000 59258
rect 67541 59200 67546 59256
rect 67602 59200 70000 59256
rect 67541 59198 70000 59200
rect 67541 59195 67607 59198
rect 69200 59168 70000 59198
rect 66989 57898 67055 57901
rect 69200 57898 70000 57928
rect 66989 57896 70000 57898
rect 66989 57840 66994 57896
rect 67050 57840 70000 57896
rect 66989 57838 70000 57840
rect 66989 57835 67055 57838
rect 69200 57808 70000 57838
rect 19570 57696 19886 57697
rect 0 57536 800 57656
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 68093 56538 68159 56541
rect 69200 56538 70000 56568
rect 68093 56536 70000 56538
rect 68093 56480 68098 56536
rect 68154 56480 70000 56536
rect 68093 56478 70000 56480
rect 68093 56475 68159 56478
rect 69200 56448 70000 56478
rect 0 56040 800 56160
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 65650 55999 65966 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 67633 55178 67699 55181
rect 69200 55178 70000 55208
rect 67633 55176 70000 55178
rect 67633 55120 67638 55176
rect 67694 55120 70000 55176
rect 67633 55118 70000 55120
rect 67633 55115 67699 55118
rect 69200 55088 70000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 0 54544 800 54664
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 67541 53818 67607 53821
rect 69200 53818 70000 53848
rect 67541 53816 70000 53818
rect 67541 53760 67546 53816
rect 67602 53760 70000 53816
rect 67541 53758 70000 53760
rect 67541 53755 67607 53758
rect 69200 53728 70000 53758
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 0 53048 800 53168
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 68093 52458 68159 52461
rect 69200 52458 70000 52488
rect 68093 52456 70000 52458
rect 68093 52400 68098 52456
rect 68154 52400 70000 52456
rect 68093 52398 70000 52400
rect 68093 52395 68159 52398
rect 69200 52368 70000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51552 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 68093 51098 68159 51101
rect 69200 51098 70000 51128
rect 68093 51096 70000 51098
rect 68093 51040 68098 51096
rect 68154 51040 70000 51096
rect 68093 51038 70000 51040
rect 68093 51035 68159 51038
rect 69200 51008 70000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 0 50056 800 50176
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 67633 49738 67699 49741
rect 69200 49738 70000 49768
rect 67633 49736 70000 49738
rect 67633 49680 67638 49736
rect 67694 49680 70000 49736
rect 67633 49678 70000 49680
rect 67633 49675 67699 49678
rect 69200 49648 70000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48560 800 48680
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 67633 48378 67699 48381
rect 69200 48378 70000 48408
rect 67633 48376 70000 48378
rect 67633 48320 67638 48376
rect 67694 48320 70000 48376
rect 67633 48318 70000 48320
rect 67633 48315 67699 48318
rect 69200 48288 70000 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 0 47064 800 47184
rect 68093 47018 68159 47021
rect 69200 47018 70000 47048
rect 68093 47016 70000 47018
rect 68093 46960 68098 47016
rect 68154 46960 70000 47016
rect 68093 46958 70000 46960
rect 68093 46955 68159 46958
rect 69200 46928 70000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 19570 45728 19886 45729
rect 0 45568 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 68093 45658 68159 45661
rect 69200 45658 70000 45688
rect 68093 45656 70000 45658
rect 68093 45600 68098 45656
rect 68154 45600 70000 45656
rect 68093 45598 70000 45600
rect 68093 45595 68159 45598
rect 69200 45568 70000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 67633 44298 67699 44301
rect 69200 44298 70000 44328
rect 67633 44296 70000 44298
rect 67633 44240 67638 44296
rect 67694 44240 70000 44296
rect 67633 44238 70000 44240
rect 67633 44235 67699 44238
rect 69200 44208 70000 44238
rect 0 44072 800 44192
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 67633 42938 67699 42941
rect 69200 42938 70000 42968
rect 67633 42936 70000 42938
rect 67633 42880 67638 42936
rect 67694 42880 70000 42936
rect 67633 42878 70000 42880
rect 67633 42875 67699 42878
rect 69200 42848 70000 42878
rect 0 42576 800 42696
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 68093 41578 68159 41581
rect 69200 41578 70000 41608
rect 68093 41576 70000 41578
rect 68093 41520 68098 41576
rect 68154 41520 70000 41576
rect 68093 41518 70000 41520
rect 68093 41515 68159 41518
rect 69200 41488 70000 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41080 800 41200
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 68093 40218 68159 40221
rect 69200 40218 70000 40248
rect 68093 40216 70000 40218
rect 68093 40160 68098 40216
rect 68154 40160 70000 40216
rect 68093 40158 70000 40160
rect 68093 40155 68159 40158
rect 69200 40128 70000 40158
rect 4210 39744 4526 39745
rect 0 39584 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 67633 38858 67699 38861
rect 69200 38858 70000 38888
rect 67633 38856 70000 38858
rect 67633 38800 67638 38856
rect 67694 38800 70000 38856
rect 67633 38798 70000 38800
rect 67633 38795 67699 38798
rect 69200 38768 70000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 0 38088 800 38208
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 67633 37498 67699 37501
rect 69200 37498 70000 37528
rect 67633 37496 70000 37498
rect 67633 37440 67638 37496
rect 67694 37440 70000 37496
rect 67633 37438 70000 37440
rect 67633 37435 67699 37438
rect 69200 37408 70000 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36592 800 36712
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 68093 36138 68159 36141
rect 69200 36138 70000 36168
rect 68093 36136 70000 36138
rect 68093 36080 68098 36136
rect 68154 36080 70000 36136
rect 68093 36078 70000 36080
rect 68093 36075 68159 36078
rect 69200 36048 70000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 0 35096 800 35216
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 68093 34778 68159 34781
rect 69200 34778 70000 34808
rect 68093 34776 70000 34778
rect 68093 34720 68098 34776
rect 68154 34720 70000 34776
rect 68093 34718 70000 34720
rect 68093 34715 68159 34718
rect 69200 34688 70000 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 19570 33760 19886 33761
rect 0 33600 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 67633 33418 67699 33421
rect 69200 33418 70000 33448
rect 67633 33416 70000 33418
rect 67633 33360 67638 33416
rect 67694 33360 70000 33416
rect 67633 33358 70000 33360
rect 67633 33355 67699 33358
rect 69200 33328 70000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32104 800 32224
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 67633 32058 67699 32061
rect 69200 32058 70000 32088
rect 67633 32056 70000 32058
rect 67633 32000 67638 32056
rect 67694 32000 70000 32056
rect 67633 31998 70000 32000
rect 67633 31995 67699 31998
rect 69200 31968 70000 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 0 30608 800 30728
rect 9765 30698 9831 30701
rect 11973 30698 12039 30701
rect 9765 30696 12039 30698
rect 9765 30640 9770 30696
rect 9826 30640 11978 30696
rect 12034 30640 12039 30696
rect 9765 30638 12039 30640
rect 9765 30635 9831 30638
rect 11973 30635 12039 30638
rect 68093 30698 68159 30701
rect 69200 30698 70000 30728
rect 68093 30696 70000 30698
rect 68093 30640 68098 30696
rect 68154 30640 70000 30696
rect 68093 30638 70000 30640
rect 68093 30635 68159 30638
rect 69200 30608 70000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 12157 29340 12223 29341
rect 12157 29336 12204 29340
rect 12268 29338 12274 29340
rect 68093 29338 68159 29341
rect 69200 29338 70000 29368
rect 12157 29280 12162 29336
rect 12157 29276 12204 29280
rect 12268 29278 12314 29338
rect 68093 29336 70000 29338
rect 68093 29280 68098 29336
rect 68154 29280 70000 29336
rect 68093 29278 70000 29280
rect 12268 29276 12274 29278
rect 12157 29275 12223 29276
rect 68093 29275 68159 29278
rect 69200 29248 70000 29278
rect 0 29112 800 29232
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 30465 28386 30531 28389
rect 30741 28386 30807 28389
rect 30465 28384 30807 28386
rect 30465 28328 30470 28384
rect 30526 28328 30746 28384
rect 30802 28328 30807 28384
rect 30465 28326 30807 28328
rect 30465 28323 30531 28326
rect 30741 28323 30807 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 30373 28250 30439 28253
rect 30833 28250 30899 28253
rect 30373 28248 30899 28250
rect 30373 28192 30378 28248
rect 30434 28192 30838 28248
rect 30894 28192 30899 28248
rect 30373 28190 30899 28192
rect 30373 28187 30439 28190
rect 30833 28187 30899 28190
rect 67633 27978 67699 27981
rect 69200 27978 70000 28008
rect 67633 27976 70000 27978
rect 67633 27920 67638 27976
rect 67694 27920 70000 27976
rect 67633 27918 70000 27920
rect 67633 27915 67699 27918
rect 69200 27888 70000 27918
rect 10317 27842 10383 27845
rect 12525 27842 12591 27845
rect 10317 27840 12591 27842
rect 10317 27784 10322 27840
rect 10378 27784 12530 27840
rect 12586 27784 12591 27840
rect 10317 27782 12591 27784
rect 10317 27779 10383 27782
rect 12525 27779 12591 27782
rect 4210 27776 4526 27777
rect 0 27616 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 10777 27706 10843 27709
rect 12157 27706 12223 27709
rect 10777 27704 12223 27706
rect 10777 27648 10782 27704
rect 10838 27648 12162 27704
rect 12218 27648 12223 27704
rect 10777 27646 12223 27648
rect 10777 27643 10843 27646
rect 12157 27643 12223 27646
rect 12801 27706 12867 27709
rect 12934 27706 12940 27708
rect 12801 27704 12940 27706
rect 12801 27648 12806 27704
rect 12862 27648 12940 27704
rect 12801 27646 12940 27648
rect 12801 27643 12867 27646
rect 12934 27644 12940 27646
rect 13004 27644 13010 27708
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 67633 26618 67699 26621
rect 69200 26618 70000 26648
rect 67633 26616 70000 26618
rect 67633 26560 67638 26616
rect 67694 26560 70000 26616
rect 67633 26558 70000 26560
rect 67633 26555 67699 26558
rect 69200 26528 70000 26558
rect 22829 26482 22895 26485
rect 24209 26482 24275 26485
rect 25773 26482 25839 26485
rect 22829 26480 25839 26482
rect 22829 26424 22834 26480
rect 22890 26424 24214 26480
rect 24270 26424 25778 26480
rect 25834 26424 25839 26480
rect 22829 26422 25839 26424
rect 22829 26419 22895 26422
rect 24209 26419 24275 26422
rect 25773 26419 25839 26422
rect 19701 26346 19767 26349
rect 27061 26346 27127 26349
rect 19701 26344 27127 26346
rect 19701 26288 19706 26344
rect 19762 26288 27066 26344
rect 27122 26288 27127 26344
rect 19701 26286 27127 26288
rect 19701 26283 19767 26286
rect 27061 26283 27127 26286
rect 0 26120 800 26240
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 68093 25258 68159 25261
rect 69200 25258 70000 25288
rect 68093 25256 70000 25258
rect 68093 25200 68098 25256
rect 68154 25200 70000 25256
rect 68093 25198 70000 25200
rect 68093 25195 68159 25198
rect 69200 25168 70000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24624 800 24744
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 19333 24036 19399 24037
rect 19333 24034 19380 24036
rect 19288 24032 19380 24034
rect 19288 23976 19338 24032
rect 19288 23974 19380 23976
rect 19333 23972 19380 23974
rect 19444 23972 19450 24036
rect 20110 23972 20116 24036
rect 20180 24034 20186 24036
rect 20345 24034 20411 24037
rect 20180 24032 20411 24034
rect 20180 23976 20350 24032
rect 20406 23976 20411 24032
rect 20180 23974 20411 23976
rect 20180 23972 20186 23974
rect 19333 23971 19399 23972
rect 20345 23971 20411 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 22461 23898 22527 23901
rect 28165 23898 28231 23901
rect 22461 23896 28231 23898
rect 22461 23840 22466 23896
rect 22522 23840 28170 23896
rect 28226 23840 28231 23896
rect 22461 23838 28231 23840
rect 22461 23835 22527 23838
rect 28165 23835 28231 23838
rect 68093 23898 68159 23901
rect 69200 23898 70000 23928
rect 68093 23896 70000 23898
rect 68093 23840 68098 23896
rect 68154 23840 70000 23896
rect 68093 23838 70000 23840
rect 68093 23835 68159 23838
rect 69200 23808 70000 23838
rect 12525 23490 12591 23493
rect 14406 23490 14412 23492
rect 12525 23488 14412 23490
rect 12525 23432 12530 23488
rect 12586 23432 14412 23488
rect 12525 23430 14412 23432
rect 12525 23427 12591 23430
rect 14406 23428 14412 23430
rect 14476 23428 14482 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 0 23128 800 23248
rect 19333 23218 19399 23221
rect 25497 23218 25563 23221
rect 19333 23216 25563 23218
rect 19333 23160 19338 23216
rect 19394 23160 25502 23216
rect 25558 23160 25563 23216
rect 19333 23158 25563 23160
rect 19333 23155 19399 23158
rect 25497 23155 25563 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 67633 22538 67699 22541
rect 69200 22538 70000 22568
rect 67633 22536 70000 22538
rect 67633 22480 67638 22536
rect 67694 22480 70000 22536
rect 67633 22478 70000 22480
rect 67633 22475 67699 22478
rect 69200 22448 70000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 23013 22266 23079 22269
rect 24853 22266 24919 22269
rect 23013 22264 24919 22266
rect 23013 22208 23018 22264
rect 23074 22208 24858 22264
rect 24914 22208 24919 22264
rect 23013 22206 24919 22208
rect 23013 22203 23079 22206
rect 24853 22203 24919 22206
rect 9673 21994 9739 21997
rect 20529 21994 20595 21997
rect 9673 21992 20595 21994
rect 9673 21936 9678 21992
rect 9734 21936 20534 21992
rect 20590 21936 20595 21992
rect 9673 21934 20595 21936
rect 9673 21931 9739 21934
rect 20529 21931 20595 21934
rect 7189 21858 7255 21861
rect 9397 21858 9463 21861
rect 7189 21856 9463 21858
rect 7189 21800 7194 21856
rect 7250 21800 9402 21856
rect 9458 21800 9463 21856
rect 7189 21798 9463 21800
rect 7189 21795 7255 21798
rect 9397 21795 9463 21798
rect 19570 21792 19886 21793
rect 0 21632 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 21541 21722 21607 21725
rect 26969 21722 27035 21725
rect 21541 21720 27035 21722
rect 21541 21664 21546 21720
rect 21602 21664 26974 21720
rect 27030 21664 27035 21720
rect 21541 21662 27035 21664
rect 21541 21659 21607 21662
rect 26969 21659 27035 21662
rect 9305 21586 9371 21589
rect 10593 21586 10659 21589
rect 16573 21586 16639 21589
rect 9305 21584 16639 21586
rect 9305 21528 9310 21584
rect 9366 21528 10598 21584
rect 10654 21528 16578 21584
rect 16634 21528 16639 21584
rect 9305 21526 16639 21528
rect 9305 21523 9371 21526
rect 10593 21523 10659 21526
rect 16573 21523 16639 21526
rect 9305 21450 9371 21453
rect 9581 21450 9647 21453
rect 9305 21448 9647 21450
rect 9305 21392 9310 21448
rect 9366 21392 9586 21448
rect 9642 21392 9647 21448
rect 9305 21390 9647 21392
rect 9305 21387 9371 21390
rect 9581 21387 9647 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 67633 21178 67699 21181
rect 69200 21178 70000 21208
rect 67633 21176 70000 21178
rect 67633 21120 67638 21176
rect 67694 21120 70000 21176
rect 67633 21118 70000 21120
rect 67633 21115 67699 21118
rect 69200 21088 70000 21118
rect 18873 20906 18939 20909
rect 23105 20906 23171 20909
rect 18873 20904 23171 20906
rect 18873 20848 18878 20904
rect 18934 20848 23110 20904
rect 23166 20848 23171 20904
rect 18873 20846 23171 20848
rect 18873 20843 18939 20846
rect 23105 20843 23171 20846
rect 17166 20708 17172 20772
rect 17236 20770 17242 20772
rect 18505 20770 18571 20773
rect 21265 20770 21331 20773
rect 17236 20768 18571 20770
rect 17236 20712 18510 20768
rect 18566 20712 18571 20768
rect 17236 20710 18571 20712
rect 17236 20708 17242 20710
rect 18505 20707 18571 20710
rect 21222 20768 21331 20770
rect 21222 20712 21270 20768
rect 21326 20712 21331 20768
rect 21222 20707 21331 20712
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 19333 20498 19399 20501
rect 21222 20498 21282 20707
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 36169 20634 36235 20637
rect 38837 20634 38903 20637
rect 36169 20632 38903 20634
rect 36169 20576 36174 20632
rect 36230 20576 38842 20632
rect 38898 20576 38903 20632
rect 36169 20574 38903 20576
rect 36169 20571 36235 20574
rect 38837 20571 38903 20574
rect 19333 20496 21282 20498
rect 19333 20440 19338 20496
rect 19394 20440 21282 20496
rect 19333 20438 21282 20440
rect 22645 20498 22711 20501
rect 26509 20498 26575 20501
rect 22645 20496 26575 20498
rect 22645 20440 22650 20496
rect 22706 20440 26514 20496
rect 26570 20440 26575 20496
rect 22645 20438 26575 20440
rect 19333 20435 19399 20438
rect 22645 20435 22711 20438
rect 26509 20435 26575 20438
rect 0 20136 800 20256
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 16297 19954 16363 19957
rect 25037 19954 25103 19957
rect 16297 19952 25103 19954
rect 16297 19896 16302 19952
rect 16358 19896 25042 19952
rect 25098 19896 25103 19952
rect 16297 19894 25103 19896
rect 16297 19891 16363 19894
rect 25037 19891 25103 19894
rect 5533 19818 5599 19821
rect 10593 19818 10659 19821
rect 13721 19818 13787 19821
rect 5533 19816 13787 19818
rect 5533 19760 5538 19816
rect 5594 19760 10598 19816
rect 10654 19760 13726 19816
rect 13782 19760 13787 19816
rect 5533 19758 13787 19760
rect 5533 19755 5599 19758
rect 10593 19755 10659 19758
rect 13721 19755 13787 19758
rect 22093 19818 22159 19821
rect 28165 19818 28231 19821
rect 22093 19816 28231 19818
rect 22093 19760 22098 19816
rect 22154 19760 28170 19816
rect 28226 19760 28231 19816
rect 22093 19758 28231 19760
rect 22093 19755 22159 19758
rect 28165 19755 28231 19758
rect 68093 19818 68159 19821
rect 69200 19818 70000 19848
rect 68093 19816 70000 19818
rect 68093 19760 68098 19816
rect 68154 19760 70000 19816
rect 68093 19758 70000 19760
rect 68093 19755 68159 19758
rect 69200 19728 70000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 13445 19546 13511 19549
rect 18229 19546 18295 19549
rect 13445 19544 18295 19546
rect 13445 19488 13450 19544
rect 13506 19488 18234 19544
rect 18290 19488 18295 19544
rect 13445 19486 18295 19488
rect 13445 19483 13511 19486
rect 18229 19483 18295 19486
rect 20437 19546 20503 19549
rect 26509 19546 26575 19549
rect 20437 19544 26575 19546
rect 20437 19488 20442 19544
rect 20498 19488 26514 19544
rect 26570 19488 26575 19544
rect 20437 19486 26575 19488
rect 20437 19483 20503 19486
rect 26509 19483 26575 19486
rect 6637 19410 6703 19413
rect 8937 19410 9003 19413
rect 6637 19408 9003 19410
rect 6637 19352 6642 19408
rect 6698 19352 8942 19408
rect 8998 19352 9003 19408
rect 6637 19350 9003 19352
rect 6637 19347 6703 19350
rect 8937 19347 9003 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 18689 19002 18755 19005
rect 20110 19002 20116 19004
rect 13172 19000 20116 19002
rect 13172 18944 18694 19000
rect 18750 18944 20116 19000
rect 13172 18942 20116 18944
rect 2589 18866 2655 18869
rect 12617 18866 12683 18869
rect 2589 18864 12683 18866
rect 2589 18808 2594 18864
rect 2650 18808 12622 18864
rect 12678 18808 12683 18864
rect 2589 18806 12683 18808
rect 2589 18803 2655 18806
rect 12617 18803 12683 18806
rect 0 18640 800 18760
rect 5441 18730 5507 18733
rect 13172 18730 13232 18942
rect 18689 18939 18755 18942
rect 20110 18940 20116 18942
rect 20180 18940 20186 19004
rect 13302 18804 13308 18868
rect 13372 18866 13378 18868
rect 23381 18866 23447 18869
rect 13372 18864 23447 18866
rect 13372 18808 23386 18864
rect 23442 18808 23447 18864
rect 13372 18806 23447 18808
rect 13372 18804 13378 18806
rect 23381 18803 23447 18806
rect 5441 18728 13232 18730
rect 5441 18672 5446 18728
rect 5502 18672 13232 18728
rect 5441 18670 13232 18672
rect 5441 18667 5507 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 68093 18458 68159 18461
rect 69200 18458 70000 18488
rect 68093 18456 70000 18458
rect 68093 18400 68098 18456
rect 68154 18400 70000 18456
rect 68093 18398 70000 18400
rect 68093 18395 68159 18398
rect 69200 18368 70000 18398
rect 22461 18186 22527 18189
rect 23197 18186 23263 18189
rect 25773 18186 25839 18189
rect 22461 18184 25839 18186
rect 22461 18128 22466 18184
rect 22522 18128 23202 18184
rect 23258 18128 25778 18184
rect 25834 18128 25839 18184
rect 22461 18126 25839 18128
rect 22461 18123 22527 18126
rect 23197 18123 23263 18126
rect 25773 18123 25839 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 14774 17716 14780 17780
rect 14844 17778 14850 17780
rect 20529 17778 20595 17781
rect 14844 17776 20595 17778
rect 14844 17720 20534 17776
rect 20590 17720 20595 17776
rect 14844 17718 20595 17720
rect 14844 17716 14850 17718
rect 20529 17715 20595 17718
rect 29085 17778 29151 17781
rect 30833 17778 30899 17781
rect 29085 17776 30899 17778
rect 29085 17720 29090 17776
rect 29146 17720 30838 17776
rect 30894 17720 30899 17776
rect 29085 17718 30899 17720
rect 29085 17715 29151 17718
rect 30833 17715 30899 17718
rect 21909 17642 21975 17645
rect 29545 17642 29611 17645
rect 21909 17640 29611 17642
rect 21909 17584 21914 17640
rect 21970 17584 29550 17640
rect 29606 17584 29611 17640
rect 21909 17582 29611 17584
rect 21909 17579 21975 17582
rect 29545 17579 29611 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 2497 17370 2563 17373
rect 18965 17370 19031 17373
rect 2497 17368 19031 17370
rect 2497 17312 2502 17368
rect 2558 17312 18970 17368
rect 19026 17312 19031 17368
rect 2497 17310 19031 17312
rect 2497 17307 2563 17310
rect 18965 17307 19031 17310
rect 0 17144 800 17264
rect 5901 17234 5967 17237
rect 12617 17234 12683 17237
rect 5901 17232 12683 17234
rect 5901 17176 5906 17232
rect 5962 17176 12622 17232
rect 12678 17176 12683 17232
rect 5901 17174 12683 17176
rect 5901 17171 5967 17174
rect 12617 17171 12683 17174
rect 19241 17234 19307 17237
rect 19374 17234 19380 17236
rect 19241 17232 19380 17234
rect 19241 17176 19246 17232
rect 19302 17176 19380 17232
rect 19241 17174 19380 17176
rect 19241 17171 19307 17174
rect 19374 17172 19380 17174
rect 19444 17234 19450 17236
rect 19977 17234 20043 17237
rect 19444 17232 20043 17234
rect 19444 17176 19982 17232
rect 20038 17176 20043 17232
rect 19444 17174 20043 17176
rect 19444 17172 19450 17174
rect 19977 17171 20043 17174
rect 67633 17098 67699 17101
rect 69200 17098 70000 17128
rect 67633 17096 70000 17098
rect 67633 17040 67638 17096
rect 67694 17040 70000 17096
rect 67633 17038 70000 17040
rect 67633 17035 67699 17038
rect 69200 17008 70000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 17902 16628 17908 16692
rect 17972 16690 17978 16692
rect 18689 16690 18755 16693
rect 17972 16688 18755 16690
rect 17972 16632 18694 16688
rect 18750 16632 18755 16688
rect 17972 16630 18755 16632
rect 17972 16628 17978 16630
rect 18689 16627 18755 16630
rect 29453 16690 29519 16693
rect 30649 16690 30715 16693
rect 32305 16690 32371 16693
rect 29453 16688 32371 16690
rect 29453 16632 29458 16688
rect 29514 16632 30654 16688
rect 30710 16632 32310 16688
rect 32366 16632 32371 16688
rect 29453 16630 32371 16632
rect 29453 16627 29519 16630
rect 30649 16627 30715 16630
rect 32305 16627 32371 16630
rect 20529 16554 20595 16557
rect 22185 16554 22251 16557
rect 20529 16552 22251 16554
rect 20529 16496 20534 16552
rect 20590 16496 22190 16552
rect 22246 16496 22251 16552
rect 20529 16494 22251 16496
rect 20529 16491 20595 16494
rect 22185 16491 22251 16494
rect 29821 16554 29887 16557
rect 36261 16554 36327 16557
rect 29821 16552 36327 16554
rect 29821 16496 29826 16552
rect 29882 16496 36266 16552
rect 36322 16496 36327 16552
rect 29821 16494 36327 16496
rect 29821 16491 29887 16494
rect 36261 16491 36327 16494
rect 7373 16420 7439 16421
rect 7373 16418 7420 16420
rect 7328 16416 7420 16418
rect 7328 16360 7378 16416
rect 7328 16358 7420 16360
rect 7373 16356 7420 16358
rect 7484 16356 7490 16420
rect 20989 16418 21055 16421
rect 25405 16418 25471 16421
rect 20989 16416 25471 16418
rect 20989 16360 20994 16416
rect 21050 16360 25410 16416
rect 25466 16360 25471 16416
rect 20989 16358 25471 16360
rect 7373 16355 7439 16356
rect 20989 16355 21055 16358
rect 25405 16355 25471 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 3785 16282 3851 16285
rect 9765 16282 9831 16285
rect 3785 16280 9831 16282
rect 3785 16224 3790 16280
rect 3846 16224 9770 16280
rect 9826 16224 9831 16280
rect 3785 16222 9831 16224
rect 3785 16219 3851 16222
rect 9765 16219 9831 16222
rect 20345 16146 20411 16149
rect 28073 16146 28139 16149
rect 20345 16144 28139 16146
rect 20345 16088 20350 16144
rect 20406 16088 28078 16144
rect 28134 16088 28139 16144
rect 20345 16086 28139 16088
rect 20345 16083 20411 16086
rect 28073 16083 28139 16086
rect 8385 16010 8451 16013
rect 21357 16010 21423 16013
rect 8385 16008 21423 16010
rect 8385 15952 8390 16008
rect 8446 15952 21362 16008
rect 21418 15952 21423 16008
rect 8385 15950 21423 15952
rect 8385 15947 8451 15950
rect 21357 15947 21423 15950
rect 20529 15876 20595 15877
rect 20478 15812 20484 15876
rect 20548 15874 20595 15876
rect 21541 15874 21607 15877
rect 32581 15874 32647 15877
rect 20548 15872 20640 15874
rect 20590 15816 20640 15872
rect 20548 15814 20640 15816
rect 21541 15872 32647 15874
rect 21541 15816 21546 15872
rect 21602 15816 32586 15872
rect 32642 15816 32647 15872
rect 21541 15814 32647 15816
rect 20548 15812 20595 15814
rect 20529 15811 20595 15812
rect 21541 15811 21607 15814
rect 32581 15811 32647 15814
rect 4210 15808 4526 15809
rect 0 15648 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 7649 15738 7715 15741
rect 20713 15738 20779 15741
rect 7649 15736 20779 15738
rect 7649 15680 7654 15736
rect 7710 15680 20718 15736
rect 20774 15680 20779 15736
rect 7649 15678 20779 15680
rect 7649 15675 7715 15678
rect 20713 15675 20779 15678
rect 22369 15738 22435 15741
rect 30741 15738 30807 15741
rect 22369 15736 30807 15738
rect 22369 15680 22374 15736
rect 22430 15680 30746 15736
rect 30802 15680 30807 15736
rect 22369 15678 30807 15680
rect 22369 15675 22435 15678
rect 30741 15675 30807 15678
rect 67633 15738 67699 15741
rect 69200 15738 70000 15768
rect 67633 15736 70000 15738
rect 67633 15680 67638 15736
rect 67694 15680 70000 15736
rect 67633 15678 70000 15680
rect 67633 15675 67699 15678
rect 69200 15648 70000 15678
rect 9489 15602 9555 15605
rect 20069 15602 20135 15605
rect 9489 15600 20135 15602
rect 9489 15544 9494 15600
rect 9550 15544 20074 15600
rect 20130 15544 20135 15600
rect 9489 15542 20135 15544
rect 9489 15539 9555 15542
rect 20069 15539 20135 15542
rect 13445 15466 13511 15469
rect 23381 15466 23447 15469
rect 13445 15464 23447 15466
rect 13445 15408 13450 15464
rect 13506 15408 23386 15464
rect 23442 15408 23447 15464
rect 13445 15406 23447 15408
rect 13445 15403 13511 15406
rect 23381 15403 23447 15406
rect 19977 15330 20043 15333
rect 22369 15330 22435 15333
rect 19977 15328 22435 15330
rect 19977 15272 19982 15328
rect 20038 15272 22374 15328
rect 22430 15272 22435 15328
rect 19977 15270 22435 15272
rect 19977 15267 20043 15270
rect 22369 15267 22435 15270
rect 23473 15330 23539 15333
rect 28625 15330 28691 15333
rect 33317 15330 33383 15333
rect 33777 15330 33843 15333
rect 23473 15328 33843 15330
rect 23473 15272 23478 15328
rect 23534 15272 28630 15328
rect 28686 15272 33322 15328
rect 33378 15272 33782 15328
rect 33838 15272 33843 15328
rect 23473 15270 33843 15272
rect 23473 15267 23539 15270
rect 28625 15267 28691 15270
rect 33317 15267 33383 15270
rect 33777 15267 33843 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 12934 15132 12940 15196
rect 13004 15194 13010 15196
rect 14273 15194 14339 15197
rect 13004 15192 14339 15194
rect 13004 15136 14278 15192
rect 14334 15136 14339 15192
rect 13004 15134 14339 15136
rect 13004 15132 13010 15134
rect 14273 15131 14339 15134
rect 20069 15194 20135 15197
rect 24393 15194 24459 15197
rect 20069 15192 24459 15194
rect 20069 15136 20074 15192
rect 20130 15136 24398 15192
rect 24454 15136 24459 15192
rect 20069 15134 24459 15136
rect 20069 15131 20135 15134
rect 24393 15131 24459 15134
rect 20161 14922 20227 14925
rect 24761 14922 24827 14925
rect 20161 14920 24827 14922
rect 20161 14864 20166 14920
rect 20222 14864 24766 14920
rect 24822 14864 24827 14920
rect 20161 14862 24827 14864
rect 20161 14859 20227 14862
rect 24761 14859 24827 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 12985 14378 13051 14381
rect 25221 14378 25287 14381
rect 12985 14376 25287 14378
rect 12985 14320 12990 14376
rect 13046 14320 25226 14376
rect 25282 14320 25287 14376
rect 12985 14318 25287 14320
rect 12985 14315 13051 14318
rect 25221 14315 25287 14318
rect 38837 14378 38903 14381
rect 40493 14378 40559 14381
rect 38837 14376 40559 14378
rect 38837 14320 38842 14376
rect 38898 14320 40498 14376
rect 40554 14320 40559 14376
rect 38837 14318 40559 14320
rect 38837 14315 38903 14318
rect 40493 14315 40559 14318
rect 68093 14378 68159 14381
rect 69200 14378 70000 14408
rect 68093 14376 70000 14378
rect 68093 14320 68098 14376
rect 68154 14320 70000 14376
rect 68093 14318 70000 14320
rect 68093 14315 68159 14318
rect 69200 14288 70000 14318
rect 0 14152 800 14272
rect 20069 14244 20135 14245
rect 20069 14242 20116 14244
rect 20024 14240 20116 14242
rect 20024 14184 20074 14240
rect 20024 14182 20116 14184
rect 20069 14180 20116 14182
rect 20180 14180 20186 14244
rect 20529 14242 20595 14245
rect 28257 14242 28323 14245
rect 20529 14240 28323 14242
rect 20529 14184 20534 14240
rect 20590 14184 28262 14240
rect 28318 14184 28323 14240
rect 20529 14182 28323 14184
rect 20069 14179 20135 14180
rect 20529 14179 20595 14182
rect 28257 14179 28323 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 20161 14106 20227 14109
rect 25497 14106 25563 14109
rect 20161 14104 25563 14106
rect 20161 14048 20166 14104
rect 20222 14048 25502 14104
rect 25558 14048 25563 14104
rect 20161 14046 25563 14048
rect 20161 14043 20227 14046
rect 25497 14043 25563 14046
rect 15837 13972 15903 13973
rect 15837 13968 15884 13972
rect 15948 13970 15954 13972
rect 17585 13970 17651 13973
rect 24342 13970 24348 13972
rect 15837 13912 15842 13968
rect 15837 13908 15884 13912
rect 15948 13910 15994 13970
rect 17585 13968 24348 13970
rect 17585 13912 17590 13968
rect 17646 13912 24348 13968
rect 17585 13910 24348 13912
rect 15948 13908 15954 13910
rect 15837 13907 15903 13908
rect 17585 13907 17651 13910
rect 24342 13908 24348 13910
rect 24412 13908 24418 13972
rect 10869 13834 10935 13837
rect 22093 13834 22159 13837
rect 10869 13832 22159 13834
rect 10869 13776 10874 13832
rect 10930 13776 22098 13832
rect 22154 13776 22159 13832
rect 10869 13774 22159 13776
rect 10869 13771 10935 13774
rect 22093 13771 22159 13774
rect 12198 13636 12204 13700
rect 12268 13698 12274 13700
rect 12801 13698 12867 13701
rect 12268 13696 12867 13698
rect 12268 13640 12806 13696
rect 12862 13640 12867 13696
rect 12268 13638 12867 13640
rect 12268 13636 12274 13638
rect 12801 13635 12867 13638
rect 14365 13700 14431 13701
rect 14365 13696 14412 13700
rect 14476 13698 14482 13700
rect 14641 13698 14707 13701
rect 14774 13698 14780 13700
rect 14365 13640 14370 13696
rect 14365 13636 14412 13640
rect 14476 13638 14522 13698
rect 14641 13696 14780 13698
rect 14641 13640 14646 13696
rect 14702 13640 14780 13696
rect 14641 13638 14780 13640
rect 14476 13636 14482 13638
rect 14365 13635 14431 13636
rect 14641 13635 14707 13638
rect 14774 13636 14780 13638
rect 14844 13636 14850 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 12893 13426 12959 13429
rect 18873 13426 18939 13429
rect 12893 13424 18939 13426
rect 12893 13368 12898 13424
rect 12954 13368 18878 13424
rect 18934 13368 18939 13424
rect 12893 13366 18939 13368
rect 12893 13363 12959 13366
rect 18873 13363 18939 13366
rect 21081 13426 21147 13429
rect 27521 13426 27587 13429
rect 21081 13424 27587 13426
rect 21081 13368 21086 13424
rect 21142 13368 27526 13424
rect 27582 13368 27587 13424
rect 21081 13366 27587 13368
rect 21081 13363 21147 13366
rect 27521 13363 27587 13366
rect 30005 13290 30071 13293
rect 36077 13290 36143 13293
rect 30005 13288 36143 13290
rect 30005 13232 30010 13288
rect 30066 13232 36082 13288
rect 36138 13232 36143 13288
rect 30005 13230 36143 13232
rect 30005 13227 30071 13230
rect 36077 13227 36143 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 17125 13020 17191 13021
rect 17125 13018 17172 13020
rect 17080 13016 17172 13018
rect 17236 13018 17242 13020
rect 17861 13018 17927 13021
rect 17236 13016 17927 13018
rect 17080 12960 17130 13016
rect 17236 12960 17866 13016
rect 17922 12960 17927 13016
rect 17080 12958 17172 12960
rect 17125 12956 17172 12958
rect 17236 12958 17927 12960
rect 17236 12956 17242 12958
rect 17125 12955 17191 12956
rect 17861 12955 17927 12958
rect 68093 13018 68159 13021
rect 69200 13018 70000 13048
rect 68093 13016 70000 13018
rect 68093 12960 68098 13016
rect 68154 12960 70000 13016
rect 68093 12958 70000 12960
rect 68093 12955 68159 12958
rect 69200 12928 70000 12958
rect 15377 12882 15443 12885
rect 21725 12882 21791 12885
rect 15377 12880 21791 12882
rect 15377 12824 15382 12880
rect 15438 12824 21730 12880
rect 21786 12824 21791 12880
rect 15377 12822 21791 12824
rect 15377 12819 15443 12822
rect 21725 12819 21791 12822
rect 0 12656 800 12776
rect 12341 12746 12407 12749
rect 28993 12746 29059 12749
rect 12341 12744 29059 12746
rect 12341 12688 12346 12744
rect 12402 12688 28998 12744
rect 29054 12688 29059 12744
rect 12341 12686 29059 12688
rect 12341 12683 12407 12686
rect 28993 12683 29059 12686
rect 14457 12610 14523 12613
rect 27429 12610 27495 12613
rect 14457 12608 27495 12610
rect 14457 12552 14462 12608
rect 14518 12552 27434 12608
rect 27490 12552 27495 12608
rect 14457 12550 27495 12552
rect 14457 12547 14523 12550
rect 27429 12547 27495 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 13077 12474 13143 12477
rect 30281 12474 30347 12477
rect 13077 12472 30347 12474
rect 13077 12416 13082 12472
rect 13138 12416 30286 12472
rect 30342 12416 30347 12472
rect 13077 12414 30347 12416
rect 13077 12411 13143 12414
rect 30281 12411 30347 12414
rect 13169 12338 13235 12341
rect 13302 12338 13308 12340
rect 13169 12336 13308 12338
rect 13169 12280 13174 12336
rect 13230 12280 13308 12336
rect 13169 12278 13308 12280
rect 13169 12275 13235 12278
rect 13302 12276 13308 12278
rect 13372 12276 13378 12340
rect 16573 12202 16639 12205
rect 25589 12202 25655 12205
rect 16573 12200 25655 12202
rect 16573 12144 16578 12200
rect 16634 12144 25594 12200
rect 25650 12144 25655 12200
rect 16573 12142 25655 12144
rect 16573 12139 16639 12142
rect 25589 12139 25655 12142
rect 19425 12068 19491 12069
rect 19374 12066 19380 12068
rect 19334 12006 19380 12066
rect 19444 12064 19491 12068
rect 19486 12008 19491 12064
rect 19374 12004 19380 12006
rect 19444 12004 19491 12008
rect 19425 12003 19491 12004
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 24342 11868 24348 11932
rect 24412 11930 24418 11932
rect 24577 11930 24643 11933
rect 24412 11928 24643 11930
rect 24412 11872 24582 11928
rect 24638 11872 24643 11928
rect 24412 11870 24643 11872
rect 24412 11868 24418 11870
rect 24577 11867 24643 11870
rect 19701 11794 19767 11797
rect 22277 11794 22343 11797
rect 19701 11792 22343 11794
rect 19701 11736 19706 11792
rect 19762 11736 22282 11792
rect 22338 11736 22343 11792
rect 19701 11734 22343 11736
rect 19701 11731 19767 11734
rect 22277 11731 22343 11734
rect 9581 11658 9647 11661
rect 25957 11658 26023 11661
rect 9581 11656 26023 11658
rect 9581 11600 9586 11656
rect 9642 11600 25962 11656
rect 26018 11600 26023 11656
rect 9581 11598 26023 11600
rect 9581 11595 9647 11598
rect 25957 11595 26023 11598
rect 67633 11658 67699 11661
rect 69200 11658 70000 11688
rect 67633 11656 70000 11658
rect 67633 11600 67638 11656
rect 67694 11600 70000 11656
rect 67633 11598 70000 11600
rect 67633 11595 67699 11598
rect 69200 11568 70000 11598
rect 10593 11522 10659 11525
rect 25037 11522 25103 11525
rect 10593 11520 25103 11522
rect 10593 11464 10598 11520
rect 10654 11464 25042 11520
rect 25098 11464 25103 11520
rect 10593 11462 25103 11464
rect 10593 11459 10659 11462
rect 25037 11459 25103 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 19793 11386 19859 11389
rect 24117 11386 24183 11389
rect 19793 11384 24183 11386
rect 19793 11328 19798 11384
rect 19854 11328 24122 11384
rect 24178 11328 24183 11384
rect 19793 11326 24183 11328
rect 19793 11323 19859 11326
rect 24117 11323 24183 11326
rect 31385 11386 31451 11389
rect 34421 11386 34487 11389
rect 31385 11384 34487 11386
rect 31385 11328 31390 11384
rect 31446 11328 34426 11384
rect 34482 11328 34487 11384
rect 31385 11326 34487 11328
rect 31385 11323 31451 11326
rect 34421 11323 34487 11326
rect 0 11160 800 11280
rect 16481 11250 16547 11253
rect 29637 11250 29703 11253
rect 16481 11248 29703 11250
rect 16481 11192 16486 11248
rect 16542 11192 29642 11248
rect 29698 11192 29703 11248
rect 16481 11190 29703 11192
rect 16481 11187 16547 11190
rect 29637 11187 29703 11190
rect 31661 11250 31727 11253
rect 37549 11250 37615 11253
rect 31661 11248 37615 11250
rect 31661 11192 31666 11248
rect 31722 11192 37554 11248
rect 37610 11192 37615 11248
rect 31661 11190 37615 11192
rect 31661 11187 31727 11190
rect 37549 11187 37615 11190
rect 11053 11116 11119 11117
rect 11053 11114 11100 11116
rect 11008 11112 11100 11114
rect 11008 11056 11058 11112
rect 11008 11054 11100 11056
rect 11053 11052 11100 11054
rect 11164 11052 11170 11116
rect 19977 11114 20043 11117
rect 20110 11114 20116 11116
rect 19977 11112 20116 11114
rect 19977 11056 19982 11112
rect 20038 11056 20116 11112
rect 19977 11054 20116 11056
rect 11053 11051 11119 11052
rect 19977 11051 20043 11054
rect 20110 11052 20116 11054
rect 20180 11052 20186 11116
rect 17309 10978 17375 10981
rect 17902 10978 17908 10980
rect 17309 10976 17908 10978
rect 17309 10920 17314 10976
rect 17370 10920 17908 10976
rect 17309 10918 17908 10920
rect 17309 10915 17375 10918
rect 17902 10916 17908 10918
rect 17972 10916 17978 10980
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 5625 10706 5691 10709
rect 14365 10706 14431 10709
rect 5625 10704 14431 10706
rect 5625 10648 5630 10704
rect 5686 10648 14370 10704
rect 14426 10648 14431 10704
rect 5625 10646 14431 10648
rect 5625 10643 5691 10646
rect 14365 10643 14431 10646
rect 17217 10706 17283 10709
rect 30005 10706 30071 10709
rect 17217 10704 30071 10706
rect 17217 10648 17222 10704
rect 17278 10648 30010 10704
rect 30066 10648 30071 10704
rect 17217 10646 30071 10648
rect 17217 10643 17283 10646
rect 30005 10643 30071 10646
rect 12065 10570 12131 10573
rect 29545 10570 29611 10573
rect 12065 10568 29611 10570
rect 12065 10512 12070 10568
rect 12126 10512 29550 10568
rect 29606 10512 29611 10568
rect 12065 10510 29611 10512
rect 12065 10507 12131 10510
rect 29545 10507 29611 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 67633 10298 67699 10301
rect 69200 10298 70000 10328
rect 67633 10296 70000 10298
rect 67633 10240 67638 10296
rect 67694 10240 70000 10296
rect 67633 10238 70000 10240
rect 67633 10235 67699 10238
rect 69200 10208 70000 10238
rect 19570 9824 19886 9825
rect 0 9664 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 15142 9284 15148 9348
rect 15212 9346 15218 9348
rect 19885 9346 19951 9349
rect 20529 9346 20595 9349
rect 15212 9344 20595 9346
rect 15212 9288 19890 9344
rect 19946 9288 20534 9344
rect 20590 9288 20595 9344
rect 15212 9286 20595 9288
rect 15212 9284 15218 9286
rect 19885 9283 19951 9286
rect 20529 9283 20595 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 22921 8938 22987 8941
rect 32489 8938 32555 8941
rect 22921 8936 32555 8938
rect 22921 8880 22926 8936
rect 22982 8880 32494 8936
rect 32550 8880 32555 8936
rect 22921 8878 32555 8880
rect 22921 8875 22987 8878
rect 32489 8875 32555 8878
rect 68093 8938 68159 8941
rect 69200 8938 70000 8968
rect 68093 8936 70000 8938
rect 68093 8880 68098 8936
rect 68154 8880 70000 8936
rect 68093 8878 70000 8880
rect 68093 8875 68159 8878
rect 69200 8848 70000 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 7649 8396 7715 8397
rect 7598 8394 7604 8396
rect 7558 8334 7604 8394
rect 7668 8392 7715 8396
rect 7710 8336 7715 8392
rect 7598 8332 7604 8334
rect 7668 8332 7715 8336
rect 7649 8331 7715 8332
rect 0 8168 800 8288
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 11094 7788 11100 7852
rect 11164 7850 11170 7852
rect 21449 7850 21515 7853
rect 11164 7848 21515 7850
rect 11164 7792 21454 7848
rect 21510 7792 21515 7848
rect 11164 7790 21515 7792
rect 11164 7788 11170 7790
rect 21449 7787 21515 7790
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 8293 7578 8359 7581
rect 11053 7578 11119 7581
rect 8293 7576 11119 7578
rect 8293 7520 8298 7576
rect 8354 7520 11058 7576
rect 11114 7520 11119 7576
rect 8293 7518 11119 7520
rect 8293 7515 8359 7518
rect 11053 7515 11119 7518
rect 68093 7578 68159 7581
rect 69200 7578 70000 7608
rect 68093 7576 70000 7578
rect 68093 7520 68098 7576
rect 68154 7520 70000 7576
rect 68093 7518 70000 7520
rect 68093 7515 68159 7518
rect 69200 7488 70000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 10961 6898 11027 6901
rect 14917 6898 14983 6901
rect 10961 6896 14983 6898
rect 10961 6840 10966 6896
rect 11022 6840 14922 6896
rect 14978 6840 14983 6896
rect 10961 6838 14983 6840
rect 10961 6835 11027 6838
rect 14917 6835 14983 6838
rect 0 6672 800 6792
rect 10685 6762 10751 6765
rect 12525 6762 12591 6765
rect 10685 6760 12591 6762
rect 10685 6704 10690 6760
rect 10746 6704 12530 6760
rect 12586 6704 12591 6760
rect 10685 6702 12591 6704
rect 10685 6699 10751 6702
rect 12525 6699 12591 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 28441 6354 28507 6357
rect 32673 6354 32739 6357
rect 28441 6352 32739 6354
rect 28441 6296 28446 6352
rect 28502 6296 32678 6352
rect 32734 6296 32739 6352
rect 28441 6294 32739 6296
rect 28441 6291 28507 6294
rect 32673 6291 32739 6294
rect 6126 6156 6132 6220
rect 6196 6218 6202 6220
rect 20069 6218 20135 6221
rect 20989 6218 21055 6221
rect 6196 6216 21055 6218
rect 6196 6160 20074 6216
rect 20130 6160 20994 6216
rect 21050 6160 21055 6216
rect 6196 6158 21055 6160
rect 6196 6156 6202 6158
rect 20069 6155 20135 6158
rect 20989 6155 21055 6158
rect 67633 6218 67699 6221
rect 69200 6218 70000 6248
rect 67633 6216 70000 6218
rect 67633 6160 67638 6216
rect 67694 6160 70000 6216
rect 67633 6158 70000 6160
rect 67633 6155 67699 6158
rect 69200 6128 70000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 8293 5810 8359 5813
rect 17585 5810 17651 5813
rect 8293 5808 17651 5810
rect 8293 5752 8298 5808
rect 8354 5752 17590 5808
rect 17646 5752 17651 5808
rect 8293 5750 17651 5752
rect 8293 5747 8359 5750
rect 17585 5747 17651 5750
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 5176 800 5296
rect 9305 5266 9371 5269
rect 17677 5266 17743 5269
rect 9305 5264 17743 5266
rect 9305 5208 9310 5264
rect 9366 5208 17682 5264
rect 17738 5208 17743 5264
rect 9305 5206 17743 5208
rect 9305 5203 9371 5206
rect 17677 5203 17743 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 10501 4858 10567 4861
rect 12341 4858 12407 4861
rect 10501 4856 12407 4858
rect 10501 4800 10506 4856
rect 10562 4800 12346 4856
rect 12402 4800 12407 4856
rect 10501 4798 12407 4800
rect 10501 4795 10567 4798
rect 12341 4795 12407 4798
rect 67633 4858 67699 4861
rect 69200 4858 70000 4888
rect 67633 4856 70000 4858
rect 67633 4800 67638 4856
rect 67694 4800 70000 4856
rect 67633 4798 70000 4800
rect 67633 4795 67699 4798
rect 69200 4768 70000 4798
rect 4705 4722 4771 4725
rect 11605 4722 11671 4725
rect 4705 4720 11671 4722
rect 4705 4664 4710 4720
rect 4766 4664 11610 4720
rect 11666 4664 11671 4720
rect 4705 4662 11671 4664
rect 4705 4659 4771 4662
rect 11605 4659 11671 4662
rect 11973 4722 12039 4725
rect 13169 4722 13235 4725
rect 11973 4720 13235 4722
rect 11973 4664 11978 4720
rect 12034 4664 13174 4720
rect 13230 4664 13235 4720
rect 11973 4662 13235 4664
rect 11973 4659 12039 4662
rect 13169 4659 13235 4662
rect 10409 4586 10475 4589
rect 14917 4586 14983 4589
rect 10409 4584 14983 4586
rect 10409 4528 10414 4584
rect 10470 4528 14922 4584
rect 14978 4528 14983 4584
rect 10409 4526 14983 4528
rect 10409 4523 10475 4526
rect 14917 4523 14983 4526
rect 8937 4450 9003 4453
rect 13813 4450 13879 4453
rect 8937 4448 13879 4450
rect 8937 4392 8942 4448
rect 8998 4392 13818 4448
rect 13874 4392 13879 4448
rect 8937 4390 13879 4392
rect 8937 4387 9003 4390
rect 13813 4387 13879 4390
rect 13997 4450 14063 4453
rect 18229 4450 18295 4453
rect 13997 4448 18295 4450
rect 13997 4392 14002 4448
rect 14058 4392 18234 4448
rect 18290 4392 18295 4448
rect 13997 4390 18295 4392
rect 13997 4387 14063 4390
rect 18229 4387 18295 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 3417 4314 3483 4317
rect 8845 4314 8911 4317
rect 3417 4312 8911 4314
rect 3417 4256 3422 4312
rect 3478 4256 8850 4312
rect 8906 4256 8911 4312
rect 3417 4254 8911 4256
rect 3417 4251 3483 4254
rect 8845 4251 8911 4254
rect 9673 4314 9739 4317
rect 15101 4314 15167 4317
rect 9673 4312 15167 4314
rect 9673 4256 9678 4312
rect 9734 4256 15106 4312
rect 15162 4256 15167 4312
rect 9673 4254 15167 4256
rect 9673 4251 9739 4254
rect 15101 4251 15167 4254
rect 9622 4116 9628 4180
rect 9692 4178 9698 4180
rect 10501 4178 10567 4181
rect 16573 4178 16639 4181
rect 9692 4176 10567 4178
rect 9692 4120 10506 4176
rect 10562 4120 10567 4176
rect 9692 4118 10567 4120
rect 9692 4116 9698 4118
rect 10501 4115 10567 4118
rect 16438 4176 16639 4178
rect 16438 4120 16578 4176
rect 16634 4120 16639 4176
rect 16438 4118 16639 4120
rect 2129 4042 2195 4045
rect 5809 4042 5875 4045
rect 10133 4042 10199 4045
rect 11789 4042 11855 4045
rect 16438 4042 16498 4118
rect 16573 4115 16639 4118
rect 2129 4040 5642 4042
rect 2129 3984 2134 4040
rect 2190 3984 5642 4040
rect 2129 3982 5642 3984
rect 2129 3979 2195 3982
rect 5582 3906 5642 3982
rect 5809 4040 11714 4042
rect 5809 3984 5814 4040
rect 5870 3984 10138 4040
rect 10194 3984 11714 4040
rect 5809 3982 11714 3984
rect 5809 3979 5875 3982
rect 10133 3979 10199 3982
rect 7414 3906 7420 3908
rect 5582 3846 7420 3906
rect 7414 3844 7420 3846
rect 7484 3906 7490 3908
rect 10593 3906 10659 3909
rect 7484 3904 10659 3906
rect 7484 3848 10598 3904
rect 10654 3848 10659 3904
rect 7484 3846 10659 3848
rect 11654 3906 11714 3982
rect 11789 4040 16498 4042
rect 11789 3984 11794 4040
rect 11850 3984 16498 4040
rect 11789 3982 16498 3984
rect 11789 3979 11855 3982
rect 12709 3906 12775 3909
rect 11654 3904 12775 3906
rect 11654 3848 12714 3904
rect 12770 3848 12775 3904
rect 11654 3846 12775 3848
rect 7484 3844 7490 3846
rect 10593 3843 10659 3846
rect 12709 3843 12775 3846
rect 13261 3906 13327 3909
rect 13905 3906 13971 3909
rect 20897 3906 20963 3909
rect 13261 3904 20963 3906
rect 13261 3848 13266 3904
rect 13322 3848 13910 3904
rect 13966 3848 20902 3904
rect 20958 3848 20963 3904
rect 13261 3846 20963 3848
rect 13261 3843 13327 3846
rect 13905 3843 13971 3846
rect 20897 3843 20963 3846
rect 4210 3840 4526 3841
rect 0 3680 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 6729 3770 6795 3773
rect 8937 3770 9003 3773
rect 6729 3768 9003 3770
rect 6729 3712 6734 3768
rect 6790 3712 8942 3768
rect 8998 3712 9003 3768
rect 6729 3710 9003 3712
rect 6729 3707 6795 3710
rect 8937 3707 9003 3710
rect 10685 3770 10751 3773
rect 19885 3770 19951 3773
rect 10685 3768 19951 3770
rect 10685 3712 10690 3768
rect 10746 3712 19890 3768
rect 19946 3712 19951 3768
rect 10685 3710 19951 3712
rect 10685 3707 10751 3710
rect 19885 3707 19951 3710
rect 7557 3636 7623 3637
rect 7557 3634 7604 3636
rect 7512 3632 7604 3634
rect 7512 3576 7562 3632
rect 7512 3574 7604 3576
rect 7557 3572 7604 3574
rect 7668 3572 7674 3636
rect 10041 3634 10107 3637
rect 13077 3634 13143 3637
rect 10041 3632 13143 3634
rect 10041 3576 10046 3632
rect 10102 3576 13082 3632
rect 13138 3576 13143 3632
rect 10041 3574 13143 3576
rect 7557 3571 7623 3572
rect 10041 3571 10107 3574
rect 13077 3571 13143 3574
rect 13721 3634 13787 3637
rect 16113 3634 16179 3637
rect 13721 3632 16179 3634
rect 13721 3576 13726 3632
rect 13782 3576 16118 3632
rect 16174 3576 16179 3632
rect 13721 3574 16179 3576
rect 13721 3571 13787 3574
rect 16113 3571 16179 3574
rect 2957 3498 3023 3501
rect 3877 3498 3943 3501
rect 9121 3498 9187 3501
rect 2957 3496 9187 3498
rect 2957 3440 2962 3496
rect 3018 3440 3882 3496
rect 3938 3440 9126 3496
rect 9182 3440 9187 3496
rect 2957 3438 9187 3440
rect 2957 3435 3023 3438
rect 3877 3435 3943 3438
rect 9121 3435 9187 3438
rect 10869 3498 10935 3501
rect 20478 3498 20484 3500
rect 10869 3496 20484 3498
rect 10869 3440 10874 3496
rect 10930 3440 20484 3496
rect 10869 3438 20484 3440
rect 10869 3435 10935 3438
rect 20478 3436 20484 3438
rect 20548 3436 20554 3500
rect 68093 3498 68159 3501
rect 69200 3498 70000 3528
rect 68093 3496 70000 3498
rect 68093 3440 68098 3496
rect 68154 3440 70000 3496
rect 68093 3438 70000 3440
rect 68093 3435 68159 3438
rect 69200 3408 70000 3438
rect 8845 3362 8911 3365
rect 14641 3362 14707 3365
rect 15142 3362 15148 3364
rect 8845 3360 15148 3362
rect 8845 3304 8850 3360
rect 8906 3304 14646 3360
rect 14702 3304 15148 3360
rect 8845 3302 15148 3304
rect 8845 3299 8911 3302
rect 14641 3299 14707 3302
rect 15142 3300 15148 3302
rect 15212 3300 15218 3364
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 6821 3226 6887 3229
rect 14365 3226 14431 3229
rect 6821 3224 14431 3226
rect 6821 3168 6826 3224
rect 6882 3168 14370 3224
rect 14426 3168 14431 3224
rect 6821 3166 14431 3168
rect 6821 3163 6887 3166
rect 14365 3163 14431 3166
rect 57881 3226 57947 3229
rect 60457 3226 60523 3229
rect 57881 3224 60523 3226
rect 57881 3168 57886 3224
rect 57942 3168 60462 3224
rect 60518 3168 60523 3224
rect 57881 3166 60523 3168
rect 57881 3163 57947 3166
rect 60457 3163 60523 3166
rect 4613 3090 4679 3093
rect 6126 3090 6132 3092
rect 4613 3088 6132 3090
rect 4613 3032 4618 3088
rect 4674 3032 6132 3088
rect 4613 3030 6132 3032
rect 4613 3027 4679 3030
rect 6126 3028 6132 3030
rect 6196 3028 6202 3092
rect 6269 3090 6335 3093
rect 10501 3090 10567 3093
rect 17166 3090 17172 3092
rect 6269 3088 10567 3090
rect 6269 3032 6274 3088
rect 6330 3032 10506 3088
rect 10562 3032 10567 3088
rect 6269 3030 10567 3032
rect 6269 3027 6335 3030
rect 10501 3027 10567 3030
rect 12390 3030 17172 3090
rect 10593 2954 10659 2957
rect 12390 2954 12450 3030
rect 17166 3028 17172 3030
rect 17236 3028 17242 3092
rect 10593 2952 12450 2954
rect 10593 2896 10598 2952
rect 10654 2896 12450 2952
rect 10593 2894 12450 2896
rect 13261 2954 13327 2957
rect 13445 2954 13511 2957
rect 14549 2954 14615 2957
rect 13261 2952 13370 2954
rect 13261 2896 13266 2952
rect 13322 2896 13370 2952
rect 10593 2891 10659 2894
rect 13261 2891 13370 2896
rect 13445 2952 14615 2954
rect 13445 2896 13450 2952
rect 13506 2896 14554 2952
rect 14610 2896 14615 2952
rect 13445 2894 14615 2896
rect 13445 2891 13511 2894
rect 14549 2891 14615 2894
rect 10409 2818 10475 2821
rect 10869 2818 10935 2821
rect 10409 2816 10935 2818
rect 10409 2760 10414 2816
rect 10470 2760 10874 2816
rect 10930 2760 10935 2816
rect 10409 2758 10935 2760
rect 13310 2818 13370 2891
rect 13445 2818 13511 2821
rect 13310 2816 13511 2818
rect 13310 2760 13450 2816
rect 13506 2760 13511 2816
rect 13310 2758 13511 2760
rect 10409 2755 10475 2758
rect 10869 2755 10935 2758
rect 13445 2755 13511 2758
rect 13813 2818 13879 2821
rect 17861 2818 17927 2821
rect 13813 2816 17927 2818
rect 13813 2760 13818 2816
rect 13874 2760 17866 2816
rect 17922 2760 17927 2816
rect 13813 2758 17927 2760
rect 13813 2755 13879 2758
rect 17861 2755 17927 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 11094 2620 11100 2684
rect 11164 2682 11170 2684
rect 11237 2682 11303 2685
rect 11164 2680 11303 2682
rect 11164 2624 11242 2680
rect 11298 2624 11303 2680
rect 11164 2622 11303 2624
rect 11164 2620 11170 2622
rect 11237 2619 11303 2622
rect 15009 2682 15075 2685
rect 19374 2682 19380 2684
rect 15009 2680 19380 2682
rect 15009 2624 15014 2680
rect 15070 2624 19380 2680
rect 15009 2622 19380 2624
rect 15009 2619 15075 2622
rect 19374 2620 19380 2622
rect 19444 2620 19450 2684
rect 15878 2484 15884 2548
rect 15948 2546 15954 2548
rect 17585 2546 17651 2549
rect 15948 2544 17651 2546
rect 15948 2488 17590 2544
rect 17646 2488 17651 2544
rect 15948 2486 17651 2488
rect 15948 2484 15954 2486
rect 17585 2483 17651 2486
rect 5257 2410 5323 2413
rect 18229 2410 18295 2413
rect 5257 2408 18295 2410
rect 5257 2352 5262 2408
rect 5318 2352 18234 2408
rect 18290 2352 18295 2408
rect 5257 2350 18295 2352
rect 5257 2347 5323 2350
rect 18229 2347 18295 2350
rect 0 2184 800 2304
rect 5165 2274 5231 2277
rect 15561 2274 15627 2277
rect 5165 2272 15627 2274
rect 5165 2216 5170 2272
rect 5226 2216 15566 2272
rect 15622 2216 15627 2272
rect 5165 2214 15627 2216
rect 5165 2211 5231 2214
rect 15561 2211 15627 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 3049 2138 3115 2141
rect 13169 2138 13235 2141
rect 3049 2136 13235 2138
rect 3049 2080 3054 2136
rect 3110 2080 13174 2136
rect 13230 2080 13235 2136
rect 3049 2078 13235 2080
rect 3049 2075 3115 2078
rect 13169 2075 13235 2078
rect 66989 2138 67055 2141
rect 69200 2138 70000 2168
rect 66989 2136 70000 2138
rect 66989 2080 66994 2136
rect 67050 2080 70000 2136
rect 66989 2078 70000 2080
rect 66989 2075 67055 2078
rect 69200 2048 70000 2078
rect 4061 2002 4127 2005
rect 13077 2002 13143 2005
rect 4061 2000 13143 2002
rect 4061 1944 4066 2000
rect 4122 1944 13082 2000
rect 13138 1944 13143 2000
rect 4061 1942 13143 1944
rect 4061 1939 4127 1942
rect 13077 1939 13143 1942
rect 1945 1866 2011 1869
rect 9622 1866 9628 1868
rect 1945 1864 9628 1866
rect 1945 1808 1950 1864
rect 2006 1808 9628 1864
rect 1945 1806 9628 1808
rect 1945 1803 2011 1806
rect 9622 1804 9628 1806
rect 9692 1804 9698 1868
rect 2405 1730 2471 1733
rect 12617 1730 12683 1733
rect 2405 1728 12683 1730
rect 2405 1672 2410 1728
rect 2466 1672 12622 1728
rect 12678 1672 12683 1728
rect 2405 1670 12683 1672
rect 2405 1667 2471 1670
rect 12617 1667 12683 1670
rect 9029 1594 9095 1597
rect 15878 1594 15884 1596
rect 9029 1592 15884 1594
rect 9029 1536 9034 1592
rect 9090 1536 15884 1592
rect 9029 1534 15884 1536
rect 9029 1531 9095 1534
rect 15878 1532 15884 1534
rect 15948 1532 15954 1596
rect 67541 778 67607 781
rect 69200 778 70000 808
rect 67541 776 70000 778
rect 67541 720 67546 776
rect 67602 720 70000 776
rect 67541 718 70000 720
rect 67541 715 67607 718
rect 69200 688 70000 718
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 12204 29336 12268 29340
rect 12204 29280 12218 29336
rect 12218 29280 12268 29336
rect 12204 29276 12268 29280
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 12940 27644 13004 27708
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19380 24032 19444 24036
rect 19380 23976 19394 24032
rect 19394 23976 19444 24032
rect 19380 23972 19444 23976
rect 20116 23972 20180 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 14412 23428 14476 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 17172 20708 17236 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 20116 18940 20180 19004
rect 13308 18804 13372 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 14780 17716 14844 17780
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 19380 17172 19444 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 17908 16628 17972 16692
rect 7420 16416 7484 16420
rect 7420 16360 7434 16416
rect 7434 16360 7484 16416
rect 7420 16356 7484 16360
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 20484 15872 20548 15876
rect 20484 15816 20534 15872
rect 20534 15816 20548 15872
rect 20484 15812 20548 15816
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 12940 15132 13004 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 20116 14240 20180 14244
rect 20116 14184 20130 14240
rect 20130 14184 20180 14240
rect 20116 14180 20180 14184
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 15884 13968 15948 13972
rect 15884 13912 15898 13968
rect 15898 13912 15948 13968
rect 15884 13908 15948 13912
rect 24348 13908 24412 13972
rect 12204 13636 12268 13700
rect 14412 13696 14476 13700
rect 14412 13640 14426 13696
rect 14426 13640 14476 13696
rect 14412 13636 14476 13640
rect 14780 13636 14844 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 17172 13016 17236 13020
rect 17172 12960 17186 13016
rect 17186 12960 17236 13016
rect 17172 12956 17236 12960
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 13308 12276 13372 12340
rect 19380 12064 19444 12068
rect 19380 12008 19430 12064
rect 19430 12008 19444 12064
rect 19380 12004 19444 12008
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 24348 11868 24412 11932
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 11100 11112 11164 11116
rect 11100 11056 11114 11112
rect 11114 11056 11164 11112
rect 11100 11052 11164 11056
rect 20116 11052 20180 11116
rect 17908 10916 17972 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 15148 9284 15212 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 7604 8392 7668 8396
rect 7604 8336 7654 8392
rect 7654 8336 7668 8392
rect 7604 8332 7668 8336
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 11100 7788 11164 7852
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 6132 6156 6196 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 9628 4116 9692 4180
rect 7420 3844 7484 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 7604 3632 7668 3636
rect 7604 3576 7618 3632
rect 7618 3576 7668 3632
rect 7604 3572 7668 3576
rect 20484 3436 20548 3500
rect 15148 3300 15212 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 6132 3028 6196 3092
rect 17172 3028 17236 3092
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 11100 2620 11164 2684
rect 19380 2620 19444 2684
rect 15884 2484 15948 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
rect 9628 1804 9692 1868
rect 15884 1532 15948 1596
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 12203 29340 12269 29341
rect 12203 29276 12204 29340
rect 12268 29276 12269 29340
rect 12203 29275 12269 29276
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 7419 16420 7485 16421
rect 7419 16356 7420 16420
rect 7484 16356 7485 16420
rect 7419 16355 7485 16356
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 6131 6220 6197 6221
rect 6131 6156 6132 6220
rect 6196 6156 6197 6220
rect 6131 6155 6197 6156
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 6134 3093 6194 6155
rect 7422 3909 7482 16355
rect 12206 13701 12266 29275
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 12939 27708 13005 27709
rect 12939 27644 12940 27708
rect 13004 27644 13005 27708
rect 12939 27643 13005 27644
rect 12942 15197 13002 27643
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19379 24036 19445 24037
rect 19379 23972 19380 24036
rect 19444 23972 19445 24036
rect 19379 23971 19445 23972
rect 14411 23492 14477 23493
rect 14411 23428 14412 23492
rect 14476 23428 14477 23492
rect 14411 23427 14477 23428
rect 13307 18868 13373 18869
rect 13307 18804 13308 18868
rect 13372 18804 13373 18868
rect 13307 18803 13373 18804
rect 12939 15196 13005 15197
rect 12939 15132 12940 15196
rect 13004 15132 13005 15196
rect 12939 15131 13005 15132
rect 12203 13700 12269 13701
rect 12203 13636 12204 13700
rect 12268 13636 12269 13700
rect 12203 13635 12269 13636
rect 13310 12341 13370 18803
rect 14414 13701 14474 23427
rect 17171 20772 17237 20773
rect 17171 20708 17172 20772
rect 17236 20708 17237 20772
rect 17171 20707 17237 20708
rect 14779 17780 14845 17781
rect 14779 17716 14780 17780
rect 14844 17716 14845 17780
rect 14779 17715 14845 17716
rect 14782 13701 14842 17715
rect 15883 13972 15949 13973
rect 15883 13908 15884 13972
rect 15948 13908 15949 13972
rect 15883 13907 15949 13908
rect 14411 13700 14477 13701
rect 14411 13636 14412 13700
rect 14476 13636 14477 13700
rect 14411 13635 14477 13636
rect 14779 13700 14845 13701
rect 14779 13636 14780 13700
rect 14844 13636 14845 13700
rect 14779 13635 14845 13636
rect 13307 12340 13373 12341
rect 13307 12276 13308 12340
rect 13372 12276 13373 12340
rect 13307 12275 13373 12276
rect 11099 11116 11165 11117
rect 11099 11052 11100 11116
rect 11164 11052 11165 11116
rect 11099 11051 11165 11052
rect 7603 8396 7669 8397
rect 7603 8332 7604 8396
rect 7668 8332 7669 8396
rect 7603 8331 7669 8332
rect 7419 3908 7485 3909
rect 7419 3844 7420 3908
rect 7484 3844 7485 3908
rect 7419 3843 7485 3844
rect 7606 3637 7666 8331
rect 11102 7853 11162 11051
rect 15147 9348 15213 9349
rect 15147 9284 15148 9348
rect 15212 9284 15213 9348
rect 15147 9283 15213 9284
rect 11099 7852 11165 7853
rect 11099 7788 11100 7852
rect 11164 7788 11165 7852
rect 11099 7787 11165 7788
rect 9627 4180 9693 4181
rect 9627 4116 9628 4180
rect 9692 4116 9693 4180
rect 9627 4115 9693 4116
rect 7603 3636 7669 3637
rect 7603 3572 7604 3636
rect 7668 3572 7669 3636
rect 7603 3571 7669 3572
rect 6131 3092 6197 3093
rect 6131 3028 6132 3092
rect 6196 3028 6197 3092
rect 6131 3027 6197 3028
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 9630 1869 9690 4115
rect 11102 2685 11162 7787
rect 15150 3365 15210 9283
rect 15147 3364 15213 3365
rect 15147 3300 15148 3364
rect 15212 3300 15213 3364
rect 15147 3299 15213 3300
rect 11099 2684 11165 2685
rect 11099 2620 11100 2684
rect 11164 2620 11165 2684
rect 11099 2619 11165 2620
rect 15886 2549 15946 13907
rect 17174 13021 17234 20707
rect 19382 17237 19442 23971
rect 19568 23968 19888 24992
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 20115 24036 20181 24037
rect 20115 23972 20116 24036
rect 20180 23972 20181 24036
rect 20115 23971 20181 23972
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 20118 19005 20178 23971
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 20115 19004 20181 19005
rect 20115 18940 20116 19004
rect 20180 18940 20181 19004
rect 20115 18939 20181 18940
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19379 17236 19445 17237
rect 19379 17172 19380 17236
rect 19444 17172 19445 17236
rect 19379 17171 19445 17172
rect 17907 16692 17973 16693
rect 17907 16628 17908 16692
rect 17972 16628 17973 16692
rect 17907 16627 17973 16628
rect 17171 13020 17237 13021
rect 17171 12956 17172 13020
rect 17236 12956 17237 13020
rect 17171 12955 17237 12956
rect 17174 3093 17234 12955
rect 17910 10981 17970 16627
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 20483 15876 20549 15877
rect 20483 15812 20484 15876
rect 20548 15812 20549 15876
rect 20483 15811 20549 15812
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 20115 14244 20181 14245
rect 20115 14180 20116 14244
rect 20180 14180 20181 14244
rect 20115 14179 20181 14180
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19379 12068 19445 12069
rect 19379 12004 19380 12068
rect 19444 12004 19445 12068
rect 19379 12003 19445 12004
rect 17907 10980 17973 10981
rect 17907 10916 17908 10980
rect 17972 10916 17973 10980
rect 17907 10915 17973 10916
rect 17171 3092 17237 3093
rect 17171 3028 17172 3092
rect 17236 3028 17237 3092
rect 17171 3027 17237 3028
rect 19382 2685 19442 12003
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 20118 11117 20178 14179
rect 20115 11116 20181 11117
rect 20115 11052 20116 11116
rect 20180 11052 20181 11116
rect 20115 11051 20181 11052
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 20486 3501 20546 15811
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 24347 13972 24413 13973
rect 24347 13908 24348 13972
rect 24412 13908 24413 13972
rect 24347 13907 24413 13908
rect 24350 11933 24410 13907
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 24347 11932 24413 11933
rect 24347 11868 24348 11932
rect 24412 11868 24413 11932
rect 24347 11867 24413 11868
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 20483 3500 20549 3501
rect 20483 3436 20484 3500
rect 20548 3436 20549 3500
rect 20483 3435 20549 3436
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19379 2684 19445 2685
rect 19379 2620 19380 2684
rect 19444 2620 19445 2684
rect 19379 2619 19445 2620
rect 15883 2548 15949 2549
rect 15883 2484 15884 2548
rect 15948 2484 15949 2548
rect 15883 2483 15949 2484
rect 9627 1868 9693 1869
rect 9627 1804 9628 1868
rect 9692 1804 9693 1868
rect 9627 1803 9693 1804
rect 15886 1597 15946 2483
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 57152 65968 57712
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 15883 1596 15949 1597
rect 15883 1532 15884 1596
rect 15948 1532 15949 1596
rect 15883 1531 15949 1532
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A0
timestamp 1649977179
transform 1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A
timestamp 1649977179
transform -1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A0
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A0
timestamp 1649977179
transform 1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A0
timestamp 1649977179
transform 1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A0
timestamp 1649977179
transform -1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A0
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A
timestamp 1649977179
transform 1 0 22264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A0
timestamp 1649977179
transform 1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A0
timestamp 1649977179
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A0
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A0
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A0
timestamp 1649977179
transform -1 0 3496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1649977179
transform 1 0 12788 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B
timestamp 1649977179
transform -1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1649977179
transform 1 0 5704 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A
timestamp 1649977179
transform 1 0 3036 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1649977179
transform 1 0 3680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1649977179
transform -1 0 1656 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A1
timestamp 1649977179
transform -1 0 1656 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1649977179
transform 1 0 4876 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A1
timestamp 1649977179
transform 1 0 3680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1649977179
transform 1 0 4784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A1
timestamp 1649977179
transform -1 0 3956 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1649977179
transform -1 0 5336 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1649977179
transform 1 0 3036 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A1
timestamp 1649977179
transform -1 0 5060 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1649977179
transform -1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1649977179
transform 1 0 3036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1649977179
transform 1 0 3956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A1
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A1
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1649977179
transform 1 0 13248 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1649977179
transform 1 0 3036 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1
timestamp 1649977179
transform 1 0 4416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1649977179
transform -1 0 1564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1649977179
transform -1 0 3864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A1
timestamp 1649977179
transform -1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A1
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1649977179
transform -1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1649977179
transform -1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1649977179
transform -1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A1
timestamp 1649977179
transform -1 0 4140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A1
timestamp 1649977179
transform -1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1649977179
transform -1 0 6900 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A1
timestamp 1649977179
transform -1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1649977179
transform 1 0 10212 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A1
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A1
timestamp 1649977179
transform -1 0 10948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A1
timestamp 1649977179
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A1
timestamp 1649977179
transform 1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__C1
timestamp 1649977179
transform -1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1649977179
transform 1 0 5704 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__C1
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__C1
timestamp 1649977179
transform -1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1649977179
transform -1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A1
timestamp 1649977179
transform -1 0 9108 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__C1
timestamp 1649977179
transform -1 0 8372 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__C1
timestamp 1649977179
transform 1 0 7636 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A1
timestamp 1649977179
transform -1 0 7360 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A1
timestamp 1649977179
transform 1 0 5704 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1649977179
transform 1 0 5704 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A1
timestamp 1649977179
transform 1 0 9568 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A1
timestamp 1649977179
transform 1 0 5704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp 1649977179
transform 1 0 12144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A1
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1649977179
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A1
timestamp 1649977179
transform -1 0 10120 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1
timestamp 1649977179
transform 1 0 14628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A1
timestamp 1649977179
transform -1 0 17572 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A1
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A1
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A1
timestamp 1649977179
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A1
timestamp 1649977179
transform 1 0 15456 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A1
timestamp 1649977179
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A1
timestamp 1649977179
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1649977179
transform 1 0 18032 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1649977179
transform -1 0 22632 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1649977179
transform -1 0 22080 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1649977179
transform 1 0 22632 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A1
timestamp 1649977179
transform 1 0 22356 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1649977179
transform 1 0 18584 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1649977179
transform 1 0 22632 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A1
timestamp 1649977179
transform 1 0 24840 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A1
timestamp 1649977179
transform 1 0 26312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A1
timestamp 1649977179
transform 1 0 26956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1649977179
transform 1 0 27876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1649977179
transform 1 0 28704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1649977179
transform 1 0 28336 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A1
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1649977179
transform 1 0 26312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1649977179
transform 1 0 28244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1649977179
transform -1 0 27140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1
timestamp 1649977179
transform 1 0 26864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1649977179
transform 1 0 23276 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A1
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1649977179
transform -1 0 24564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1649977179
transform 1 0 23184 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__C1
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1649977179
transform 1 0 24196 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1649977179
transform 1 0 25208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B
timestamp 1649977179
transform -1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A1
timestamp 1649977179
transform 1 0 30084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__C1
timestamp 1649977179
transform 1 0 29532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A1
timestamp 1649977179
transform 1 0 31188 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__C1
timestamp 1649977179
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1649977179
transform -1 0 33120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1649977179
transform -1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A1
timestamp 1649977179
transform 1 0 32384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__C1
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1649977179
transform -1 0 28980 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A1
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1649977179
transform 1 0 27876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A1
timestamp 1649977179
transform 1 0 31188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A1
timestamp 1649977179
transform -1 0 26404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A1
timestamp 1649977179
transform 1 0 27416 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1649977179
transform 1 0 26312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A1
timestamp 1649977179
transform 1 0 28704 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1649977179
transform 1 0 18584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1649977179
transform 1 0 32936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1649977179
transform 1 0 30636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1649977179
transform 1 0 36064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A1
timestamp 1649977179
transform 1 0 39652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A1
timestamp 1649977179
transform -1 0 41308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A1
timestamp 1649977179
transform 1 0 36156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A1
timestamp 1649977179
transform -1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A1
timestamp 1649977179
transform -1 0 35972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A1
timestamp 1649977179
transform 1 0 34684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A1
timestamp 1649977179
transform -1 0 34224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A1
timestamp 1649977179
transform 1 0 32936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1649977179
transform -1 0 33488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform 1 0 21160 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A
timestamp 1649977179
transform -1 0 30360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1649977179
transform -1 0 30636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A1
timestamp 1649977179
transform 1 0 32292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A1
timestamp 1649977179
transform 1 0 34040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1649977179
transform 1 0 39192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A1
timestamp 1649977179
transform -1 0 40204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A1
timestamp 1649977179
transform -1 0 39836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A1
timestamp 1649977179
transform 1 0 36340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A1
timestamp 1649977179
transform 1 0 36156 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A
timestamp 1649977179
transform -1 0 27232 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A1
timestamp 1649977179
transform -1 0 32292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A1
timestamp 1649977179
transform 1 0 30176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A1
timestamp 1649977179
transform -1 0 31372 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A1
timestamp 1649977179
transform -1 0 34868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1649977179
transform 1 0 31464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A
timestamp 1649977179
transform -1 0 33304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A1
timestamp 1649977179
transform 1 0 34224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 1649977179
transform 1 0 34040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A1
timestamp 1649977179
transform 1 0 35512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A1
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A1
timestamp 1649977179
transform 1 0 37628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1649977179
transform 1 0 35328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A1
timestamp 1649977179
transform 1 0 35328 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A1
timestamp 1649977179
transform -1 0 37444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1649977179
transform -1 0 34132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A1
timestamp 1649977179
transform -1 0 34868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A1
timestamp 1649977179
transform -1 0 33028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A
timestamp 1649977179
transform -1 0 22080 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1649977179
transform -1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1649977179
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A
timestamp 1649977179
transform 1 0 20516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A
timestamp 1649977179
transform -1 0 26772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A1
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A
timestamp 1649977179
transform -1 0 21252 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1
timestamp 1649977179
transform 1 0 20424 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A
timestamp 1649977179
transform 1 0 19044 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1
timestamp 1649977179
transform 1 0 20608 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A
timestamp 1649977179
transform 1 0 18584 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A1
timestamp 1649977179
transform -1 0 24564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A
timestamp 1649977179
transform -1 0 20516 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A1
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1649977179
transform -1 0 19412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A
timestamp 1649977179
transform 1 0 25852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A1
timestamp 1649977179
transform 1 0 24748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A
timestamp 1649977179
transform -1 0 18768 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1
timestamp 1649977179
transform -1 0 26404 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A
timestamp 1649977179
transform 1 0 16744 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A1
timestamp 1649977179
transform 1 0 25668 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1
timestamp 1649977179
transform -1 0 24564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__A
timestamp 1649977179
transform 1 0 21988 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1
timestamp 1649977179
transform 1 0 21160 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A
timestamp 1649977179
transform 1 0 18032 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A
timestamp 1649977179
transform 1 0 18584 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1
timestamp 1649977179
transform 1 0 21160 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A_N
timestamp 1649977179
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A
timestamp 1649977179
transform 1 0 29348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1649977179
transform -1 0 28244 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1649977179
transform -1 0 29992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A1
timestamp 1649977179
transform 1 0 29716 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A1
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A1
timestamp 1649977179
transform 1 0 30820 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A1
timestamp 1649977179
transform 1 0 32292 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A1
timestamp 1649977179
transform -1 0 33764 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1649977179
transform -1 0 32384 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1649977179
transform 1 0 31464 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1
timestamp 1649977179
transform -1 0 29072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__C1
timestamp 1649977179
transform 1 0 27600 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A1
timestamp 1649977179
transform 1 0 28152 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__C1
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A_N
timestamp 1649977179
transform -1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A
timestamp 1649977179
transform 1 0 14904 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A1
timestamp 1649977179
transform -1 0 15824 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__C1
timestamp 1649977179
transform 1 0 15824 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1649977179
transform -1 0 17940 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__C1
timestamp 1649977179
transform 1 0 18124 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A1
timestamp 1649977179
transform -1 0 18124 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__C1
timestamp 1649977179
transform 1 0 16928 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A1
timestamp 1649977179
transform 1 0 17480 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A1
timestamp 1649977179
transform 1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A1
timestamp 1649977179
transform -1 0 16928 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A1
timestamp 1649977179
transform 1 0 18032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A1
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A1
timestamp 1649977179
transform 1 0 17572 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1649977179
transform 1 0 17756 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A1
timestamp 1649977179
transform 1 0 16744 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A_N
timestamp 1649977179
transform -1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1649977179
transform -1 0 12144 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A1
timestamp 1649977179
transform 1 0 10212 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1649977179
transform 1 0 12420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A
timestamp 1649977179
transform -1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A1
timestamp 1649977179
transform 1 0 10028 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A1
timestamp 1649977179
transform -1 0 13524 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__A1
timestamp 1649977179
transform 1 0 13984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A1
timestamp 1649977179
transform 1 0 12788 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A1
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A
timestamp 1649977179
transform 1 0 21160 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A1
timestamp 1649977179
transform -1 0 15456 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1649977179
transform 1 0 14076 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A1
timestamp 1649977179
transform -1 0 13616 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A1
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__A
timestamp 1649977179
transform 1 0 21160 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A
timestamp 1649977179
transform 1 0 21344 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__B
timestamp 1649977179
transform -1 0 20332 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1649977179
transform 1 0 22632 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A
timestamp 1649977179
transform 1 0 21896 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__A1
timestamp 1649977179
transform 1 0 23000 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1649977179
transform -1 0 26496 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A1
timestamp 1649977179
transform 1 0 25208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__A1
timestamp 1649977179
transform 1 0 24656 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A1
timestamp 1649977179
transform 1 0 24656 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__A1
timestamp 1649977179
transform 1 0 27600 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A1
timestamp 1649977179
transform 1 0 27784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__A1
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A1
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__A1
timestamp 1649977179
transform -1 0 22908 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1649977179
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 1649977179
transform -1 0 22632 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__A
timestamp 1649977179
transform -1 0 19412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__A
timestamp 1649977179
transform 1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A1
timestamp 1649977179
transform 1 0 17112 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A1
timestamp 1649977179
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__A1
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A1
timestamp 1649977179
transform -1 0 20700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__A1
timestamp 1649977179
transform 1 0 18032 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__A
timestamp 1649977179
transform -1 0 23644 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A1
timestamp 1649977179
transform 1 0 27416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A1
timestamp 1649977179
transform 1 0 28796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__A1
timestamp 1649977179
transform 1 0 26864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A1
timestamp 1649977179
transform 1 0 24656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A1
timestamp 1649977179
transform -1 0 25116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A
timestamp 1649977179
transform -1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A1
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__A1
timestamp 1649977179
transform 1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__C
timestamp 1649977179
transform -1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__B
timestamp 1649977179
transform -1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A
timestamp 1649977179
transform -1 0 14720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__D
timestamp 1649977179
transform 1 0 29624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A
timestamp 1649977179
transform 1 0 21896 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__C
timestamp 1649977179
transform -1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__D
timestamp 1649977179
transform -1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A
timestamp 1649977179
transform 1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__A
timestamp 1649977179
transform -1 0 25944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__C
timestamp 1649977179
transform -1 0 14812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__D
timestamp 1649977179
transform -1 0 30728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__B1
timestamp 1649977179
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1561__B1
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__A2
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__B1
timestamp 1649977179
transform 1 0 18032 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__B1
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__A2
timestamp 1649977179
transform 1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__B1
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__A
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 20424 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_wb_clk_i_A
timestamp 1649977179
transform -1 0 30452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 11868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1649977179
transform 1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1649977179
transform 1 0 7728 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1649977179
transform 1 0 11316 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1649977179
transform 1 0 17112 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1649977179
transform 1 0 19872 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1649977179
transform -1 0 28060 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1649977179
transform 1 0 33396 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1649977179
transform 1 0 34776 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1649977179
transform 1 0 29072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1649977179
transform 1 0 33396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1649977179
transform 1 0 37352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1649977179
transform -1 0 35052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1649977179
transform 1 0 29624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1649977179
transform 1 0 26312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1649977179
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 23000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 22448 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 4048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 21988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 6808 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 4692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 12880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 2208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31
timestamp 1649977179
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_151 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_255
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_283
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_318
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_346
timestamp 1649977179
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_353
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_627
timestamp 1649977179
transform 1 0 58788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_634
timestamp 1649977179
transform 1 0 59432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 1649977179
transform 1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_648
timestamp 1649977179
transform 1 0 60720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_655
timestamp 1649977179
transform 1 0 61364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_662
timestamp 1649977179
transform 1 0 62008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_670
timestamp 1649977179
transform 1 0 62744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_676
timestamp 1649977179
transform 1 0 63296 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_683 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 63940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_695
timestamp 1649977179
transform 1 0 65044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1649977179
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_717
timestamp 1649977179
transform 1 0 67068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_724
timestamp 1649977179
transform 1 0 67712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_16
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_24
timestamp 1649977179
transform 1 0 3312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_41
timestamp 1649977179
transform 1 0 4876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_127
timestamp 1649977179
transform 1 0 12788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_227
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_290
timestamp 1649977179
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1649977179
transform 1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1649977179
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_318
timestamp 1649977179
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1649977179
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_346
timestamp 1649977179
transform 1 0 32936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_353
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_360
timestamp 1649977179
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_367
timestamp 1649977179
transform 1 0 34868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_376
timestamp 1649977179
transform 1 0 35696 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_627
timestamp 1649977179
transform 1 0 58788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_634
timestamp 1649977179
transform 1 0 59432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_641
timestamp 1649977179
transform 1 0 60076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_648
timestamp 1649977179
transform 1 0 60720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_655
timestamp 1649977179
transform 1 0 61364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_662
timestamp 1649977179
transform 1 0 62008 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_670
timestamp 1649977179
transform 1 0 62744 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_676
timestamp 1649977179
transform 1 0 63296 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_688
timestamp 1649977179
transform 1 0 64400 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_700
timestamp 1649977179
transform 1 0 65504 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_712
timestamp 1649977179
transform 1 0 66608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_724
timestamp 1649977179
transform 1 0 67712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_5
timestamp 1649977179
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_14
timestamp 1649977179
transform 1 0 2392 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1649977179
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_89
timestamp 1649977179
transform 1 0 9292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1649977179
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_120
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_149
timestamp 1649977179
transform 1 0 14812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_219
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_225
timestamp 1649977179
transform 1 0 21804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_229
timestamp 1649977179
transform 1 0 22172 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_238
timestamp 1649977179
transform 1 0 23000 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1649977179
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_256
timestamp 1649977179
transform 1 0 24656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_274
timestamp 1649977179
transform 1 0 26312 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_283
timestamp 1649977179
transform 1 0 27140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_292
timestamp 1649977179
transform 1 0 27968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_316
timestamp 1649977179
transform 1 0 30176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_325
timestamp 1649977179
transform 1 0 31004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_334
timestamp 1649977179
transform 1 0 31832 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_343
timestamp 1649977179
transform 1 0 32660 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_352
timestamp 1649977179
transform 1 0 33488 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_424
timestamp 1649977179
transform 1 0 40112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_431
timestamp 1649977179
transform 1 0 40756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_438
timestamp 1649977179
transform 1 0 41400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1649977179
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_461
timestamp 1649977179
transform 1 0 43516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1649977179
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_481
timestamp 1649977179
transform 1 0 45356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_488
timestamp 1649977179
transform 1 0 46000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_495
timestamp 1649977179
transform 1 0 46644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_502
timestamp 1649977179
transform 1 0 47288 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_511
timestamp 1649977179
transform 1 0 48116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_519
timestamp 1649977179
transform 1 0 48852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_523
timestamp 1649977179
transform 1 0 49220 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_538
timestamp 1649977179
transform 1 0 50600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_552
timestamp 1649977179
transform 1 0 51888 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_560
timestamp 1649977179
transform 1 0 52624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1649977179
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_620
timestamp 1649977179
transform 1 0 58144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_627
timestamp 1649977179
transform 1 0 58788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_634
timestamp 1649977179
transform 1 0 59432 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_642
timestamp 1649977179
transform 1 0 60168 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_648
timestamp 1649977179
transform 1 0 60720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_655
timestamp 1649977179
transform 1 0 61364 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_662
timestamp 1649977179
transform 1 0 62008 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_674
timestamp 1649977179
transform 1 0 63112 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_686
timestamp 1649977179
transform 1 0 64216 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_698
timestamp 1649977179
transform 1 0 65320 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_729
timestamp 1649977179
transform 1 0 68172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_40
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_59
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1649977179
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1649977179
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_123
timestamp 1649977179
transform 1 0 12420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_158
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1649977179
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1649977179
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_210
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1649977179
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_248
timestamp 1649977179
transform 1 0 23920 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1649977179
transform 1 0 24840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_270
timestamp 1649977179
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1649977179
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_297
timestamp 1649977179
transform 1 0 28428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_303
timestamp 1649977179
transform 1 0 28980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_307
timestamp 1649977179
transform 1 0 29348 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_324
timestamp 1649977179
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_371
timestamp 1649977179
transform 1 0 35236 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_379
timestamp 1649977179
transform 1 0 35972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_602
timestamp 1649977179
transform 1 0 56488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_620
timestamp 1649977179
transform 1 0 58144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_627
timestamp 1649977179
transform 1 0 58788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_634
timestamp 1649977179
transform 1 0 59432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_648
timestamp 1649977179
transform 1 0 60720 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_655
timestamp 1649977179
transform 1 0 61364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_667
timestamp 1649977179
transform 1 0 62468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_6
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1649977179
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_35
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_66
timestamp 1649977179
transform 1 0 7176 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_113
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_126
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_161
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1649977179
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_212
timestamp 1649977179
transform 1 0 20608 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_226
timestamp 1649977179
transform 1 0 21896 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1649977179
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_238
timestamp 1649977179
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_242
timestamp 1649977179
transform 1 0 23368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_269
timestamp 1649977179
transform 1 0 25852 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_278
timestamp 1649977179
transform 1 0 26680 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_290
timestamp 1649977179
transform 1 0 27784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_294
timestamp 1649977179
transform 1 0 28152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1649977179
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_329
timestamp 1649977179
transform 1 0 31372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_353
timestamp 1649977179
transform 1 0 33580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1649977179
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_369
timestamp 1649977179
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_409
timestamp 1649977179
transform 1 0 38732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 1649977179
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_609
timestamp 1649977179
transform 1 0 57132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_620
timestamp 1649977179
transform 1 0 58144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_627
timestamp 1649977179
transform 1 0 58788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_634
timestamp 1649977179
transform 1 0 59432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_642
timestamp 1649977179
transform 1 0 60168 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_648
timestamp 1649977179
transform 1 0 60720 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_660
timestamp 1649977179
transform 1 0 61824 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_672
timestamp 1649977179
transform 1 0 62928 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_684
timestamp 1649977179
transform 1 0 64032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_696
timestamp 1649977179
transform 1 0 65136 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_12
timestamp 1649977179
transform 1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1649977179
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_63
timestamp 1649977179
transform 1 0 6900 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_70
timestamp 1649977179
transform 1 0 7544 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_91
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_121
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_155
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_186
timestamp 1649977179
transform 1 0 18216 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_204
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_241
timestamp 1649977179
transform 1 0 23276 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp 1649977179
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_269
timestamp 1649977179
transform 1 0 25852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1649977179
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_289
timestamp 1649977179
transform 1 0 27692 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_298
timestamp 1649977179
transform 1 0 28520 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_312
timestamp 1649977179
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1649977179
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_339
timestamp 1649977179
transform 1 0 32292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_351
timestamp 1649977179
transform 1 0 33396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_360
timestamp 1649977179
transform 1 0 34224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_364
timestamp 1649977179
transform 1 0 34592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_387
timestamp 1649977179
transform 1 0 36708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_398
timestamp 1649977179
transform 1 0 37720 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_407
timestamp 1649977179
transform 1 0 38548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_419
timestamp 1649977179
transform 1 0 39652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_431
timestamp 1649977179
transform 1 0 40756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1649977179
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_625
timestamp 1649977179
transform 1 0 58604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_630
timestamp 1649977179
transform 1 0 59064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_637
timestamp 1649977179
transform 1 0 59708 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_644
timestamp 1649977179
transform 1 0 60352 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_656
timestamp 1649977179
transform 1 0 61456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_668
timestamp 1649977179
transform 1 0 62560 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_724
timestamp 1649977179
transform 1 0 67712 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_6
timestamp 1649977179
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_45
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_57
timestamp 1649977179
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_69
timestamp 1649977179
transform 1 0 7452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_73
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_95
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_120
timestamp 1649977179
transform 1 0 12144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_132
timestamp 1649977179
transform 1 0 13248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_156
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_176
timestamp 1649977179
transform 1 0 17296 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_205
timestamp 1649977179
transform 1 0 19964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_226
timestamp 1649977179
transform 1 0 21896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_232
timestamp 1649977179
transform 1 0 22448 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_236
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1649977179
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_261
timestamp 1649977179
transform 1 0 25116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1649977179
transform 1 0 25944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1649977179
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_282
timestamp 1649977179
transform 1 0 27048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1649977179
transform 1 0 27600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_300
timestamp 1649977179
transform 1 0 28704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_325
timestamp 1649977179
transform 1 0 31004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_337
timestamp 1649977179
transform 1 0 32108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_348
timestamp 1649977179
transform 1 0 33120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1649977179
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_393
timestamp 1649977179
transform 1 0 37260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_410
timestamp 1649977179
transform 1 0 38824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1649977179
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1649977179
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_16
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_25
timestamp 1649977179
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_37
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_45
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_73
timestamp 1649977179
transform 1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_80
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1649977179
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_101
timestamp 1649977179
transform 1 0 10396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1649977179
transform 1 0 15456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_160
timestamp 1649977179
transform 1 0 15824 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_171
timestamp 1649977179
transform 1 0 16836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_183
timestamp 1649977179
transform 1 0 17940 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_194
timestamp 1649977179
transform 1 0 18952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1649977179
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_243
timestamp 1649977179
transform 1 0 23460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_267
timestamp 1649977179
transform 1 0 25668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1649977179
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_283
timestamp 1649977179
transform 1 0 27140 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_291
timestamp 1649977179
transform 1 0 27876 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_312
timestamp 1649977179
transform 1 0 29808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_328
timestamp 1649977179
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_347
timestamp 1649977179
transform 1 0 33028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_351
timestamp 1649977179
transform 1 0 33396 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_357
timestamp 1649977179
transform 1 0 33948 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_367
timestamp 1649977179
transform 1 0 34868 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_379
timestamp 1649977179
transform 1 0 35972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_724
timestamp 1649977179
transform 1 0 67712 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1649977179
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1649977179
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_50
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_58
timestamp 1649977179
transform 1 0 6440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1649977179
transform 1 0 9660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_100
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_113
timestamp 1649977179
transform 1 0 11500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_120
timestamp 1649977179
transform 1 0 12144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_127
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_155
timestamp 1649977179
transform 1 0 15364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_159
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_176
timestamp 1649977179
transform 1 0 17296 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_182
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_213
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_230
timestamp 1649977179
transform 1 0 22264 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_260
timestamp 1649977179
transform 1 0 25024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1649977179
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_300
timestamp 1649977179
transform 1 0 28704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_325
timestamp 1649977179
transform 1 0 31004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_334
timestamp 1649977179
transform 1 0 31832 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_356
timestamp 1649977179
transform 1 0 33856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_371
timestamp 1649977179
transform 1 0 35236 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_383
timestamp 1649977179
transform 1 0 36340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_405
timestamp 1649977179
transform 1 0 38364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_414
timestamp 1649977179
transform 1 0 39192 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1649977179
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_21
timestamp 1649977179
transform 1 0 3036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_64
timestamp 1649977179
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_77
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_99
timestamp 1649977179
transform 1 0 10212 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp 1649977179
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_190
timestamp 1649977179
transform 1 0 18584 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_197
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_214
timestamp 1649977179
transform 1 0 20792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_230
timestamp 1649977179
transform 1 0 22264 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_238
timestamp 1649977179
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_243
timestamp 1649977179
transform 1 0 23460 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_267
timestamp 1649977179
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_285
timestamp 1649977179
transform 1 0 27324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_291
timestamp 1649977179
transform 1 0 27876 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_297
timestamp 1649977179
transform 1 0 28428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_309
timestamp 1649977179
transform 1 0 29532 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_315
timestamp 1649977179
transform 1 0 30084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_318
timestamp 1649977179
transform 1 0 30360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1649977179
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_345
timestamp 1649977179
transform 1 0 32844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_353
timestamp 1649977179
transform 1 0 33580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_358
timestamp 1649977179
transform 1 0 34040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_372
timestamp 1649977179
transform 1 0 35328 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_386
timestamp 1649977179
transform 1 0 36616 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_401
timestamp 1649977179
transform 1 0 37996 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_413
timestamp 1649977179
transform 1 0 39100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_425
timestamp 1649977179
transform 1 0 40204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_437
timestamp 1649977179
transform 1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1649977179
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_5
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_11
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_17
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_31
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1649977179
transform 1 0 5336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_95
timestamp 1649977179
transform 1 0 9844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_104
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_111
timestamp 1649977179
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_115
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1649977179
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1649977179
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp 1649977179
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_205
timestamp 1649977179
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_216
timestamp 1649977179
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_220
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1649977179
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_232
timestamp 1649977179
transform 1 0 22448 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1649977179
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_264
timestamp 1649977179
transform 1 0 25392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_276
timestamp 1649977179
transform 1 0 26496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_282
timestamp 1649977179
transform 1 0 27048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_286
timestamp 1649977179
transform 1 0 27416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_295
timestamp 1649977179
transform 1 0 28244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1649977179
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_329
timestamp 1649977179
transform 1 0 31372 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_337
timestamp 1649977179
transform 1 0 32108 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_349
timestamp 1649977179
transform 1 0 33212 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_352
timestamp 1649977179
transform 1 0 33488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_356
timestamp 1649977179
transform 1 0 33856 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_376
timestamp 1649977179
transform 1 0 35696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_380
timestamp 1649977179
transform 1 0 36064 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_729
timestamp 1649977179
transform 1 0 68172 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_21
timestamp 1649977179
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_41
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1649977179
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1649977179
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_77
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_88
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_148
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_176
timestamp 1649977179
transform 1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_196
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_204
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_241
timestamp 1649977179
transform 1 0 23276 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1649977179
transform 1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_260
timestamp 1649977179
transform 1 0 25024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_263
timestamp 1649977179
transform 1 0 25300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1649977179
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_289
timestamp 1649977179
transform 1 0 27692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_301
timestamp 1649977179
transform 1 0 28796 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_323
timestamp 1649977179
transform 1 0 30820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_344
timestamp 1649977179
transform 1 0 32752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_352
timestamp 1649977179
transform 1 0 33488 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_358
timestamp 1649977179
transform 1 0 34040 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_370
timestamp 1649977179
transform 1 0 35144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_379
timestamp 1649977179
transform 1 0 35972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_410
timestamp 1649977179
transform 1 0 38824 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_422
timestamp 1649977179
transform 1 0 39928 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_434
timestamp 1649977179
transform 1 0 41032 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1649977179
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_17
timestamp 1649977179
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1649977179
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_34
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_46
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_101
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp 1649977179
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_122
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_132
timestamp 1649977179
transform 1 0 13248 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 1649977179
transform 1 0 14720 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1649977179
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_173
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_203
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_227
timestamp 1649977179
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_239
timestamp 1649977179
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_260
timestamp 1649977179
transform 1 0 25024 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_273
timestamp 1649977179
transform 1 0 26220 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_285
timestamp 1649977179
transform 1 0 27324 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_292
timestamp 1649977179
transform 1 0 27968 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1649977179
transform 1 0 31004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_336
timestamp 1649977179
transform 1 0 32016 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_340
timestamp 1649977179
transform 1 0 32384 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_348
timestamp 1649977179
transform 1 0 33120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1649977179
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_367
timestamp 1649977179
transform 1 0 34868 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_387
timestamp 1649977179
transform 1 0 36708 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_399
timestamp 1649977179
transform 1 0 37812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_411
timestamp 1649977179
transform 1 0 38916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_729
timestamp 1649977179
transform 1 0 68172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_25
timestamp 1649977179
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_29
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_77
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_83
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_101
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_120
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_135
timestamp 1649977179
transform 1 0 13524 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_147
timestamp 1649977179
transform 1 0 14628 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_191
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_199
timestamp 1649977179
transform 1 0 19412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_207
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_213
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_228
timestamp 1649977179
transform 1 0 22080 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_234
timestamp 1649977179
transform 1 0 22632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_240
timestamp 1649977179
transform 1 0 23184 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_246
timestamp 1649977179
transform 1 0 23736 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_258
timestamp 1649977179
transform 1 0 24840 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_264
timestamp 1649977179
transform 1 0 25392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1649977179
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_287
timestamp 1649977179
transform 1 0 27508 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_296
timestamp 1649977179
transform 1 0 28336 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_302
timestamp 1649977179
transform 1 0 28888 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_314
timestamp 1649977179
transform 1 0 29992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_318
timestamp 1649977179
transform 1 0 30360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1649977179
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_340
timestamp 1649977179
transform 1 0 32384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_354
timestamp 1649977179
transform 1 0 33672 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_368
timestamp 1649977179
transform 1 0 34960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1649977179
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_412
timestamp 1649977179
transform 1 0 39008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_418
timestamp 1649977179
transform 1 0 39560 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_421
timestamp 1649977179
transform 1 0 39836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_433
timestamp 1649977179
transform 1 0 40940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1649977179
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_10
timestamp 1649977179
transform 1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_31
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_43
timestamp 1649977179
transform 1 0 5060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_55
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_71
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_112
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_149
timestamp 1649977179
transform 1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_169
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_181
timestamp 1649977179
transform 1 0 17756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1649977179
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_213
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1649977179
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1649977179
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_266
timestamp 1649977179
transform 1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_280
timestamp 1649977179
transform 1 0 26864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_290
timestamp 1649977179
transform 1 0 27784 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_296
timestamp 1649977179
transform 1 0 28336 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_316
timestamp 1649977179
transform 1 0 30176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_338
timestamp 1649977179
transform 1 0 32200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_356
timestamp 1649977179
transform 1 0 33856 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_370
timestamp 1649977179
transform 1 0 35144 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_378
timestamp 1649977179
transform 1 0 35880 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_390
timestamp 1649977179
transform 1 0 36984 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_402
timestamp 1649977179
transform 1 0 38088 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_410
timestamp 1649977179
transform 1 0 38824 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1649977179
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_429
timestamp 1649977179
transform 1 0 40572 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_441
timestamp 1649977179
transform 1 0 41676 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_453
timestamp 1649977179
transform 1 0 42780 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_465
timestamp 1649977179
transform 1 0 43884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1649977179
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_8
timestamp 1649977179
transform 1 0 1840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_63
timestamp 1649977179
transform 1 0 6900 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_83
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_94
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_120
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_132
timestamp 1649977179
transform 1 0 13248 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_150
timestamp 1649977179
transform 1 0 14904 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1649977179
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1649977179
transform 1 0 17388 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_183
timestamp 1649977179
transform 1 0 17940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_186
timestamp 1649977179
transform 1 0 18216 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1649977179
transform 1 0 19044 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_204
timestamp 1649977179
transform 1 0 19872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_228
timestamp 1649977179
transform 1 0 22080 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_234
timestamp 1649977179
transform 1 0 22632 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_242
timestamp 1649977179
transform 1 0 23368 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_255
timestamp 1649977179
transform 1 0 24564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_266
timestamp 1649977179
transform 1 0 25576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1649977179
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_289
timestamp 1649977179
transform 1 0 27692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_301
timestamp 1649977179
transform 1 0 28796 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_315
timestamp 1649977179
transform 1 0 30084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_321
timestamp 1649977179
transform 1 0 30636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1649977179
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_344
timestamp 1649977179
transform 1 0 32752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_353
timestamp 1649977179
transform 1 0 33580 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_369
timestamp 1649977179
transform 1 0 35052 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_377
timestamp 1649977179
transform 1 0 35788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_383
timestamp 1649977179
transform 1 0 36340 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_413
timestamp 1649977179
transform 1 0 39100 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_419
timestamp 1649977179
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_425
timestamp 1649977179
transform 1 0 40204 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_437
timestamp 1649977179
transform 1 0 41308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1649977179
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_724
timestamp 1649977179
transform 1 0 67712 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1649977179
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_103
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_116
timestamp 1649977179
transform 1 0 11776 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_124
timestamp 1649977179
transform 1 0 12512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1649977179
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_169
timestamp 1649977179
transform 1 0 16652 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1649977179
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_213
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_239
timestamp 1649977179
transform 1 0 23092 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_255
timestamp 1649977179
transform 1 0 24564 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_269
timestamp 1649977179
transform 1 0 25852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_297
timestamp 1649977179
transform 1 0 28428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1649977179
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1649977179
transform 1 0 30176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_322
timestamp 1649977179
transform 1 0 30728 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_344
timestamp 1649977179
transform 1 0 32752 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1649977179
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_372
timestamp 1649977179
transform 1 0 35328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_392
timestamp 1649977179
transform 1 0 37168 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_412
timestamp 1649977179
transform 1 0 39008 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_429
timestamp 1649977179
transform 1 0 40572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_441
timestamp 1649977179
transform 1 0 41676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_453
timestamp 1649977179
transform 1 0 42780 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_465
timestamp 1649977179
transform 1 0 43884 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_473
timestamp 1649977179
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_18
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_33
timestamp 1649977179
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1649977179
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1649977179
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_70
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_78
timestamp 1649977179
transform 1 0 8280 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_85
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_104
timestamp 1649977179
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1649977179
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_146
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1649977179
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_211
timestamp 1649977179
transform 1 0 20516 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_228
timestamp 1649977179
transform 1 0 22080 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_242
timestamp 1649977179
transform 1 0 23368 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1649977179
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_289
timestamp 1649977179
transform 1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_304
timestamp 1649977179
transform 1 0 29072 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_308
timestamp 1649977179
transform 1 0 29440 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_315
timestamp 1649977179
transform 1 0 30084 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_323
timestamp 1649977179
transform 1 0 30820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1649977179
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_341
timestamp 1649977179
transform 1 0 32476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_347
timestamp 1649977179
transform 1 0 33028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_356
timestamp 1649977179
transform 1 0 33856 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_364
timestamp 1649977179
transform 1 0 34592 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_410
timestamp 1649977179
transform 1 0 38824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_418
timestamp 1649977179
transform 1 0 39560 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_426
timestamp 1649977179
transform 1 0 40296 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_438
timestamp 1649977179
transform 1 0 41400 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1649977179
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_724
timestamp 1649977179
transform 1 0 67712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_47
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_75
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_119
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1649977179
transform 1 0 14536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_175
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_179
timestamp 1649977179
transform 1 0 17572 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1649977179
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_199
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_211
timestamp 1649977179
transform 1 0 20516 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_231
timestamp 1649977179
transform 1 0 22356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_235
timestamp 1649977179
transform 1 0 22724 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1649977179
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1649977179
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1649977179
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_268
timestamp 1649977179
transform 1 0 25760 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_283
timestamp 1649977179
transform 1 0 27140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_295
timestamp 1649977179
transform 1 0 28244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1649977179
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_318
timestamp 1649977179
transform 1 0 30360 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_340
timestamp 1649977179
transform 1 0 32384 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_348
timestamp 1649977179
transform 1 0 33120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1649977179
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_368
timestamp 1649977179
transform 1 0 34960 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_392
timestamp 1649977179
transform 1 0 37168 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1649977179
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_431
timestamp 1649977179
transform 1 0 40756 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_437
timestamp 1649977179
transform 1 0 41308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_449
timestamp 1649977179
transform 1 0 42412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_461
timestamp 1649977179
transform 1 0 43516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1649977179
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1649977179
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_16
timestamp 1649977179
transform 1 0 2576 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_22
timestamp 1649977179
transform 1 0 3128 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1649977179
transform 1 0 3680 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_45
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_72
timestamp 1649977179
transform 1 0 7728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_76
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_102
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1649977179
transform 1 0 12420 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_134
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_187
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1649977179
transform 1 0 19136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_227
timestamp 1649977179
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_233
timestamp 1649977179
transform 1 0 22540 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_236
timestamp 1649977179
transform 1 0 22816 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_244
timestamp 1649977179
transform 1 0 23552 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_253
timestamp 1649977179
transform 1 0 24380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_259
timestamp 1649977179
transform 1 0 24932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_268
timestamp 1649977179
transform 1 0 25760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1649977179
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_289
timestamp 1649977179
transform 1 0 27692 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_295
timestamp 1649977179
transform 1 0 28244 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_298
timestamp 1649977179
transform 1 0 28520 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1649977179
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_312
timestamp 1649977179
transform 1 0 29808 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_324
timestamp 1649977179
transform 1 0 30912 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1649977179
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_344
timestamp 1649977179
transform 1 0 32752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_350
timestamp 1649977179
transform 1 0 33304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_381
timestamp 1649977179
transform 1 0 36156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1649977179
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_396
timestamp 1649977179
transform 1 0 37536 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_408
timestamp 1649977179
transform 1 0 38640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_414
timestamp 1649977179
transform 1 0 39192 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_428
timestamp 1649977179
transform 1 0 40480 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_440
timestamp 1649977179
transform 1 0 41584 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1649977179
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_10
timestamp 1649977179
transform 1 0 2024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1649977179
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1649977179
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_68
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_74
timestamp 1649977179
transform 1 0 7912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_95
timestamp 1649977179
transform 1 0 9844 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_103
timestamp 1649977179
transform 1 0 10580 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_124
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_147
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_171
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_175
timestamp 1649977179
transform 1 0 17204 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_202
timestamp 1649977179
transform 1 0 19688 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_228
timestamp 1649977179
transform 1 0 22080 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1649977179
transform 1 0 22816 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1649977179
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_260
timestamp 1649977179
transform 1 0 25024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_280
timestamp 1649977179
transform 1 0 26864 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_286
timestamp 1649977179
transform 1 0 27416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1649977179
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1649977179
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_332
timestamp 1649977179
transform 1 0 31648 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_338
timestamp 1649977179
transform 1 0 32200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_341
timestamp 1649977179
transform 1 0 32476 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_352
timestamp 1649977179
transform 1 0 33488 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_367
timestamp 1649977179
transform 1 0 34868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_376
timestamp 1649977179
transform 1 0 35696 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_382
timestamp 1649977179
transform 1 0 36248 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_394
timestamp 1649977179
transform 1 0 37352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_412
timestamp 1649977179
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_429
timestamp 1649977179
transform 1 0 40572 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_438
timestamp 1649977179
transform 1 0 41400 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_450
timestamp 1649977179
transform 1 0 42504 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_462
timestamp 1649977179
transform 1 0 43608 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_474
timestamp 1649977179
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_725
timestamp 1649977179
transform 1 0 67804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_729
timestamp 1649977179
transform 1 0 68172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_33
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_41
timestamp 1649977179
transform 1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_61
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_130
timestamp 1649977179
transform 1 0 13064 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_138
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_151
timestamp 1649977179
transform 1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_206
timestamp 1649977179
transform 1 0 20056 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_212
timestamp 1649977179
transform 1 0 20608 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1649977179
transform 1 0 22540 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1649977179
transform 1 0 23644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1649977179
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_260
timestamp 1649977179
transform 1 0 25024 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_272
timestamp 1649977179
transform 1 0 26128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1649977179
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_290
timestamp 1649977179
transform 1 0 27784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_307
timestamp 1649977179
transform 1 0 29348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_321
timestamp 1649977179
transform 1 0 30636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1649977179
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_352
timestamp 1649977179
transform 1 0 33488 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_356
timestamp 1649977179
transform 1 0 33856 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_377
timestamp 1649977179
transform 1 0 35788 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_386
timestamp 1649977179
transform 1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_413
timestamp 1649977179
transform 1 0 39100 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_416
timestamp 1649977179
transform 1 0 39376 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_425
timestamp 1649977179
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1649977179
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1649977179
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1649977179
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1649977179
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1649977179
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1649977179
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_47
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_58
timestamp 1649977179
transform 1 0 6440 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_64
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1649977179
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1649977179
transform 1 0 9200 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_106
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 1649977179
transform 1 0 12972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1649977179
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1649977179
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1649977179
transform 1 0 15640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_161
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_170
timestamp 1649977179
transform 1 0 16744 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_176
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_182
timestamp 1649977179
transform 1 0 17848 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_199
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_205
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1649977179
transform 1 0 20700 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_216
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1649977179
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_229
timestamp 1649977179
transform 1 0 22172 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1649977179
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1649977179
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_259
timestamp 1649977179
transform 1 0 24932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_271
timestamp 1649977179
transform 1 0 26036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_279
timestamp 1649977179
transform 1 0 26772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_285
timestamp 1649977179
transform 1 0 27324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1649977179
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_292
timestamp 1649977179
transform 1 0 27968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_297
timestamp 1649977179
transform 1 0 28428 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1649977179
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_325
timestamp 1649977179
transform 1 0 31004 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_331
timestamp 1649977179
transform 1 0 31556 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_339
timestamp 1649977179
transform 1 0 32292 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 1649977179
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1649977179
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_370
timestamp 1649977179
transform 1 0 35144 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_392
timestamp 1649977179
transform 1 0 37168 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1649977179
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_429
timestamp 1649977179
transform 1 0 40572 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_441
timestamp 1649977179
transform 1 0 41676 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_453
timestamp 1649977179
transform 1 0 42780 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_465
timestamp 1649977179
transform 1 0 43884 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1649977179
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1649977179
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1649977179
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1649977179
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1649977179
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_725
timestamp 1649977179
transform 1 0 67804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_729
timestamp 1649977179
transform 1 0 68172 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_11
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_24
timestamp 1649977179
transform 1 0 3312 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_36
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_42
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_67
timestamp 1649977179
transform 1 0 7268 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_87
timestamp 1649977179
transform 1 0 9108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1649977179
transform 1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_117
timestamp 1649977179
transform 1 0 11868 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1649977179
transform 1 0 12420 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1649977179
transform 1 0 17112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_198
timestamp 1649977179
transform 1 0 19320 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1649977179
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_213
timestamp 1649977179
transform 1 0 20700 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1649977179
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_251
timestamp 1649977179
transform 1 0 24196 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_289
timestamp 1649977179
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_310
timestamp 1649977179
transform 1 0 29624 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_316
timestamp 1649977179
transform 1 0 30176 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_319
timestamp 1649977179
transform 1 0 30452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1649977179
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_353
timestamp 1649977179
transform 1 0 33580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_377
timestamp 1649977179
transform 1 0 35788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_386
timestamp 1649977179
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_421
timestamp 1649977179
transform 1 0 39836 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_433
timestamp 1649977179
transform 1 0 40940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_445
timestamp 1649977179
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1649977179
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1649977179
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_9
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1649977179
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_58
timestamp 1649977179
transform 1 0 6440 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1649977179
transform 1 0 6992 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_72
timestamp 1649977179
transform 1 0 7728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_92
timestamp 1649977179
transform 1 0 9568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1649977179
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1649977179
transform 1 0 12972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1649977179
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_143
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_158
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1649977179
transform 1 0 20424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1649977179
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_224
timestamp 1649977179
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1649977179
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_242
timestamp 1649977179
transform 1 0 23368 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1649977179
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_255
timestamp 1649977179
transform 1 0 24564 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_267
timestamp 1649977179
transform 1 0 25668 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_275
timestamp 1649977179
transform 1 0 26404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1649977179
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_296
timestamp 1649977179
transform 1 0 28336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1649977179
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_319
timestamp 1649977179
transform 1 0 30452 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_347
timestamp 1649977179
transform 1 0 33028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1649977179
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_367
timestamp 1649977179
transform 1 0 34868 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_379
timestamp 1649977179
transform 1 0 35972 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_391
timestamp 1649977179
transform 1 0 37076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_395
timestamp 1649977179
transform 1 0 37444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_412
timestamp 1649977179
transform 1 0 39008 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1649977179
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1649977179
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1649977179
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_24
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_30
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_63
timestamp 1649977179
transform 1 0 6900 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_71
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_88
timestamp 1649977179
transform 1 0 9200 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_127
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_143
timestamp 1649977179
transform 1 0 14260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_155
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_179
timestamp 1649977179
transform 1 0 17572 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_189
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_195
timestamp 1649977179
transform 1 0 19044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_212
timestamp 1649977179
transform 1 0 20608 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_233
timestamp 1649977179
transform 1 0 22540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_239
timestamp 1649977179
transform 1 0 23092 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1649977179
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_253
timestamp 1649977179
transform 1 0 24380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_264
timestamp 1649977179
transform 1 0 25392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 1649977179
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_301
timestamp 1649977179
transform 1 0 28796 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_321
timestamp 1649977179
transform 1 0 30636 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1649977179
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_367
timestamp 1649977179
transform 1 0 34868 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_371
timestamp 1649977179
transform 1 0 35236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_374
timestamp 1649977179
transform 1 0 35512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_386
timestamp 1649977179
transform 1 0 36616 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_398
timestamp 1649977179
transform 1 0 37720 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_410
timestamp 1649977179
transform 1 0 38824 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_422
timestamp 1649977179
transform 1 0 39928 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_434
timestamp 1649977179
transform 1 0 41032 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1649977179
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_724
timestamp 1649977179
transform 1 0 67712 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_17
timestamp 1649977179
transform 1 0 2668 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_34
timestamp 1649977179
transform 1 0 4232 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_64
timestamp 1649977179
transform 1 0 6992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1649977179
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_95
timestamp 1649977179
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_101
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1649977179
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_146
timestamp 1649977179
transform 1 0 14536 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1649977179
transform 1 0 15272 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_158
timestamp 1649977179
transform 1 0 15640 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1649977179
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_184
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1649977179
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_218
timestamp 1649977179
transform 1 0 21160 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1649977179
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1649977179
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_269
timestamp 1649977179
transform 1 0 25852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_276
timestamp 1649977179
transform 1 0 26496 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1649977179
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_316
timestamp 1649977179
transform 1 0 30176 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_332
timestamp 1649977179
transform 1 0 31648 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_338
timestamp 1649977179
transform 1 0 32200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_344
timestamp 1649977179
transform 1 0 32752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_350
timestamp 1649977179
transform 1 0 33304 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_356
timestamp 1649977179
transform 1 0 33856 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1649977179
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_370
timestamp 1649977179
transform 1 0 35144 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_394
timestamp 1649977179
transform 1 0 37352 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_414
timestamp 1649977179
transform 1 0 39192 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1649977179
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_14
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_63
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_75
timestamp 1649977179
transform 1 0 8004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1649977179
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1649977179
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1649977179
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1649977179
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1649977179
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_180
timestamp 1649977179
transform 1 0 17664 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_263
timestamp 1649977179
transform 1 0 25300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1649977179
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_300
timestamp 1649977179
transform 1 0 28704 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1649977179
transform 1 0 29256 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1649977179
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_341
timestamp 1649977179
transform 1 0 32476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_350
timestamp 1649977179
transform 1 0 33304 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_358
timestamp 1649977179
transform 1 0 34040 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_362
timestamp 1649977179
transform 1 0 34408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_376
timestamp 1649977179
transform 1 0 35696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1649977179
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_395
timestamp 1649977179
transform 1 0 37444 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_403
timestamp 1649977179
transform 1 0 38180 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_411
timestamp 1649977179
transform 1 0 38916 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_423
timestamp 1649977179
transform 1 0 40020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_435
timestamp 1649977179
transform 1 0 41124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1649977179
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1649977179
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_724
timestamp 1649977179
transform 1 0 67712 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_5
timestamp 1649977179
transform 1 0 1564 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_17
timestamp 1649977179
transform 1 0 2668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1649977179
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_45
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_62
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1649977179
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1649977179
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_119
timestamp 1649977179
transform 1 0 12052 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_125
timestamp 1649977179
transform 1 0 12604 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1649977179
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_151
timestamp 1649977179
transform 1 0 14996 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_164
timestamp 1649977179
transform 1 0 16192 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_172
timestamp 1649977179
transform 1 0 16928 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_181
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_206
timestamp 1649977179
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_217
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_223
timestamp 1649977179
transform 1 0 21620 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1649977179
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_255
timestamp 1649977179
transform 1 0 24564 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_261
timestamp 1649977179
transform 1 0 25116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_273
timestamp 1649977179
transform 1 0 26220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_282
timestamp 1649977179
transform 1 0 27048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_290
timestamp 1649977179
transform 1 0 27784 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_293
timestamp 1649977179
transform 1 0 28060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1649977179
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_316
timestamp 1649977179
transform 1 0 30176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_322
timestamp 1649977179
transform 1 0 30728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_339
timestamp 1649977179
transform 1 0 32292 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_347
timestamp 1649977179
transform 1 0 33028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1649977179
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_368
timestamp 1649977179
transform 1 0 34960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_374
timestamp 1649977179
transform 1 0 35512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_388
timestamp 1649977179
transform 1 0 36800 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_396
timestamp 1649977179
transform 1 0 37536 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_399
timestamp 1649977179
transform 1 0 37812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_411
timestamp 1649977179
transform 1 0 38916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1649977179
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1649977179
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1649977179
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1649977179
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_19
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1649977179
transform 1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_66
timestamp 1649977179
transform 1 0 7176 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_72
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_79
timestamp 1649977179
transform 1 0 8372 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_87
timestamp 1649977179
transform 1 0 9108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_90
timestamp 1649977179
transform 1 0 9384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_133
timestamp 1649977179
transform 1 0 13340 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1649977179
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1649977179
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_178
timestamp 1649977179
transform 1 0 17480 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_186
timestamp 1649977179
transform 1 0 18216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1649977179
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_228
timestamp 1649977179
transform 1 0 22080 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_242
timestamp 1649977179
transform 1 0 23368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_253
timestamp 1649977179
transform 1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_264
timestamp 1649977179
transform 1 0 25392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1649977179
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1649977179
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_291
timestamp 1649977179
transform 1 0 27876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_297
timestamp 1649977179
transform 1 0 28428 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_308
timestamp 1649977179
transform 1 0 29440 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_314
timestamp 1649977179
transform 1 0 29992 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_323
timestamp 1649977179
transform 1 0 30820 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_339
timestamp 1649977179
transform 1 0 32292 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_347
timestamp 1649977179
transform 1 0 33028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_359
timestamp 1649977179
transform 1 0 34132 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_362
timestamp 1649977179
transform 1 0 34408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_376
timestamp 1649977179
transform 1 0 35696 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_397
timestamp 1649977179
transform 1 0 37628 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_414
timestamp 1649977179
transform 1 0 39192 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_426
timestamp 1649977179
transform 1 0 40296 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_438
timestamp 1649977179
transform 1 0 41400 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1649977179
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_17
timestamp 1649977179
transform 1 0 2668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1649977179
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_57
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_66
timestamp 1649977179
transform 1 0 7176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1649977179
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_95
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_106
timestamp 1649977179
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_112
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_129
timestamp 1649977179
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1649977179
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_143
timestamp 1649977179
transform 1 0 14260 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_181
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1649977179
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_231
timestamp 1649977179
transform 1 0 22356 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_237
timestamp 1649977179
transform 1 0 22908 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1649977179
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_283
timestamp 1649977179
transform 1 0 27140 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_303
timestamp 1649977179
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_319
timestamp 1649977179
transform 1 0 30452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_326
timestamp 1649977179
transform 1 0 31096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_330
timestamp 1649977179
transform 1 0 31464 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_347
timestamp 1649977179
transform 1 0 33028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1649977179
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_373
timestamp 1649977179
transform 1 0 35420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_397
timestamp 1649977179
transform 1 0 37628 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_403
timestamp 1649977179
transform 1 0 38180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_415
timestamp 1649977179
transform 1 0 39284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_729
timestamp 1649977179
transform 1 0 68172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_12
timestamp 1649977179
transform 1 0 2208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_32
timestamp 1649977179
transform 1 0 4048 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_101
timestamp 1649977179
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1649977179
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_118
timestamp 1649977179
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1649977179
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_134
timestamp 1649977179
transform 1 0 13432 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_138
timestamp 1649977179
transform 1 0 13800 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_147
timestamp 1649977179
transform 1 0 14628 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1649977179
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1649977179
transform 1 0 16928 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_196
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_199
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1649977179
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_233
timestamp 1649977179
transform 1 0 22540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_242
timestamp 1649977179
transform 1 0 23368 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_248
timestamp 1649977179
transform 1 0 23920 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_256
timestamp 1649977179
transform 1 0 24656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1649977179
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1649977179
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1649977179
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_339
timestamp 1649977179
transform 1 0 32292 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_351
timestamp 1649977179
transform 1 0 33396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_369
timestamp 1649977179
transform 1 0 35052 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_377
timestamp 1649977179
transform 1 0 35788 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_386
timestamp 1649977179
transform 1 0 36616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_398
timestamp 1649977179
transform 1 0 37720 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_410
timestamp 1649977179
transform 1 0 38824 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_422
timestamp 1649977179
transform 1 0 39928 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_434
timestamp 1649977179
transform 1 0 41032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1649977179
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1649977179
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1649977179
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_39
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_42
timestamp 1649977179
transform 1 0 4968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_50
timestamp 1649977179
transform 1 0 5704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_54
timestamp 1649977179
transform 1 0 6072 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1649977179
transform 1 0 6900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_94
timestamp 1649977179
transform 1 0 9752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_143
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_155
timestamp 1649977179
transform 1 0 15364 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_175
timestamp 1649977179
transform 1 0 17204 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_181
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_186
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_213
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_235
timestamp 1649977179
transform 1 0 22724 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1649977179
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_260
timestamp 1649977179
transform 1 0 25024 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_268
timestamp 1649977179
transform 1 0 25760 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_292
timestamp 1649977179
transform 1 0 27968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_322
timestamp 1649977179
transform 1 0 30728 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_342
timestamp 1649977179
transform 1 0 32568 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_354
timestamp 1649977179
transform 1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1649977179
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_368
timestamp 1649977179
transform 1 0 34960 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1649977179
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_385
timestamp 1649977179
transform 1 0 36524 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_729
timestamp 1649977179
transform 1 0 68172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_6
timestamp 1649977179
transform 1 0 1656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_18
timestamp 1649977179
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_30
timestamp 1649977179
transform 1 0 3864 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_36
timestamp 1649977179
transform 1 0 4416 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_48
timestamp 1649977179
transform 1 0 5520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1649977179
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1649977179
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_67
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_71
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_80
timestamp 1649977179
transform 1 0 8464 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_86
timestamp 1649977179
transform 1 0 9016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_92
timestamp 1649977179
transform 1 0 9568 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_98
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_115
timestamp 1649977179
transform 1 0 11684 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_143
timestamp 1649977179
transform 1 0 14260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_174
timestamp 1649977179
transform 1 0 17112 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_196
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1649977179
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_227
timestamp 1649977179
transform 1 0 21988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_231
timestamp 1649977179
transform 1 0 22356 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_248
timestamp 1649977179
transform 1 0 23920 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_256
timestamp 1649977179
transform 1 0 24656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1649977179
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1649977179
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_289
timestamp 1649977179
transform 1 0 27692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_297
timestamp 1649977179
transform 1 0 28428 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1649977179
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_342
timestamp 1649977179
transform 1 0 32568 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_364
timestamp 1649977179
transform 1 0 34592 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1649977179
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_395
timestamp 1649977179
transform 1 0 37444 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_407
timestamp 1649977179
transform 1 0 38548 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_419
timestamp 1649977179
transform 1 0 39652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_431
timestamp 1649977179
transform 1 0 40756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1649977179
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_7
timestamp 1649977179
transform 1 0 1748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1649977179
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1649977179
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_45
timestamp 1649977179
transform 1 0 5244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_57
timestamp 1649977179
transform 1 0 6348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_90
timestamp 1649977179
transform 1 0 9384 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_98
timestamp 1649977179
transform 1 0 10120 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_104
timestamp 1649977179
transform 1 0 10672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_116
timestamp 1649977179
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_122
timestamp 1649977179
transform 1 0 12328 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_128
timestamp 1649977179
transform 1 0 12880 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1649977179
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1649977179
transform 1 0 14812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1649977179
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_173
timestamp 1649977179
transform 1 0 17020 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_179
timestamp 1649977179
transform 1 0 17572 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_183
timestamp 1649977179
transform 1 0 17940 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_186
timestamp 1649977179
transform 1 0 18216 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1649977179
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_201
timestamp 1649977179
transform 1 0 19596 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1649977179
transform 1 0 20056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_210
timestamp 1649977179
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1649977179
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_237
timestamp 1649977179
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1649977179
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_258
timestamp 1649977179
transform 1 0 24840 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_270
timestamp 1649977179
transform 1 0 25944 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_290
timestamp 1649977179
transform 1 0 27784 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1649977179
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_323
timestamp 1649977179
transform 1 0 30820 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1649977179
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_338
timestamp 1649977179
transform 1 0 32200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_350
timestamp 1649977179
transform 1 0 33304 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1649977179
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_374
timestamp 1649977179
transform 1 0 35512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_388
timestamp 1649977179
transform 1 0 36800 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_400
timestamp 1649977179
transform 1 0 37904 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_412
timestamp 1649977179
transform 1 0 39008 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1649977179
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1649977179
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_45
timestamp 1649977179
transform 1 0 5244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1649977179
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1649977179
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_62
timestamp 1649977179
transform 1 0 6808 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_74
timestamp 1649977179
transform 1 0 7912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_86
timestamp 1649977179
transform 1 0 9016 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_104
timestamp 1649977179
transform 1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_138
timestamp 1649977179
transform 1 0 13800 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1649977179
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_189
timestamp 1649977179
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_194
timestamp 1649977179
transform 1 0 18952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1649977179
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_238
timestamp 1649977179
transform 1 0 23000 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_247
timestamp 1649977179
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_259
timestamp 1649977179
transform 1 0 24932 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_268
timestamp 1649977179
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_289
timestamp 1649977179
transform 1 0 27692 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_296
timestamp 1649977179
transform 1 0 28336 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_308
timestamp 1649977179
transform 1 0 29440 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_311
timestamp 1649977179
transform 1 0 29716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_344
timestamp 1649977179
transform 1 0 32752 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_368
timestamp 1649977179
transform 1 0 34960 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_372
timestamp 1649977179
transform 1 0 35328 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_375
timestamp 1649977179
transform 1 0 35604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1649977179
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_411
timestamp 1649977179
transform 1 0 38916 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_423
timestamp 1649977179
transform 1 0 40020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_435
timestamp 1649977179
transform 1 0 41124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_724
timestamp 1649977179
transform 1 0 67712 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_8
timestamp 1649977179
transform 1 0 1840 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_17
timestamp 1649977179
transform 1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1649977179
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1649977179
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1649977179
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1649977179
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1649977179
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_95
timestamp 1649977179
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 1649977179
transform 1 0 10212 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1649977179
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_122
timestamp 1649977179
transform 1 0 12328 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1649977179
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_157
timestamp 1649977179
transform 1 0 15548 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_169
timestamp 1649977179
transform 1 0 16652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_183
timestamp 1649977179
transform 1 0 17940 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_204
timestamp 1649977179
transform 1 0 19872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1649977179
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_219
timestamp 1649977179
transform 1 0 21252 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_222
timestamp 1649977179
transform 1 0 21528 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1649977179
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_244
timestamp 1649977179
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_261
timestamp 1649977179
transform 1 0 25116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_282
timestamp 1649977179
transform 1 0 27048 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_290
timestamp 1649977179
transform 1 0 27784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1649977179
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_325
timestamp 1649977179
transform 1 0 31004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_342
timestamp 1649977179
transform 1 0 32568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_354
timestamp 1649977179
transform 1 0 33672 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1649977179
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_383
timestamp 1649977179
transform 1 0 36340 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_395
timestamp 1649977179
transform 1 0 37444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_407
timestamp 1649977179
transform 1 0 38548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_16
timestamp 1649977179
transform 1 0 2576 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_38
timestamp 1649977179
transform 1 0 4600 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_46
timestamp 1649977179
transform 1 0 5336 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1649977179
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_90
timestamp 1649977179
transform 1 0 9384 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1649977179
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1649977179
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_140
timestamp 1649977179
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_143
timestamp 1649977179
transform 1 0 14260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_155
timestamp 1649977179
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1649977179
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_201
timestamp 1649977179
transform 1 0 19596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_209
timestamp 1649977179
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1649977179
transform 1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1649977179
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_228
timestamp 1649977179
transform 1 0 22080 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_242
timestamp 1649977179
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_248
timestamp 1649977179
transform 1 0 23920 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_260
timestamp 1649977179
transform 1 0 25024 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_272
timestamp 1649977179
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_309
timestamp 1649977179
transform 1 0 29532 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_325
timestamp 1649977179
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_342
timestamp 1649977179
transform 1 0 32568 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_348
timestamp 1649977179
transform 1 0 33120 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_360
timestamp 1649977179
transform 1 0 34224 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_372
timestamp 1649977179
transform 1 0 35328 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_384
timestamp 1649977179
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_409
timestamp 1649977179
transform 1 0 38732 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_421
timestamp 1649977179
transform 1 0 39836 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_433
timestamp 1649977179
transform 1 0 40940 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_445
timestamp 1649977179
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_724
timestamp 1649977179
transform 1 0 67712 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_19
timestamp 1649977179
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_33
timestamp 1649977179
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_50
timestamp 1649977179
transform 1 0 5704 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_56
timestamp 1649977179
transform 1 0 6256 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_88
timestamp 1649977179
transform 1 0 9200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_94
timestamp 1649977179
transform 1 0 9752 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_100
timestamp 1649977179
transform 1 0 10304 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_108
timestamp 1649977179
transform 1 0 11040 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_116
timestamp 1649977179
transform 1 0 11776 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_130
timestamp 1649977179
transform 1 0 13064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1649977179
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_157
timestamp 1649977179
transform 1 0 15548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_169
timestamp 1649977179
transform 1 0 16652 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_181
timestamp 1649977179
transform 1 0 17756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1649977179
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_199
timestamp 1649977179
transform 1 0 19412 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_218
timestamp 1649977179
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_227
timestamp 1649977179
transform 1 0 21988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1649977179
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_257
timestamp 1649977179
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_263
timestamp 1649977179
transform 1 0 25300 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_269
timestamp 1649977179
transform 1 0 25852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_297
timestamp 1649977179
transform 1 0 28428 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1649977179
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_314
timestamp 1649977179
transform 1 0 29992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_334
timestamp 1649977179
transform 1 0 31832 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_346
timestamp 1649977179
transform 1 0 32936 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_355
timestamp 1649977179
transform 1 0 33764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_17
timestamp 1649977179
transform 1 0 2668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_23
timestamp 1649977179
transform 1 0 3220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_45
timestamp 1649977179
transform 1 0 5244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_49
timestamp 1649977179
transform 1 0 5612 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1649977179
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_64
timestamp 1649977179
transform 1 0 6992 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_84
timestamp 1649977179
transform 1 0 8832 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1649977179
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_141
timestamp 1649977179
transform 1 0 14076 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_147
timestamp 1649977179
transform 1 0 14628 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1649977179
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1649977179
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_182
timestamp 1649977179
transform 1 0 17848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_191
timestamp 1649977179
transform 1 0 18676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_197
timestamp 1649977179
transform 1 0 19228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_214
timestamp 1649977179
transform 1 0 20792 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1649977179
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1649977179
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_242
timestamp 1649977179
transform 1 0 23368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_254
timestamp 1649977179
transform 1 0 24472 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_270
timestamp 1649977179
transform 1 0 25944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1649977179
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_296
timestamp 1649977179
transform 1 0 28336 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_308
timestamp 1649977179
transform 1 0 29440 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_319
timestamp 1649977179
transform 1 0 30452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1649977179
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_348
timestamp 1649977179
transform 1 0 33120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_368
timestamp 1649977179
transform 1 0 34960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1649977179
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_10
timestamp 1649977179
transform 1 0 2024 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1649977179
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_37
timestamp 1649977179
transform 1 0 4508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_43
timestamp 1649977179
transform 1 0 5060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_47
timestamp 1649977179
transform 1 0 5428 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_68
timestamp 1649977179
transform 1 0 7360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1649977179
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1649977179
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1649977179
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_95
timestamp 1649977179
transform 1 0 9844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1649977179
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_112
timestamp 1649977179
transform 1 0 11408 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_124
timestamp 1649977179
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1649977179
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_150
timestamp 1649977179
transform 1 0 14904 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_156
timestamp 1649977179
transform 1 0 15456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_168
timestamp 1649977179
transform 1 0 16560 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_183
timestamp 1649977179
transform 1 0 17940 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_186
timestamp 1649977179
transform 1 0 18216 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1649977179
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1649977179
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_211
timestamp 1649977179
transform 1 0 20516 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1649977179
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_226
timestamp 1649977179
transform 1 0 21896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1649977179
transform 1 0 22908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1649977179
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1649977179
transform 1 0 24564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_259
timestamp 1649977179
transform 1 0 24932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1649977179
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_291
timestamp 1649977179
transform 1 0 27876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_295
timestamp 1649977179
transform 1 0 28244 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1649977179
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_325
timestamp 1649977179
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_334
timestamp 1649977179
transform 1 0 31832 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_340
timestamp 1649977179
transform 1 0 32384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_349
timestamp 1649977179
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1649977179
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_729
timestamp 1649977179
transform 1 0 68172 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_20
timestamp 1649977179
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_32
timestamp 1649977179
transform 1 0 4048 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_37
timestamp 1649977179
transform 1 0 4508 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1649977179
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_60
timestamp 1649977179
transform 1 0 6624 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_64
timestamp 1649977179
transform 1 0 6992 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_75
timestamp 1649977179
transform 1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_95
timestamp 1649977179
transform 1 0 9844 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_107
timestamp 1649977179
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_121
timestamp 1649977179
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_127
timestamp 1649977179
transform 1 0 12788 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1649977179
transform 1 0 13156 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_140
timestamp 1649977179
transform 1 0 13984 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1649977179
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_172
timestamp 1649977179
transform 1 0 16928 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1649977179
transform 1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_191
timestamp 1649977179
transform 1 0 18676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1649977179
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_209
timestamp 1649977179
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1649977179
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_230
timestamp 1649977179
transform 1 0 22264 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_252
timestamp 1649977179
transform 1 0 24288 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_256
timestamp 1649977179
transform 1 0 24656 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_259
timestamp 1649977179
transform 1 0 24932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_271
timestamp 1649977179
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_289
timestamp 1649977179
transform 1 0 27692 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_295
timestamp 1649977179
transform 1 0 28244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_307
timestamp 1649977179
transform 1 0 29348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_315
timestamp 1649977179
transform 1 0 30084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_320
timestamp 1649977179
transform 1 0 30544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1649977179
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_341
timestamp 1649977179
transform 1 0 32476 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_355
timestamp 1649977179
transform 1 0 33764 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_363
timestamp 1649977179
transform 1 0 34500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_381
timestamp 1649977179
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1649977179
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1649977179
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_31
timestamp 1649977179
transform 1 0 3956 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_51
timestamp 1649977179
transform 1 0 5796 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_59
timestamp 1649977179
transform 1 0 6532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_66
timestamp 1649977179
transform 1 0 7176 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1649977179
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_101
timestamp 1649977179
transform 1 0 10396 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_118
timestamp 1649977179
transform 1 0 11960 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_130
timestamp 1649977179
transform 1 0 13064 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1649977179
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1649977179
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_152
timestamp 1649977179
transform 1 0 15088 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_160
timestamp 1649977179
transform 1 0 15824 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_170
timestamp 1649977179
transform 1 0 16744 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_178
timestamp 1649977179
transform 1 0 17480 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_184
timestamp 1649977179
transform 1 0 18032 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1649977179
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_213
timestamp 1649977179
transform 1 0 20700 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_217
timestamp 1649977179
transform 1 0 21068 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_220
timestamp 1649977179
transform 1 0 21344 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_227
timestamp 1649977179
transform 1 0 21988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_239
timestamp 1649977179
transform 1 0 23092 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1649977179
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1649977179
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_275
timestamp 1649977179
transform 1 0 26404 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_295
timestamp 1649977179
transform 1 0 28244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_319
timestamp 1649977179
transform 1 0 30452 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_327
timestamp 1649977179
transform 1 0 31188 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_339
timestamp 1649977179
transform 1 0 32292 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_353
timestamp 1649977179
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1649977179
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1649977179
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_729
timestamp 1649977179
transform 1 0 68172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_12
timestamp 1649977179
transform 1 0 2208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_24
timestamp 1649977179
transform 1 0 3312 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_30
timestamp 1649977179
transform 1 0 3864 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_42
timestamp 1649977179
transform 1 0 4968 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1649977179
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_65
timestamp 1649977179
transform 1 0 7084 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_118
timestamp 1649977179
transform 1 0 11960 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_126
timestamp 1649977179
transform 1 0 12696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_129
timestamp 1649977179
transform 1 0 12972 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1649977179
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_154
timestamp 1649977179
transform 1 0 15272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_158
timestamp 1649977179
transform 1 0 15640 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1649977179
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_191
timestamp 1649977179
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_213
timestamp 1649977179
transform 1 0 20700 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1649977179
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_251
timestamp 1649977179
transform 1 0 24196 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_255
timestamp 1649977179
transform 1 0 24564 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1649977179
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_283
timestamp 1649977179
transform 1 0 27140 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_291
timestamp 1649977179
transform 1 0 27876 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_302
timestamp 1649977179
transform 1 0 28888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_322
timestamp 1649977179
transform 1 0 30728 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1649977179
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_11
timestamp 1649977179
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_17
timestamp 1649977179
transform 1 0 2668 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1649977179
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_45
timestamp 1649977179
transform 1 0 5244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_57
timestamp 1649977179
transform 1 0 6348 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_61
timestamp 1649977179
transform 1 0 6716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_78
timestamp 1649977179
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_106
timestamp 1649977179
transform 1 0 10856 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_118
timestamp 1649977179
transform 1 0 11960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_127
timestamp 1649977179
transform 1 0 12788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1649977179
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_144
timestamp 1649977179
transform 1 0 14352 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_158
timestamp 1649977179
transform 1 0 15640 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_169
timestamp 1649977179
transform 1 0 16652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_172
timestamp 1649977179
transform 1 0 16928 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_180
timestamp 1649977179
transform 1 0 17664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1649977179
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_201
timestamp 1649977179
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_212
timestamp 1649977179
transform 1 0 20608 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_232
timestamp 1649977179
transform 1 0 22448 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1649977179
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_269
timestamp 1649977179
transform 1 0 25852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_278
timestamp 1649977179
transform 1 0 26680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_284
timestamp 1649977179
transform 1 0 27232 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_290
timestamp 1649977179
transform 1 0 27784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_298
timestamp 1649977179
transform 1 0 28520 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1649977179
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_317
timestamp 1649977179
transform 1 0 30268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1649977179
transform 1 0 31372 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_349
timestamp 1649977179
transform 1 0 33212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp 1649977179
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_11
timestamp 1649977179
transform 1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_21
timestamp 1649977179
transform 1 0 3036 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_41
timestamp 1649977179
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1649977179
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_67
timestamp 1649977179
transform 1 0 7268 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_73
timestamp 1649977179
transform 1 0 7820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_85
timestamp 1649977179
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_97
timestamp 1649977179
transform 1 0 10028 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1649977179
transform 1 0 10948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_117
timestamp 1649977179
transform 1 0 11868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_120
timestamp 1649977179
transform 1 0 12144 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_129
timestamp 1649977179
transform 1 0 12972 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_143
timestamp 1649977179
transform 1 0 14260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_151
timestamp 1649977179
transform 1 0 14996 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_159
timestamp 1649977179
transform 1 0 15732 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1649977179
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_179
timestamp 1649977179
transform 1 0 17572 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_213
timestamp 1649977179
transform 1 0 20700 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1649977179
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_230
timestamp 1649977179
transform 1 0 22264 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1649977179
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_263
timestamp 1649977179
transform 1 0 25300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_267
timestamp 1649977179
transform 1 0 25668 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1649977179
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_299
timestamp 1649977179
transform 1 0 28612 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_308
timestamp 1649977179
transform 1 0 29440 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_319
timestamp 1649977179
transform 1 0 30452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_325
timestamp 1649977179
transform 1 0 31004 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_333
timestamp 1649977179
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1649977179
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1649977179
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1649977179
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1649977179
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1649977179
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1649977179
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_724
timestamp 1649977179
transform 1 0 67712 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1649977179
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_18
timestamp 1649977179
transform 1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1649977179
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_61
timestamp 1649977179
transform 1 0 6716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_68
timestamp 1649977179
transform 1 0 7360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1649977179
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_101
timestamp 1649977179
transform 1 0 10396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_105
timestamp 1649977179
transform 1 0 10764 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_114
timestamp 1649977179
transform 1 0 11592 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_122
timestamp 1649977179
transform 1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1649977179
transform 1 0 12788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1649977179
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_149
timestamp 1649977179
transform 1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_157
timestamp 1649977179
transform 1 0 15548 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_168
timestamp 1649977179
transform 1 0 16560 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_176
timestamp 1649977179
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_190
timestamp 1649977179
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_202
timestamp 1649977179
transform 1 0 19688 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_212
timestamp 1649977179
transform 1 0 20608 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_222
timestamp 1649977179
transform 1 0 21528 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_226
timestamp 1649977179
transform 1 0 21896 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1649977179
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1649977179
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1649977179
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_264
timestamp 1649977179
transform 1 0 25392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_273
timestamp 1649977179
transform 1 0 26220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_279
timestamp 1649977179
transform 1 0 26772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_287
timestamp 1649977179
transform 1 0 27508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1649977179
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_311
timestamp 1649977179
transform 1 0 29716 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_323
timestamp 1649977179
transform 1 0 30820 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_335
timestamp 1649977179
transform 1 0 31924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_347
timestamp 1649977179
transform 1 0 33028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1649977179
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1649977179
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1649977179
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1649977179
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1649977179
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1649977179
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1649977179
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1649977179
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1649977179
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_12
timestamp 1649977179
transform 1 0 2208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_24
timestamp 1649977179
transform 1 0 3312 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_30
timestamp 1649977179
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_42
timestamp 1649977179
transform 1 0 4968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_46
timestamp 1649977179
transform 1 0 5336 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1649977179
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_63
timestamp 1649977179
transform 1 0 6900 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_71
timestamp 1649977179
transform 1 0 7636 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_77
timestamp 1649977179
transform 1 0 8188 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_92
timestamp 1649977179
transform 1 0 9568 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1649977179
transform 1 0 12328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_136
timestamp 1649977179
transform 1 0 13616 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_156
timestamp 1649977179
transform 1 0 15456 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1649977179
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_183
timestamp 1649977179
transform 1 0 17940 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_189
timestamp 1649977179
transform 1 0 18492 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_197
timestamp 1649977179
transform 1 0 19228 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_211
timestamp 1649977179
transform 1 0 20516 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1649977179
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_232
timestamp 1649977179
transform 1 0 22448 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1649977179
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_258
timestamp 1649977179
transform 1 0 24840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_270
timestamp 1649977179
transform 1 0 25944 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1649977179
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_289
timestamp 1649977179
transform 1 0 27692 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_295
timestamp 1649977179
transform 1 0 28244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_299
timestamp 1649977179
transform 1 0 28612 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_308
timestamp 1649977179
transform 1 0 29440 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_314
timestamp 1649977179
transform 1 0 29992 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_318
timestamp 1649977179
transform 1 0 30360 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_324
timestamp 1649977179
transform 1 0 30912 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_353
timestamp 1649977179
transform 1 0 33580 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_365
timestamp 1649977179
transform 1 0 34684 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_377
timestamp 1649977179
transform 1 0 35788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1649977179
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1649977179
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1649977179
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1649977179
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1649977179
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1649977179
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1649977179
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1649977179
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1649977179
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1649977179
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_724
timestamp 1649977179
transform 1 0 67712 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1649977179
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_14
timestamp 1649977179
transform 1 0 2392 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1649977179
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_48
timestamp 1649977179
transform 1 0 5520 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_56
timestamp 1649977179
transform 1 0 6256 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_67
timestamp 1649977179
transform 1 0 7268 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1649977179
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_87
timestamp 1649977179
transform 1 0 9108 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1649977179
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_113
timestamp 1649977179
transform 1 0 11500 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_119
timestamp 1649977179
transform 1 0 12052 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_128
timestamp 1649977179
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_160
timestamp 1649977179
transform 1 0 15824 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_172
timestamp 1649977179
transform 1 0 16928 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1649977179
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_218
timestamp 1649977179
transform 1 0 21160 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_226
timestamp 1649977179
transform 1 0 21896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_230
timestamp 1649977179
transform 1 0 22264 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_236
timestamp 1649977179
transform 1 0 22816 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1649977179
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_261
timestamp 1649977179
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_267
timestamp 1649977179
transform 1 0 25668 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_291
timestamp 1649977179
transform 1 0 27876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_303
timestamp 1649977179
transform 1 0 28980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_313
timestamp 1649977179
transform 1 0 29900 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_325
timestamp 1649977179
transform 1 0 31004 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_337
timestamp 1649977179
transform 1 0 32108 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_349
timestamp 1649977179
transform 1 0 33212 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1649977179
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1649977179
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1649977179
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1649977179
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1649977179
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1649977179
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1649977179
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1649977179
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1649977179
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1649977179
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1649977179
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1649977179
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1649977179
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_73
timestamp 1649977179
transform 1 0 7820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_79
timestamp 1649977179
transform 1 0 8372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_85
timestamp 1649977179
transform 1 0 8924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1649977179
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_121
timestamp 1649977179
transform 1 0 12236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_130
timestamp 1649977179
transform 1 0 13064 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_152
timestamp 1649977179
transform 1 0 15088 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1649977179
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_174
timestamp 1649977179
transform 1 0 17112 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_180
timestamp 1649977179
transform 1 0 17664 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_192
timestamp 1649977179
transform 1 0 18768 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_204
timestamp 1649977179
transform 1 0 19872 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_228
timestamp 1649977179
transform 1 0 22080 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_256
timestamp 1649977179
transform 1 0 24656 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_268
timestamp 1649977179
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_289
timestamp 1649977179
transform 1 0 27692 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_299
timestamp 1649977179
transform 1 0 28612 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_327
timestamp 1649977179
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_353
timestamp 1649977179
transform 1 0 33580 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_365
timestamp 1649977179
transform 1 0 34684 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_377
timestamp 1649977179
transform 1 0 35788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1649977179
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1649977179
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1649977179
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1649977179
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1649977179
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1649977179
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1649977179
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1649977179
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1649977179
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1649977179
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1649977179
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1649977179
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1649977179
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_45
timestamp 1649977179
transform 1 0 5244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_57
timestamp 1649977179
transform 1 0 6348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_69
timestamp 1649977179
transform 1 0 7452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_81
timestamp 1649977179
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_117
timestamp 1649977179
transform 1 0 11868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_129
timestamp 1649977179
transform 1 0 12972 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1649977179
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_169
timestamp 1649977179
transform 1 0 16652 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_175
timestamp 1649977179
transform 1 0 17204 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_214
timestamp 1649977179
transform 1 0 20792 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_226
timestamp 1649977179
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_235
timestamp 1649977179
transform 1 0 22724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_239
timestamp 1649977179
transform 1 0 23092 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1649977179
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_255
timestamp 1649977179
transform 1 0 24564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_275
timestamp 1649977179
transform 1 0 26404 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_295
timestamp 1649977179
transform 1 0 28244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1649977179
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1649977179
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1649977179
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1649977179
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1649977179
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1649977179
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1649977179
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1649977179
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1649977179
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1649977179
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1649977179
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_725
timestamp 1649977179
transform 1 0 67804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_729
timestamp 1649977179
transform 1 0 68172 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_35
timestamp 1649977179
transform 1 0 4324 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1649977179
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_61
timestamp 1649977179
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_78
timestamp 1649977179
transform 1 0 8280 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_84
timestamp 1649977179
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_99
timestamp 1649977179
transform 1 0 10212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_118
timestamp 1649977179
transform 1 0 11960 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_124
timestamp 1649977179
transform 1 0 12512 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_141
timestamp 1649977179
transform 1 0 14076 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_153
timestamp 1649977179
transform 1 0 15180 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_159
timestamp 1649977179
transform 1 0 15732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_174
timestamp 1649977179
transform 1 0 17112 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_194
timestamp 1649977179
transform 1 0 18952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1649977179
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1649977179
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_241
timestamp 1649977179
transform 1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_250
timestamp 1649977179
transform 1 0 24104 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_258
timestamp 1649977179
transform 1 0 24840 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1649977179
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_310
timestamp 1649977179
transform 1 0 29624 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_322
timestamp 1649977179
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1649977179
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1649977179
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1649977179
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1649977179
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1649977179
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1649977179
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1649977179
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1649977179
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1649977179
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1649977179
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1649977179
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1649977179
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1649977179
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_73
timestamp 1649977179
transform 1 0 7820 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1649977179
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_95
timestamp 1649977179
transform 1 0 9844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_101
timestamp 1649977179
transform 1 0 10396 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_119
timestamp 1649977179
transform 1 0 12052 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_125
timestamp 1649977179
transform 1 0 12604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1649977179
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_149
timestamp 1649977179
transform 1 0 14812 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_158
timestamp 1649977179
transform 1 0 15640 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1649977179
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_179
timestamp 1649977179
transform 1 0 17572 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_185
timestamp 1649977179
transform 1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1649977179
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_205
timestamp 1649977179
transform 1 0 19964 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_213
timestamp 1649977179
transform 1 0 20700 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_225
timestamp 1649977179
transform 1 0 21804 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1649977179
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1649977179
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_255
timestamp 1649977179
transform 1 0 24564 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_267
timestamp 1649977179
transform 1 0 25668 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_279
timestamp 1649977179
transform 1 0 26772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_291
timestamp 1649977179
transform 1 0 27876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1649977179
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1649977179
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1649977179
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1649977179
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1649977179
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1649977179
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1649977179
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1649977179
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1649977179
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1649977179
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1649977179
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1649977179
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_725
timestamp 1649977179
transform 1 0 67804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_729
timestamp 1649977179
transform 1 0 68172 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_86
timestamp 1649977179
transform 1 0 9016 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_98
timestamp 1649977179
transform 1 0 10120 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1649977179
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_124
timestamp 1649977179
transform 1 0 12512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1649977179
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_142
timestamp 1649977179
transform 1 0 14168 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_150
timestamp 1649977179
transform 1 0 14904 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_156
timestamp 1649977179
transform 1 0 15456 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1649977179
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_187
timestamp 1649977179
transform 1 0 18308 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_199
timestamp 1649977179
transform 1 0 19412 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_207
timestamp 1649977179
transform 1 0 20148 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1649977179
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_227
timestamp 1649977179
transform 1 0 21988 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_239
timestamp 1649977179
transform 1 0 23092 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_246
timestamp 1649977179
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_258
timestamp 1649977179
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1649977179
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1649977179
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1649977179
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1649977179
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1649977179
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1649977179
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1649977179
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1649977179
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1649977179
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1649977179
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1649977179
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1649977179
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1649977179
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1649977179
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_157
timestamp 1649977179
transform 1 0 15548 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_160
timestamp 1649977179
transform 1 0 15824 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_172
timestamp 1649977179
transform 1 0 16928 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_180
timestamp 1649977179
transform 1 0 17664 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_183
timestamp 1649977179
transform 1 0 17940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1649977179
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1649977179
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1649977179
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1649977179
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1649977179
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1649977179
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1649977179
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1649977179
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1649977179
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1649977179
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1649977179
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_725
timestamp 1649977179
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1649977179
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1649977179
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1649977179
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1649977179
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1649977179
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1649977179
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1649977179
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1649977179
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1649977179
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_724
timestamp 1649977179
transform 1 0 67712 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1649977179
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1649977179
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1649977179
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1649977179
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1649977179
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1649977179
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1649977179
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1649977179
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1649977179
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1649977179
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1649977179
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1649977179
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_725
timestamp 1649977179
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1649977179
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1649977179
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1649977179
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1649977179
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1649977179
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1649977179
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1649977179
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1649977179
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1649977179
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_724
timestamp 1649977179
transform 1 0 67712 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1649977179
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1649977179
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1649977179
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1649977179
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1649977179
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1649977179
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1649977179
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1649977179
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1649977179
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1649977179
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1649977179
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1649977179
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_725
timestamp 1649977179
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1649977179
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1649977179
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1649977179
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1649977179
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1649977179
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1649977179
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1649977179
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1649977179
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1649977179
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1649977179
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1649977179
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1649977179
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1649977179
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1649977179
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1649977179
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1649977179
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1649977179
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1649977179
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1649977179
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1649977179
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1649977179
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1649977179
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1649977179
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_725
timestamp 1649977179
transform 1 0 67804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_729
timestamp 1649977179
transform 1 0 68172 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1649977179
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1649977179
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1649977179
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1649977179
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1649977179
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1649977179
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1649977179
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1649977179
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1649977179
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1649977179
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1649977179
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1649977179
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1649977179
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1649977179
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1649977179
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1649977179
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1649977179
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1649977179
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1649977179
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1649977179
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1649977179
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1649977179
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1649977179
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_725
timestamp 1649977179
transform 1 0 67804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_729
timestamp 1649977179
transform 1 0 68172 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_629
timestamp 1649977179
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_641
timestamp 1649977179
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_653
timestamp 1649977179
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1649977179
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1649977179
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1649977179
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1649977179
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1649977179
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1649977179
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1649977179
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1649977179
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1649977179
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_625
timestamp 1649977179
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1649977179
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1649977179
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1649977179
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1649977179
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_669
timestamp 1649977179
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_681
timestamp 1649977179
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1649977179
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1649977179
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1649977179
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1649977179
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1649977179
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1649977179
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1649977179
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1649977179
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1649977179
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1649977179
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1649977179
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1649977179
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1649977179
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_709
timestamp 1649977179
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_724
timestamp 1649977179
transform 1 0 67712 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1649977179
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_625
timestamp 1649977179
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1649977179
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1649977179
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1649977179
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_657
timestamp 1649977179
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_669
timestamp 1649977179
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_681
timestamp 1649977179
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1649977179
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1649977179
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1649977179
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_713
timestamp 1649977179
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_725
timestamp 1649977179
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1649977179
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_641
timestamp 1649977179
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_653
timestamp 1649977179
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1649977179
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1649977179
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_673
timestamp 1649977179
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_685
timestamp 1649977179
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_697
timestamp 1649977179
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_709
timestamp 1649977179
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_724
timestamp 1649977179
transform 1 0 67712 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1649977179
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_625
timestamp 1649977179
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1649977179
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1649977179
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_645
timestamp 1649977179
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_657
timestamp 1649977179
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_669
timestamp 1649977179
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_681
timestamp 1649977179
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1649977179
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1649977179
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1649977179
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_713
timestamp 1649977179
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_725
timestamp 1649977179
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1649977179
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_641
timestamp 1649977179
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_653
timestamp 1649977179
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1649977179
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1649977179
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1649977179
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1649977179
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1649977179
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_709
timestamp 1649977179
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_721
timestamp 1649977179
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1649977179
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1649977179
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_625
timestamp 1649977179
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1649977179
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1649977179
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1649977179
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1649977179
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1649977179
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1649977179
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1649977179
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1649977179
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1649977179
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_713
timestamp 1649977179
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_725
timestamp 1649977179
transform 1 0 67804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_729
timestamp 1649977179
transform 1 0 68172 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_629
timestamp 1649977179
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_641
timestamp 1649977179
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_653
timestamp 1649977179
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1649977179
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1649977179
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1649977179
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1649977179
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1649977179
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1649977179
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1649977179
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1649977179
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1649977179
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1649977179
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1649977179
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1649977179
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1649977179
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1649977179
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1649977179
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1649977179
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1649977179
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1649977179
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1649977179
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_713
timestamp 1649977179
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_725
timestamp 1649977179
transform 1 0 67804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_729
timestamp 1649977179
transform 1 0 68172 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1649977179
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1649977179
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1649977179
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1649977179
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1649977179
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1649977179
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1649977179
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1649977179
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1649977179
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1649977179
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1649977179
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1649977179
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_625
timestamp 1649977179
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1649977179
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1649977179
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1649977179
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1649977179
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1649977179
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1649977179
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1649977179
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1649977179
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1649977179
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1649977179
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_725
timestamp 1649977179
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1649977179
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1649977179
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1649977179
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1649977179
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1649977179
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1649977179
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1649977179
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1649977179
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1649977179
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_724
timestamp 1649977179
transform 1 0 67712 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1649977179
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1649977179
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1649977179
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1649977179
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1649977179
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1649977179
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1649977179
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1649977179
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1649977179
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1649977179
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1649977179
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_713
timestamp 1649977179
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_725
timestamp 1649977179
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1649977179
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1649977179
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1649977179
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1649977179
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1649977179
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1649977179
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1649977179
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1649977179
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1649977179
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_724
timestamp 1649977179
transform 1 0 67712 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1649977179
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1649977179
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1649977179
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1649977179
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1649977179
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1649977179
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1649977179
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1649977179
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1649977179
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1649977179
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1649977179
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_713
timestamp 1649977179
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_725
timestamp 1649977179
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1649977179
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1649977179
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1649977179
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1649977179
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1649977179
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1649977179
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1649977179
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1649977179
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_709
timestamp 1649977179
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1649977179
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1649977179
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1649977179
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1649977179
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1649977179
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1649977179
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1649977179
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1649977179
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1649977179
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1649977179
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1649977179
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1649977179
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1649977179
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1649977179
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_725
timestamp 1649977179
transform 1 0 67804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_729
timestamp 1649977179
transform 1 0 68172 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1649977179
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1649977179
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1649977179
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1649977179
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1649977179
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1649977179
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1649977179
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1649977179
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1649977179
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1649977179
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1649977179
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1649977179
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1649977179
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1649977179
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1649977179
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1649977179
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1649977179
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1649977179
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1649977179
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1649977179
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1649977179
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_701
timestamp 1649977179
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_713
timestamp 1649977179
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_725
timestamp 1649977179
transform 1 0 67804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_729
timestamp 1649977179
transform 1 0 68172 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1649977179
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1649977179
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1649977179
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1649977179
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1649977179
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1649977179
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_685
timestamp 1649977179
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_697
timestamp 1649977179
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_709
timestamp 1649977179
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1649977179
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1649977179
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1649977179
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1649977179
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1649977179
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1649977179
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1649977179
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1649977179
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1649977179
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1649977179
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1649977179
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1649977179
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1649977179
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1649977179
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_725
timestamp 1649977179
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1649977179
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1649977179
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1649977179
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1649977179
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1649977179
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1649977179
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1649977179
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1649977179
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_709
timestamp 1649977179
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_724
timestamp 1649977179
transform 1 0 67712 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1649977179
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1649977179
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1649977179
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1649977179
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1649977179
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1649977179
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1649977179
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1649977179
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1649977179
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1649977179
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1649977179
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1649977179
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1649977179
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1649977179
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1649977179
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1649977179
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1649977179
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1649977179
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_673
timestamp 1649977179
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_685
timestamp 1649977179
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_697
timestamp 1649977179
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_709
timestamp 1649977179
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_724
timestamp 1649977179
transform 1 0 67712 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1649977179
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1649977179
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1649977179
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1649977179
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1649977179
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1649977179
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_669
timestamp 1649977179
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_681
timestamp 1649977179
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1649977179
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1649977179
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1649977179
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1649977179
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_725
timestamp 1649977179
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1649977179
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1649977179
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1649977179
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1649977179
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1649977179
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_673
timestamp 1649977179
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_685
timestamp 1649977179
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_697
timestamp 1649977179
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_709
timestamp 1649977179
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1649977179
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1649977179
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1649977179
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1649977179
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1649977179
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1649977179
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1649977179
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1649977179
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1649977179
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1649977179
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1649977179
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1649977179
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1649977179
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1649977179
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_725
timestamp 1649977179
transform 1 0 67804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_729
timestamp 1649977179
transform 1 0 68172 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1649977179
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1649977179
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1649977179
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1649977179
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1649977179
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1649977179
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1649977179
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1649977179
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1649977179
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1649977179
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1649977179
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1649977179
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1649977179
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1649977179
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1649977179
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1649977179
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1649977179
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1649977179
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1649977179
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1649977179
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1649977179
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1649977179
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1649977179
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_725
timestamp 1649977179
transform 1 0 67804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_729
timestamp 1649977179
transform 1 0 68172 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1649977179
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1649977179
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1649977179
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1649977179
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1649977179
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1649977179
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1649977179
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1649977179
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1649977179
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1649977179
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1649977179
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1649977179
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1649977179
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1649977179
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1649977179
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1649977179
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1649977179
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1649977179
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1649977179
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1649977179
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1649977179
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_701
timestamp 1649977179
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_713
timestamp 1649977179
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_725
timestamp 1649977179
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1649977179
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1649977179
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1649977179
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1649977179
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1649977179
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1649977179
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1649977179
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1649977179
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1649977179
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_724
timestamp 1649977179
transform 1 0 67712 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1649977179
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_625
timestamp 1649977179
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1649977179
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1649977179
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1649977179
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1649977179
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1649977179
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1649977179
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1649977179
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1649977179
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1649977179
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1649977179
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_725
timestamp 1649977179
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_629
timestamp 1649977179
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_641
timestamp 1649977179
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_653
timestamp 1649977179
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1649977179
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1649977179
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1649977179
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1649977179
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1649977179
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1649977179
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_724
timestamp 1649977179
transform 1 0 67712 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1649977179
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_625
timestamp 1649977179
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1649977179
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1649977179
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_645
timestamp 1649977179
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_657
timestamp 1649977179
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_669
timestamp 1649977179
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_681
timestamp 1649977179
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1649977179
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1649977179
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1649977179
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1649977179
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_725
timestamp 1649977179
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1649977179
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_629
timestamp 1649977179
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_641
timestamp 1649977179
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_653
timestamp 1649977179
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1649977179
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1649977179
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1649977179
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1649977179
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1649977179
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_709
timestamp 1649977179
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1649977179
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1649977179
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1649977179
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1649977179
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1649977179
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1649977179
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1649977179
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1649977179
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1649977179
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1649977179
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1649977179
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_625
timestamp 1649977179
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1649977179
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1649977179
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_645
timestamp 1649977179
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_657
timestamp 1649977179
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_669
timestamp 1649977179
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_681
timestamp 1649977179
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1649977179
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1649977179
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1649977179
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1649977179
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_725
timestamp 1649977179
transform 1 0 67804 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_729
timestamp 1649977179
transform 1 0 68172 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1649977179
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1649977179
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_29
timestamp 1649977179
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_41
timestamp 1649977179
transform 1 0 4876 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_48
timestamp 1649977179
transform 1 0 5520 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1649977179
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1649977179
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1649977179
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1649977179
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1649977179
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1649977179
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 1649977179
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_156
timestamp 1649977179
transform 1 0 15456 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1649977179
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1649977179
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_197
timestamp 1649977179
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1649977179
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1649977179
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1649977179
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1649977179
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_253
timestamp 1649977179
transform 1 0 24380 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_264
timestamp 1649977179
transform 1 0 25392 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_276
timestamp 1649977179
transform 1 0 26496 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1649977179
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1649977179
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_321
timestamp 1649977179
transform 1 0 30636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1649977179
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1649977179
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1649977179
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_365
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_372
timestamp 1649977179
transform 1 0 35328 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_384
timestamp 1649977179
transform 1 0 36432 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1649977179
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1649977179
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_421
timestamp 1649977179
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_433
timestamp 1649977179
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1649977179
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1649977179
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1649977179
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_480
timestamp 1649977179
transform 1 0 45264 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_492
timestamp 1649977179
transform 1 0 46368 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1649977179
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1649977179
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_533
timestamp 1649977179
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_545
timestamp 1649977179
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1649977179
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1649977179
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1649977179
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_592
timestamp 1649977179
transform 1 0 55568 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_604
timestamp 1649977179
transform 1 0 56672 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_629
timestamp 1649977179
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_641
timestamp 1649977179
transform 1 0 60076 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_645
timestamp 1649977179
transform 1 0 60444 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_657
timestamp 1649977179
transform 1 0 61548 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_669
timestamp 1649977179
transform 1 0 62652 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_673
timestamp 1649977179
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_685
timestamp 1649977179
transform 1 0 64124 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_696
timestamp 1649977179
transform 1 0 65136 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_701
timestamp 1649977179
transform 1 0 65596 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_713
timestamp 1649977179
transform 1 0 66700 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_717
timestamp 1649977179
transform 1 0 67068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_724
timestamp 1649977179
transform 1 0 67712 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1649977179
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1649977179
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1649977179
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1649977179
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1649977179
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1649977179
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1649977179
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1649977179
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1649977179
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1649977179
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1649977179
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1649977179
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1649977179
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1649977179
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1649977179
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1649977179
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1649977179
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1649977179
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1649977179
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1649977179
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1649977179
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1649977179
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1649977179
transform 1 0 60352 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1649977179
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1649977179
transform 1 0 65504 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1649977179
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0791_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0792_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0793_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11868 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0794_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0795_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0796_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10856 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0797_
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0798_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10764 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0799_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0800_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0801_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8004 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0802_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0803_
timestamp 1649977179
transform -1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0804_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1649977179
transform -1 0 2484 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0806_
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0809_
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 1649977179
transform -1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0812_
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 1649977179
transform -1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1649977179
transform 1 0 4140 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0816_
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0817_
timestamp 1649977179
transform 1 0 5520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1649977179
transform 1 0 7176 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0819_
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 1649977179
transform -1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0821_
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0823_
timestamp 1649977179
transform 1 0 20148 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1649977179
transform -1 0 21252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1649977179
transform -1 0 21344 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0826_
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0827_
timestamp 1649977179
transform -1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0829_
timestamp 1649977179
transform -1 0 8372 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0830_
timestamp 1649977179
transform -1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0832_
timestamp 1649977179
transform -1 0 17756 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0833_
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0834_
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0835_
timestamp 1649977179
transform -1 0 8096 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0837_
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0838_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0839_
timestamp 1649977179
transform -1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_4  _0840_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12788 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0841_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13432 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0842_
timestamp 1649977179
transform -1 0 11224 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0843_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0844_
timestamp 1649977179
transform -1 0 3312 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1649977179
transform -1 0 5888 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 1649977179
transform 1 0 1748 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0847_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0848_
timestamp 1649977179
transform -1 0 8280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0849_
timestamp 1649977179
transform -1 0 2668 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0850_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3312 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0851_
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1649977179
transform 1 0 2208 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0853_
timestamp 1649977179
transform -1 0 3036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0854_
timestamp 1649977179
transform 1 0 1564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0855_
timestamp 1649977179
transform 1 0 1932 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0856_
timestamp 1649977179
transform -1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0857_
timestamp 1649977179
transform 1 0 4140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0858_
timestamp 1649977179
transform 1 0 1748 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0859_
timestamp 1649977179
transform -1 0 3312 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0860_
timestamp 1649977179
transform 1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0861_
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0862_
timestamp 1649977179
transform -1 0 3312 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0864_
timestamp 1649977179
transform 1 0 2668 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 1649977179
transform 1 0 2668 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1649977179
transform 1 0 2116 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0867_
timestamp 1649977179
transform -1 0 2668 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0868_
timestamp 1649977179
transform -1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0869_
timestamp 1649977179
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1649977179
transform -1 0 2668 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0871_
timestamp 1649977179
transform -1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0872_
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1649977179
transform -1 0 1840 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0874_
timestamp 1649977179
transform -1 0 2300 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0875_
timestamp 1649977179
transform 1 0 15364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 1649977179
transform 1 0 1840 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0877_
timestamp 1649977179
transform -1 0 2760 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0878_
timestamp 1649977179
transform -1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0880_
timestamp 1649977179
transform -1 0 3036 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0881_
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0883_
timestamp 1649977179
transform -1 0 2668 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0884_
timestamp 1649977179
transform -1 0 3864 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0885_
timestamp 1649977179
transform -1 0 12512 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0886_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0887_
timestamp 1649977179
transform 1 0 9568 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0888_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0890_
timestamp 1649977179
transform -1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1649977179
transform -1 0 2760 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0892_
timestamp 1649977179
transform 1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0893_
timestamp 1649977179
transform 1 0 1472 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0894_
timestamp 1649977179
transform -1 0 3036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1649977179
transform 1 0 1932 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0896_
timestamp 1649977179
transform -1 0 2852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0897_
timestamp 1649977179
transform -1 0 3220 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0898_
timestamp 1649977179
transform -1 0 2668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0899_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0900_
timestamp 1649977179
transform -1 0 3312 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 1649977179
transform 1 0 1564 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0902_
timestamp 1649977179
transform -1 0 2668 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0903_
timestamp 1649977179
transform -1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0904_
timestamp 1649977179
transform 1 0 2392 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1649977179
transform -1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1649977179
transform 1 0 1656 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0907_
timestamp 1649977179
transform -1 0 2760 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0909_
timestamp 1649977179
transform -1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0910_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0911_
timestamp 1649977179
transform -1 0 3036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1649977179
transform 1 0 1564 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0913_
timestamp 1649977179
transform -1 0 3128 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0914_
timestamp 1649977179
transform -1 0 3588 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0915_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0916_
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0917_
timestamp 1649977179
transform 1 0 7176 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0918_
timestamp 1649977179
transform -1 0 3312 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1649977179
transform 1 0 2668 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0920_
timestamp 1649977179
transform -1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0921_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0922_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10212 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0923_
timestamp 1649977179
transform 1 0 8924 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0924_
timestamp 1649977179
transform -1 0 9200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0925_
timestamp 1649977179
transform -1 0 8280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0926_
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1649977179
transform -1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1649977179
transform -1 0 6440 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0929_
timestamp 1649977179
transform -1 0 4416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0930_
timestamp 1649977179
transform -1 0 6900 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0931_
timestamp 1649977179
transform -1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1649977179
transform -1 0 8280 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0933_
timestamp 1649977179
transform -1 0 8004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0935_
timestamp 1649977179
transform -1 0 9844 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0936_
timestamp 1649977179
transform -1 0 11040 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1649977179
transform 1 0 8648 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0938_
timestamp 1649977179
transform -1 0 11040 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0939_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0940_
timestamp 1649977179
transform -1 0 8096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1649977179
transform -1 0 9752 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0942_
timestamp 1649977179
transform -1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0944_
timestamp 1649977179
transform 1 0 8832 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0945_
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0946_
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0947_
timestamp 1649977179
transform -1 0 6900 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0948_
timestamp 1649977179
transform -1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0949_
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1649977179
transform -1 0 7360 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0952_
timestamp 1649977179
transform -1 0 8464 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0953_
timestamp 1649977179
transform -1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1649977179
transform -1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1649977179
transform -1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1649977179
transform -1 0 12144 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 1649977179
transform -1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _0958_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15364 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0959_
timestamp 1649977179
transform -1 0 15456 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0960_
timestamp 1649977179
transform -1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0961_
timestamp 1649977179
transform -1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0962_
timestamp 1649977179
transform -1 0 8004 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1649977179
transform -1 0 9384 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0965_
timestamp 1649977179
transform 1 0 6440 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0966_
timestamp 1649977179
transform 1 0 6532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1649977179
transform -1 0 5888 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0968_
timestamp 1649977179
transform 1 0 6532 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1649977179
transform 1 0 7728 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0970_
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0971_
timestamp 1649977179
transform -1 0 8464 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0972_
timestamp 1649977179
transform -1 0 7176 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0973_
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0974_
timestamp 1649977179
transform 1 0 6532 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0975_
timestamp 1649977179
transform 1 0 6348 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0976_
timestamp 1649977179
transform -1 0 7544 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1649977179
transform -1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0978_
timestamp 1649977179
transform -1 0 7268 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0979_
timestamp 1649977179
transform -1 0 8188 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1649977179
transform -1 0 7268 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0981_
timestamp 1649977179
transform 1 0 6164 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0982_
timestamp 1649977179
transform 1 0 10212 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0983_
timestamp 1649977179
transform 1 0 7544 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0984_
timestamp 1649977179
transform -1 0 11776 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0985_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0986_
timestamp 1649977179
transform -1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1649977179
transform -1 0 10764 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0988_
timestamp 1649977179
transform -1 0 10856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0989_
timestamp 1649977179
transform -1 0 7728 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0990_
timestamp 1649977179
transform 1 0 6440 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0991_
timestamp 1649977179
transform 1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0992_
timestamp 1649977179
transform 1 0 20424 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0993_
timestamp 1649977179
transform -1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0994_
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0995_
timestamp 1649977179
transform 1 0 14536 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0996_
timestamp 1649977179
transform -1 0 15548 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1649977179
transform -1 0 9384 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0999_
timestamp 1649977179
transform 1 0 9108 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1000_
timestamp 1649977179
transform 1 0 19504 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1001_
timestamp 1649977179
transform -1 0 16928 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1002_
timestamp 1649977179
transform 1 0 9016 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1649977179
transform 1 0 14352 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 1649977179
transform -1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1006_
timestamp 1649977179
transform -1 0 17020 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1007_
timestamp 1649977179
transform -1 0 15640 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1008_
timestamp 1649977179
transform -1 0 15364 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1009_
timestamp 1649977179
transform 1 0 12696 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1649977179
transform -1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1011_
timestamp 1649977179
transform -1 0 16192 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1012_
timestamp 1649977179
transform -1 0 16192 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 1649977179
transform 1 0 17020 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1014_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1015_
timestamp 1649977179
transform -1 0 17756 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1649977179
transform -1 0 18032 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1019_
timestamp 1649977179
transform -1 0 17664 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1649977179
transform -1 0 15916 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1021_
timestamp 1649977179
transform -1 0 14260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1022_
timestamp 1649977179
transform -1 0 15456 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1023_
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1024_
timestamp 1649977179
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1025_
timestamp 1649977179
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1026_
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1027_
timestamp 1649977179
transform -1 0 23368 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1028_
timestamp 1649977179
transform -1 0 24012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1029_
timestamp 1649977179
transform 1 0 24656 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1649977179
transform 1 0 22816 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1032_
timestamp 1649977179
transform -1 0 23368 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1033_
timestamp 1649977179
transform 1 0 24840 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1034_
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1035_
timestamp 1649977179
transform 1 0 19688 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1649977179
transform -1 0 24472 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1037_
timestamp 1649977179
transform 1 0 23184 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1038_
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1039_
timestamp 1649977179
transform 1 0 24564 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1040_
timestamp 1649977179
transform -1 0 25760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1041_
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1649977179
transform -1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1044_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1045_
timestamp 1649977179
transform 1 0 26128 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1046_
timestamp 1649977179
transform -1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1047_
timestamp 1649977179
transform 1 0 28060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1048_
timestamp 1649977179
transform 1 0 24656 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1649977179
transform -1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1649977179
transform 1 0 27508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1051_
timestamp 1649977179
transform 1 0 24932 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1052_
timestamp 1649977179
transform -1 0 28336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1053_
timestamp 1649977179
transform 1 0 28888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1649977179
transform 1 0 27232 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1055_
timestamp 1649977179
transform -1 0 28796 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1056_
timestamp 1649977179
transform 1 0 27324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1649977179
transform 1 0 27416 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1058_
timestamp 1649977179
transform 1 0 27508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1059_
timestamp 1649977179
transform 1 0 26036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1060_
timestamp 1649977179
transform 1 0 26036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1061_
timestamp 1649977179
transform 1 0 25760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1649977179
transform 1 0 24656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1649977179
transform 1 0 24196 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1064_
timestamp 1649977179
transform 1 0 24656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1065_
timestamp 1649977179
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1649977179
transform 1 0 23276 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1067_
timestamp 1649977179
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1068_
timestamp 1649977179
transform 1 0 23184 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1069_
timestamp 1649977179
transform -1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1070_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16100 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1649977179
transform -1 0 25300 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1649977179
transform 1 0 26220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1073_
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1074_
timestamp 1649977179
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1075_
timestamp 1649977179
transform 1 0 25668 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1649977179
transform -1 0 31096 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 1649977179
transform 1 0 30544 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1078_
timestamp 1649977179
transform 1 0 30636 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1649977179
transform -1 0 32568 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1080_
timestamp 1649977179
transform -1 0 32568 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1649977179
transform 1 0 32292 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1649977179
transform -1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1649977179
transform -1 0 33304 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1649977179
transform 1 0 30268 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1086_
timestamp 1649977179
transform 1 0 28428 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1649977179
transform -1 0 30636 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1088_
timestamp 1649977179
transform -1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1089_
timestamp 1649977179
transform 1 0 28520 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1649977179
transform 1 0 26680 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1649977179
transform -1 0 27876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1093_
timestamp 1649977179
transform 1 0 29716 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1094_
timestamp 1649977179
transform -1 0 30820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1095_
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1096_
timestamp 1649977179
transform -1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1097_
timestamp 1649977179
transform 1 0 26772 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1098_
timestamp 1649977179
transform -1 0 28336 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1649977179
transform 1 0 26312 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1100_
timestamp 1649977179
transform -1 0 34316 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1649977179
transform 1 0 25760 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1103_
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _1104_
timestamp 1649977179
transform -1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1105_
timestamp 1649977179
transform 1 0 19320 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1106_
timestamp 1649977179
transform 1 0 32936 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1107_
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1108_
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1109_
timestamp 1649977179
transform 1 0 31188 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1110_
timestamp 1649977179
transform 1 0 34132 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1649977179
transform -1 0 35144 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1649977179
transform -1 0 35420 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1113_
timestamp 1649977179
transform 1 0 35236 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1649977179
transform 1 0 35880 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1115_
timestamp 1649977179
transform 1 0 39744 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1116_
timestamp 1649977179
transform -1 0 40572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1117_
timestamp 1649977179
transform 1 0 39836 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1649977179
transform -1 0 39192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1119_
timestamp 1649977179
transform -1 0 40756 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1120_
timestamp 1649977179
transform 1 0 34868 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1649977179
transform -1 0 36524 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1122_
timestamp 1649977179
transform -1 0 35328 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1123_
timestamp 1649977179
transform -1 0 34040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1124_
timestamp 1649977179
transform 1 0 38732 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1125_
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1649977179
transform -1 0 38548 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1127_
timestamp 1649977179
transform -1 0 36708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1649977179
transform -1 0 37720 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1129_
timestamp 1649977179
transform 1 0 35236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1649977179
transform 1 0 33488 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1131_
timestamp 1649977179
transform -1 0 34316 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1132_
timestamp 1649977179
transform -1 0 35420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1133_
timestamp 1649977179
transform 1 0 33764 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1134_
timestamp 1649977179
transform 1 0 33488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1649977179
transform 1 0 33580 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1649977179
transform 1 0 33488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1137_
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1138_
timestamp 1649977179
transform 1 0 32752 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1139_
timestamp 1649977179
transform -1 0 32384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1649977179
transform 1 0 35512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1141_
timestamp 1649977179
transform 1 0 33120 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1142_
timestamp 1649977179
transform -1 0 34224 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1649977179
transform 1 0 33396 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1144_
timestamp 1649977179
transform 1 0 33488 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1649977179
transform -1 0 33028 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1146_
timestamp 1649977179
transform -1 0 35420 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1148_
timestamp 1649977179
transform 1 0 39560 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1649977179
transform 1 0 39192 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1151_
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1649977179
transform 1 0 38916 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1153_
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1154_
timestamp 1649977179
transform -1 0 35696 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1649977179
transform -1 0 34224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1156_
timestamp 1649977179
transform 1 0 35512 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1157_
timestamp 1649977179
transform -1 0 36892 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1158_
timestamp 1649977179
transform 1 0 35328 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1159_
timestamp 1649977179
transform -1 0 36616 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1160_
timestamp 1649977179
transform -1 0 32844 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1161_
timestamp 1649977179
transform 1 0 28152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1162_
timestamp 1649977179
transform 1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1163_
timestamp 1649977179
transform -1 0 33028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1164_
timestamp 1649977179
transform -1 0 31188 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1165_
timestamp 1649977179
transform 1 0 30544 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1166_
timestamp 1649977179
transform 1 0 31372 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1649977179
transform 1 0 31372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1168_
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1169_
timestamp 1649977179
transform -1 0 34960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1170_
timestamp 1649977179
transform 1 0 21988 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1171_
timestamp 1649977179
transform 1 0 30728 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1172_
timestamp 1649977179
transform 1 0 32200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1649977179
transform 1 0 34776 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1174_
timestamp 1649977179
transform 1 0 32292 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1649977179
transform -1 0 34960 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1649977179
transform -1 0 34224 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1177_
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1178_
timestamp 1649977179
transform 1 0 36064 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1179_
timestamp 1649977179
transform 1 0 35880 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1180_
timestamp 1649977179
transform 1 0 35880 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1181_
timestamp 1649977179
transform 1 0 35052 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1649977179
transform -1 0 36708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1649977179
transform 1 0 36064 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1184_
timestamp 1649977179
transform -1 0 37904 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1186_
timestamp 1649977179
transform 1 0 38088 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1187_
timestamp 1649977179
transform 1 0 34776 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1649977179
transform 1 0 34132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1649977179
transform 1 0 38456 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1190_
timestamp 1649977179
transform 1 0 38180 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1191_
timestamp 1649977179
transform -1 0 37720 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1192_
timestamp 1649977179
transform 1 0 35880 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1193_
timestamp 1649977179
transform -1 0 36616 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1195_
timestamp 1649977179
transform 1 0 36064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1649977179
transform -1 0 34224 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1649977179
transform 1 0 34132 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1649977179
transform -1 0 36616 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1199_
timestamp 1649977179
transform -1 0 35972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1649977179
transform 1 0 32844 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1201_
timestamp 1649977179
transform 1 0 33396 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1202_
timestamp 1649977179
transform 1 0 22080 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1203_
timestamp 1649977179
transform -1 0 23644 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _1204_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1205_
timestamp 1649977179
transform -1 0 21344 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1206_
timestamp 1649977179
transform 1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1207_
timestamp 1649977179
transform 1 0 21988 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1208_
timestamp 1649977179
transform 1 0 20700 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1649977179
transform -1 0 22264 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1210_
timestamp 1649977179
transform -1 0 20700 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1211_
timestamp 1649977179
transform -1 0 25300 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1212_
timestamp 1649977179
transform 1 0 20240 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1213_
timestamp 1649977179
transform -1 0 20700 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1214_
timestamp 1649977179
transform 1 0 20608 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1215_
timestamp 1649977179
transform 1 0 20608 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1216_
timestamp 1649977179
transform -1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1217_
timestamp 1649977179
transform -1 0 22724 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1218_
timestamp 1649977179
transform -1 0 21896 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1219_
timestamp 1649977179
transform -1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1649977179
transform 1 0 23644 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1221_
timestamp 1649977179
transform 1 0 23184 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1222_
timestamp 1649977179
transform -1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1649977179
transform 1 0 23276 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1224_
timestamp 1649977179
transform -1 0 24840 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1225_
timestamp 1649977179
transform -1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1226_
timestamp 1649977179
transform -1 0 22908 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1649977179
transform -1 0 21344 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1649977179
transform 1 0 23460 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1229_
timestamp 1649977179
transform -1 0 25852 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1230_
timestamp 1649977179
transform -1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1231_
timestamp 1649977179
transform 1 0 19504 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1649977179
transform 1 0 25024 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1649977179
transform -1 0 27692 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1234_
timestamp 1649977179
transform -1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1649977179
transform 1 0 24840 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1236_
timestamp 1649977179
transform -1 0 25944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1237_
timestamp 1649977179
transform -1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1238_
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1649977179
transform -1 0 24472 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1240_
timestamp 1649977179
transform -1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1241_
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1242_
timestamp 1649977179
transform -1 0 23092 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1243_
timestamp 1649977179
transform -1 0 18952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1244_
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1245_
timestamp 1649977179
transform 1 0 19688 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1246_
timestamp 1649977179
transform 1 0 27784 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1247_
timestamp 1649977179
transform 1 0 22172 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _1248_
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1249_
timestamp 1649977179
transform 1 0 17572 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1250_
timestamp 1649977179
transform -1 0 30268 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1251_
timestamp 1649977179
transform -1 0 29072 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1252_
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1253_
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1649977179
transform -1 0 31188 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1649977179
transform -1 0 29164 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1257_
timestamp 1649977179
transform 1 0 28244 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1649977179
transform 1 0 28980 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1649977179
transform -1 0 29440 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1260_
timestamp 1649977179
transform -1 0 30912 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1261_
timestamp 1649977179
transform -1 0 31004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1262_
timestamp 1649977179
transform 1 0 29992 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1263_
timestamp 1649977179
transform -1 0 30820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1264_
timestamp 1649977179
transform 1 0 31096 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1265_
timestamp 1649977179
transform 1 0 27968 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1266_
timestamp 1649977179
transform -1 0 31372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1267_
timestamp 1649977179
transform 1 0 29532 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1268_
timestamp 1649977179
transform -1 0 30544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1269_
timestamp 1649977179
transform 1 0 32384 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1270_
timestamp 1649977179
transform -1 0 33212 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1271_
timestamp 1649977179
transform 1 0 32752 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1272_
timestamp 1649977179
transform -1 0 33764 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1649977179
transform 1 0 33304 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1649977179
transform -1 0 33120 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1649977179
transform 1 0 31188 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1649977179
transform -1 0 32936 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1277_
timestamp 1649977179
transform -1 0 31740 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1278_
timestamp 1649977179
transform 1 0 21160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1279_
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1280_
timestamp 1649977179
transform 1 0 31372 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1281_
timestamp 1649977179
transform -1 0 29072 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1282_
timestamp 1649977179
transform -1 0 14628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1283_
timestamp 1649977179
transform 1 0 14720 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1284_
timestamp 1649977179
transform 1 0 16008 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1285_
timestamp 1649977179
transform -1 0 16560 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1286_
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1649977179
transform -1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1288_
timestamp 1649977179
transform 1 0 14996 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1289_
timestamp 1649977179
transform 1 0 14904 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1290_
timestamp 1649977179
transform 1 0 17112 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1291_
timestamp 1649977179
transform -1 0 17756 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1292_
timestamp 1649977179
transform 1 0 15272 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1293_
timestamp 1649977179
transform -1 0 16744 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1649977179
transform 1 0 15364 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1295_
timestamp 1649977179
transform -1 0 18584 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1296_
timestamp 1649977179
transform 1 0 16192 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1297_
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1298_
timestamp 1649977179
transform -1 0 17940 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1299_
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1300_
timestamp 1649977179
transform -1 0 16192 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1301_
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1302_
timestamp 1649977179
transform -1 0 18768 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1303_
timestamp 1649977179
transform 1 0 17572 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1304_
timestamp 1649977179
transform -1 0 18676 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1305_
timestamp 1649977179
transform 1 0 18216 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1306_
timestamp 1649977179
transform -1 0 19964 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1307_
timestamp 1649977179
transform 1 0 16928 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1308_
timestamp 1649977179
transform -1 0 17664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1309_
timestamp 1649977179
transform 1 0 17112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1649977179
transform -1 0 18584 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1649977179
transform -1 0 17756 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1649977179
transform 1 0 15732 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1313_
timestamp 1649977179
transform -1 0 16744 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1314_
timestamp 1649977179
transform 1 0 13064 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1315_
timestamp 1649977179
transform 1 0 13524 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1316_
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1317_
timestamp 1649977179
transform -1 0 13616 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1649977179
transform 1 0 12512 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 1649977179
transform 1 0 12512 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1320_
timestamp 1649977179
transform -1 0 8464 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1321_
timestamp 1649977179
transform 1 0 9108 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1649977179
transform 1 0 11316 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1324_
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1325_
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1326_
timestamp 1649977179
transform -1 0 11776 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1327_
timestamp 1649977179
transform 1 0 8924 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1329_
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1330_
timestamp 1649977179
transform 1 0 12052 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1331_
timestamp 1649977179
transform -1 0 13616 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1332_
timestamp 1649977179
transform -1 0 14260 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1333_
timestamp 1649977179
transform -1 0 13432 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1335_
timestamp 1649977179
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1336_
timestamp 1649977179
transform -1 0 9844 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1337_
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1338_
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1339_
timestamp 1649977179
transform -1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1340_
timestamp 1649977179
transform -1 0 14904 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1649977179
transform 1 0 13156 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1649977179
transform -1 0 14076 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1343_
timestamp 1649977179
transform 1 0 12788 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1344_
timestamp 1649977179
transform 1 0 13248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1345_
timestamp 1649977179
transform 1 0 13156 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1346_
timestamp 1649977179
transform -1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1347_
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1348_
timestamp 1649977179
transform -1 0 23368 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1349_
timestamp 1649977179
transform -1 0 23552 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1350_
timestamp 1649977179
transform 1 0 23276 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1351_
timestamp 1649977179
transform 1 0 21528 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1352_
timestamp 1649977179
transform -1 0 21988 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1649977179
transform -1 0 24840 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1649977179
transform 1 0 23184 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1649977179
transform -1 0 24012 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1356_
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1357_
timestamp 1649977179
transform -1 0 23920 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1358_
timestamp 1649977179
transform 1 0 25760 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1359_
timestamp 1649977179
transform -1 0 27692 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1649977179
transform 1 0 26220 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1361_
timestamp 1649977179
transform -1 0 26496 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1362_
timestamp 1649977179
transform 1 0 25208 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1363_
timestamp 1649977179
transform 1 0 25208 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1364_
timestamp 1649977179
transform -1 0 23552 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1365_
timestamp 1649977179
transform -1 0 23000 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1649977179
transform -1 0 26496 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1367_
timestamp 1649977179
transform -1 0 25944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1649977179
transform 1 0 27876 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1369_
timestamp 1649977179
transform 1 0 21804 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1370_
timestamp 1649977179
transform -1 0 28888 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1371_
timestamp 1649977179
transform 1 0 27968 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1372_
timestamp 1649977179
transform -1 0 29072 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1373_
timestamp 1649977179
transform -1 0 23368 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1374_
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1375_
timestamp 1649977179
transform -1 0 20240 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1376_
timestamp 1649977179
transform 1 0 20608 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1377_
timestamp 1649977179
transform 1 0 23368 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1378_
timestamp 1649977179
transform -1 0 22816 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1379_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1649977179
transform -1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1382_
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1383_
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1384_
timestamp 1649977179
transform 1 0 19412 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1385_
timestamp 1649977179
transform 1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1386_
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1387_
timestamp 1649977179
transform -1 0 18768 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1388_
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1649977179
transform -1 0 19688 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1390_
timestamp 1649977179
transform 1 0 17572 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1391_
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1392_
timestamp 1649977179
transform -1 0 20516 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1393_
timestamp 1649977179
transform 1 0 19688 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1394_
timestamp 1649977179
transform -1 0 20516 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1395_
timestamp 1649977179
transform -1 0 17664 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1396_
timestamp 1649977179
transform -1 0 18768 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1397_
timestamp 1649977179
transform 1 0 22908 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1398_
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1399_
timestamp 1649977179
transform -1 0 28520 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1400_
timestamp 1649977179
transform 1 0 23644 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1649977179
transform -1 0 28704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1649977179
transform 1 0 28244 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1403_
timestamp 1649977179
transform -1 0 29072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1649977179
transform 1 0 26036 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1405_
timestamp 1649977179
transform -1 0 27692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1406_
timestamp 1649977179
transform -1 0 26680 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1407_
timestamp 1649977179
transform 1 0 25208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1408_
timestamp 1649977179
transform -1 0 25944 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1409_
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1410_
timestamp 1649977179
transform -1 0 21252 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1411_
timestamp 1649977179
transform 1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1412_
timestamp 1649977179
transform -1 0 20884 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1649977179
transform -1 0 21528 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1414_
timestamp 1649977179
transform -1 0 21344 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1415_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14904 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1416_
timestamp 1649977179
transform -1 0 13524 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1417_
timestamp 1649977179
transform -1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1418_
timestamp 1649977179
transform -1 0 11132 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1419_
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1420_
timestamp 1649977179
transform -1 0 13892 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _1421_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1422_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1423_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1424_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33488 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1425_
timestamp 1649977179
transform -1 0 30176 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1426_
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1428_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1429_
timestamp 1649977179
transform 1 0 8924 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1430_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1431_
timestamp 1649977179
transform 1 0 20240 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1432_
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1433_
timestamp 1649977179
transform -1 0 13064 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1434_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1435_
timestamp 1649977179
transform -1 0 33488 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1436_
timestamp 1649977179
transform -1 0 30176 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1437_
timestamp 1649977179
transform 1 0 20792 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1438_
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1439_
timestamp 1649977179
transform -1 0 21344 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1440_
timestamp 1649977179
transform 1 0 10120 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 1649977179
transform 1 0 11592 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1442_
timestamp 1649977179
transform -1 0 19964 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1443_
timestamp 1649977179
transform 1 0 24288 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1444_
timestamp 1649977179
transform -1 0 20332 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1445_
timestamp 1649977179
transform -1 0 9752 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1447_
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1448_
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1649977179
transform -1 0 33580 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1450_
timestamp 1649977179
transform -1 0 30268 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1451_
timestamp 1649977179
transform 1 0 20148 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1452_
timestamp 1649977179
transform 1 0 25484 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1453_
timestamp 1649977179
transform 1 0 23736 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1454_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1455_
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1649977179
transform 1 0 7820 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1457_
timestamp 1649977179
transform 1 0 12144 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1458_
timestamp 1649977179
transform 1 0 20332 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1459_
timestamp 1649977179
transform -1 0 25760 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1460_
timestamp 1649977179
transform -1 0 14536 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1461_
timestamp 1649977179
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1462_
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1463_
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1464_
timestamp 1649977179
transform -1 0 32200 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1465_
timestamp 1649977179
transform -1 0 31648 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1466_
timestamp 1649977179
transform -1 0 31740 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1467_
timestamp 1649977179
transform 1 0 30728 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1468_
timestamp 1649977179
transform 1 0 30084 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1469_
timestamp 1649977179
transform -1 0 30360 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1470_
timestamp 1649977179
transform 1 0 25944 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1471_
timestamp 1649977179
transform 1 0 28428 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1472_
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1473_
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1474_
timestamp 1649977179
transform 1 0 11592 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1475_
timestamp 1649977179
transform 1 0 29808 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1476_
timestamp 1649977179
transform -1 0 11040 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1477_
timestamp 1649977179
transform -1 0 13064 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1478_
timestamp 1649977179
transform 1 0 10304 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1479_
timestamp 1649977179
transform 1 0 10856 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1480_
timestamp 1649977179
transform 1 0 21988 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1481_
timestamp 1649977179
transform 1 0 23000 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1482_
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1483_
timestamp 1649977179
transform -1 0 25668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1484_
timestamp 1649977179
transform -1 0 13248 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1485_
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1486_
timestamp 1649977179
transform 1 0 12696 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1487_
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1488_
timestamp 1649977179
transform -1 0 32752 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1489_
timestamp 1649977179
transform -1 0 32752 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1490_
timestamp 1649977179
transform 1 0 28428 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1491_
timestamp 1649977179
transform 1 0 11776 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1492_
timestamp 1649977179
transform 1 0 29532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1493_
timestamp 1649977179
transform -1 0 13616 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1649977179
transform 1 0 14628 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1495_
timestamp 1649977179
transform 1 0 10212 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1496_
timestamp 1649977179
transform 1 0 11868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1497_
timestamp 1649977179
transform 1 0 22816 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1498_
timestamp 1649977179
transform 1 0 22448 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1499_
timestamp 1649977179
transform 1 0 23276 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1500_
timestamp 1649977179
transform 1 0 25852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1501_
timestamp 1649977179
transform -1 0 14628 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1502_
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1503_
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1504_
timestamp 1649977179
transform -1 0 32752 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp 1649977179
transform -1 0 30452 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1506_
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1507_
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1508_
timestamp 1649977179
transform -1 0 30176 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1509_
timestamp 1649977179
transform 1 0 10212 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1510_
timestamp 1649977179
transform 1 0 11868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1511_
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1512_
timestamp 1649977179
transform -1 0 26496 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1513_
timestamp 1649977179
transform -1 0 16652 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1514_
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1515_
timestamp 1649977179
transform -1 0 15916 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1516_
timestamp 1649977179
transform -1 0 31648 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1517_
timestamp 1649977179
transform -1 0 31648 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1518_
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1519_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1520_
timestamp 1649977179
transform 1 0 29532 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1521_
timestamp 1649977179
transform 1 0 9936 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1522_
timestamp 1649977179
transform 1 0 11592 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1523_
timestamp 1649977179
transform 1 0 23736 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1524_
timestamp 1649977179
transform -1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1525_
timestamp 1649977179
transform -1 0 17388 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1526_
timestamp 1649977179
transform 1 0 13432 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1527_
timestamp 1649977179
transform -1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1528_
timestamp 1649977179
transform -1 0 18768 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1529_
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1530_
timestamp 1649977179
transform -1 0 32016 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1531_
timestamp 1649977179
transform -1 0 32292 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1649977179
transform 1 0 25576 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1534_
timestamp 1649977179
transform 1 0 27232 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1535_
timestamp 1649977179
transform -1 0 11040 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1536_
timestamp 1649977179
transform 1 0 15916 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1537_
timestamp 1649977179
transform 1 0 24748 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1538_
timestamp 1649977179
transform -1 0 26220 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1539_
timestamp 1649977179
transform -1 0 19044 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1540_
timestamp 1649977179
transform -1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1541_
timestamp 1649977179
transform 1 0 17940 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1542_
timestamp 1649977179
transform -1 0 32108 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1649977179
transform -1 0 31464 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1649977179
transform -1 0 26312 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1546_
timestamp 1649977179
transform -1 0 26036 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1649977179
transform 1 0 13156 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1548_
timestamp 1649977179
transform 1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1549_
timestamp 1649977179
transform 1 0 20700 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1550_
timestamp 1649977179
transform -1 0 22448 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1649977179
transform -1 0 16744 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1552_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1553_
timestamp 1649977179
transform 1 0 15088 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1554_
timestamp 1649977179
transform -1 0 32752 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1555_
timestamp 1649977179
transform -1 0 31648 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1556_
timestamp 1649977179
transform -1 0 25024 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1557_
timestamp 1649977179
transform 1 0 10028 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1558_
timestamp 1649977179
transform -1 0 25116 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1559_
timestamp 1649977179
transform 1 0 12328 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1560_
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1561_
timestamp 1649977179
transform -1 0 20056 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1562_
timestamp 1649977179
transform -1 0 20424 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1563_
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1564_
timestamp 1649977179
transform 1 0 17204 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1565_
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1566_
timestamp 1649977179
transform -1 0 33120 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1567_
timestamp 1649977179
transform -1 0 31372 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1568_
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1569_
timestamp 1649977179
transform 1 0 10304 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1570_
timestamp 1649977179
transform 1 0 22080 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1571_
timestamp 1649977179
transform 1 0 12972 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1572_
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1573_
timestamp 1649977179
transform 1 0 20424 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1574_
timestamp 1649977179
transform -1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1575_
timestamp 1649977179
transform -1 0 15640 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1576_
timestamp 1649977179
transform -1 0 15456 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1577_
timestamp 1649977179
transform 1 0 14536 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1578_
timestamp 1649977179
transform 1 0 20056 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1579_
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1580_
timestamp 1649977179
transform -1 0 10120 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1581_
timestamp 1649977179
transform -1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1582_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5704 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1649977179
transform -1 0 5244 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1649977179
transform -1 0 23276 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1649977179
transform -1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1649977179
transform 1 0 5336 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1649977179
transform 1 0 4048 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1649977179
transform 1 0 3404 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1649977179
transform 1 0 4324 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1649977179
transform 1 0 3772 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1649977179
transform 1 0 4232 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1649977179
transform 1 0 3128 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1649977179
transform -1 0 4048 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1649977179
transform 1 0 4968 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1649977179
transform 1 0 5336 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1649977179
transform 1 0 3864 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1649977179
transform 1 0 3404 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1649977179
transform -1 0 4048 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1649977179
transform 1 0 3772 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1649977179
transform 1 0 4968 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1649977179
transform 1 0 7728 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1649977179
transform 1 0 10948 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1649977179
transform -1 0 12972 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1649977179
transform 1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1649977179
transform -1 0 6716 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1649977179
transform 1 0 6808 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1649977179
transform 1 0 7360 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1649977179
transform 1 0 7912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1649977179
transform 1 0 12788 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1649977179
transform 1 0 11592 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1649977179
transform 1 0 8924 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1649977179
transform 1 0 6716 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1649977179
transform 1 0 9200 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1649977179
transform -1 0 18124 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1649977179
transform 1 0 17664 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1649977179
transform 1 0 15732 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1649977179
transform 1 0 17296 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1649977179
transform 1 0 18584 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1649977179
transform 1 0 17848 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1649977179
transform 1 0 13156 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1649977179
transform 1 0 18584 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1649977179
transform 1 0 22724 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1649977179
transform -1 0 26864 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1649977179
transform 1 0 27508 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1649977179
transform 1 0 26956 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1649977179
transform -1 0 30820 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1649977179
transform -1 0 28704 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1649977179
transform 1 0 25392 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1649977179
transform 1 0 22448 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1649977179
transform -1 0 23920 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1649977179
transform -1 0 31832 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1649977179
transform -1 0 34960 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1649977179
transform -1 0 36340 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1649977179
transform -1 0 34592 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1649977179
transform -1 0 32568 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1649977179
transform 1 0 27508 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1649977179
transform -1 0 33028 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1649977179
transform -1 0 28704 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1649977179
transform 1 0 28152 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1649977179
transform -1 0 26220 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1649977179
transform -1 0 25852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1649977179
transform -1 0 37168 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1649977179
transform -1 0 37168 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1649977179
transform -1 0 39192 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1649977179
transform -1 0 37168 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1649977179
transform 1 0 37352 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1649977179
transform 1 0 37260 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1649977179
transform 1 0 35420 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1649977179
transform -1 0 33580 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1649977179
transform -1 0 35236 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1649977179
transform -1 0 36708 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1649977179
transform -1 0 32384 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1649977179
transform -1 0 36156 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1649977179
transform -1 0 39008 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1649977179
transform -1 0 39008 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1649977179
transform -1 0 39008 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1687_
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1649977179
transform -1 0 33856 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1649977179
transform -1 0 31648 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1649977179
transform -1 0 36800 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1649977179
transform -1 0 35052 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1649977179
transform -1 0 37628 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1649977179
transform 1 0 37444 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1649977179
transform 1 0 37628 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1649977179
transform 1 0 37720 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1649977179
transform -1 0 39192 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1649977179
transform 1 0 35880 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1649977179
transform -1 0 33764 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1649977179
transform -1 0 39008 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1649977179
transform -1 0 32292 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1649977179
transform 1 0 19320 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1649977179
transform -1 0 21160 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1649977179
transform 1 0 23184 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1649977179
transform -1 0 26496 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1649977179
transform -1 0 28244 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1649977179
transform -1 0 27876 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1649977179
transform 1 0 26956 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1649977179
transform 1 0 25576 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1649977179
transform -1 0 24288 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1649977179
transform -1 0 22448 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1649977179
transform 1 0 28152 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1649977179
transform -1 0 31188 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1649977179
transform -1 0 33580 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1649977179
transform -1 0 33580 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1649977179
transform -1 0 33212 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1649977179
transform 1 0 35420 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1649977179
transform 1 0 34684 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1649977179
transform -1 0 34960 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1649977179
transform 1 0 35328 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1649977179
transform 1 0 29256 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1649977179
transform 1 0 13616 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1649977179
transform -1 0 18952 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1649977179
transform -1 0 18768 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1649977179
transform -1 0 16652 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1649977179
transform -1 0 18768 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1649977179
transform 1 0 19228 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1649977179
transform 1 0 19320 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1649977179
transform -1 0 16192 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1649977179
transform -1 0 19596 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1649977179
transform -1 0 18676 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1649977179
transform 1 0 6808 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1649977179
transform -1 0 11868 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1649977179
transform 1 0 4416 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1649977179
transform -1 0 10948 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1649977179
transform -1 0 14076 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1649977179
transform 1 0 8188 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1649977179
transform 1 0 8372 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1649977179
transform -1 0 16192 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1649977179
transform -1 0 15548 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1649977179
transform 1 0 10488 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1649977179
transform -1 0 15456 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1649977179
transform 1 0 22816 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1649977179
transform -1 0 25852 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1649977179
transform -1 0 28244 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1649977179
transform -1 0 28612 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1649977179
transform 1 0 24932 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1649977179
transform -1 0 27784 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1649977179
transform -1 0 31004 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1649977179
transform -1 0 30268 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1649977179
transform -1 0 20700 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1649977179
transform 1 0 22448 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1649977179
transform 1 0 15364 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1649977179
transform 1 0 20884 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1649977179
transform -1 0 31004 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1649977179
transform -1 0 30912 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1649977179
transform -1 0 28428 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1649977179
transform 1 0 24196 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1649977179
transform -1 0 23276 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1649977179
transform -1 0 23460 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1649977179
transform -1 0 11040 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1649977179
transform -1 0 12972 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1649977179
transform -1 0 14352 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1649977179
transform -1 0 13616 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1649977179
transform 1 0 14352 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1649977179
transform -1 0 18676 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1649977179
transform -1 0 19136 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1649977179
transform -1 0 18584 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1649977179
transform -1 0 17296 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1649977179
transform -1 0 10212 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1649977179
transform 1 0 8188 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22172 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 12236 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1649977179
transform 1 0 31188 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1649977179
transform 1 0 6716 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1649977179
transform 1 0 5520 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1649977179
transform -1 0 10856 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1649977179
transform 1 0 18124 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1649977179
transform 1 0 20516 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1649977179
transform 1 0 24656 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1649977179
transform 1 0 26036 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1649977179
transform 1 0 33580 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1649977179
transform 1 0 34960 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1649977179
transform -1 0 29072 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1649977179
transform 1 0 33948 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1649977179
transform 1 0 37536 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1649977179
transform 1 0 35052 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1649977179
transform 1 0 27968 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1649977179
transform -1 0 25668 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1649977179
transform -1 0 7176 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1649977179
transform 1 0 5428 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1649977179
transform 1 0 11224 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 19228 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 19872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 11040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1649977179
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input18 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1649977179
transform -1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform -1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1649977179
transform -1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1649977179
transform -1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform -1 0 9292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform -1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform -1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 15640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform -1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_43 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 45264 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_44
timestamp 1649977179
transform -1 0 55568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_45
timestamp 1649977179
transform -1 0 65136 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_46
timestamp 1649977179
transform -1 0 25392 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_47
timestamp 1649977179
transform -1 0 35328 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_48
timestamp 1649977179
transform -1 0 5520 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_49
timestamp 1649977179
transform -1 0 15456 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_50
timestamp 1649977179
transform 1 0 67896 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_51
timestamp 1649977179
transform 1 0 67436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_52
timestamp 1649977179
transform 1 0 66792 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_53
timestamp 1649977179
transform 1 0 67436 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_54
timestamp 1649977179
transform -1 0 58788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_55
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_56
timestamp 1649977179
transform -1 0 56488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_57
timestamp 1649977179
transform -1 0 57500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_58
timestamp 1649977179
transform -1 0 57132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_59
timestamp 1649977179
transform -1 0 59432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_60
timestamp 1649977179
transform -1 0 58144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_61
timestamp 1649977179
transform -1 0 58788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_62
timestamp 1649977179
transform -1 0 58788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_63
timestamp 1649977179
transform -1 0 59432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_64
timestamp 1649977179
transform -1 0 60720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_65
timestamp 1649977179
transform -1 0 58144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_66
timestamp 1649977179
transform -1 0 60076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_67
timestamp 1649977179
transform -1 0 57500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_68
timestamp 1649977179
transform -1 0 58144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_69
timestamp 1649977179
transform -1 0 59432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_70
timestamp 1649977179
transform -1 0 61364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_71
timestamp 1649977179
transform -1 0 58788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_72
timestamp 1649977179
transform -1 0 58788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_73
timestamp 1649977179
transform -1 0 60720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_74
timestamp 1649977179
transform -1 0 59432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_75
timestamp 1649977179
transform -1 0 60720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_76
timestamp 1649977179
transform -1 0 60076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_77
timestamp 1649977179
transform -1 0 62008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_78
timestamp 1649977179
transform -1 0 61364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_79
timestamp 1649977179
transform -1 0 59432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_80
timestamp 1649977179
transform -1 0 61364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_81
timestamp 1649977179
transform -1 0 62008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_82
timestamp 1649977179
transform -1 0 63296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_83
timestamp 1649977179
transform -1 0 60720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_84
timestamp 1649977179
transform -1 0 59064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_85
timestamp 1649977179
transform -1 0 59708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_86
timestamp 1649977179
transform -1 0 60720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_87
timestamp 1649977179
transform -1 0 62008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_88
timestamp 1649977179
transform -1 0 63940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_89
timestamp 1649977179
transform -1 0 61364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_90
timestamp 1649977179
transform -1 0 60352 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_91
timestamp 1649977179
transform -1 0 63296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_92
timestamp 1649977179
transform 1 0 67436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_93
timestamp 1649977179
transform 1 0 66792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_94
timestamp 1649977179
transform 1 0 67896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_95
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_96
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_97
timestamp 1649977179
transform 1 0 67896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_98
timestamp 1649977179
transform 1 0 67896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_99
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_100
timestamp 1649977179
transform 1 0 67436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_101
timestamp 1649977179
transform 1 0 67896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_102
timestamp 1649977179
transform 1 0 67896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103
timestamp 1649977179
transform 1 0 67436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform 1 0 67436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform 1 0 67896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform 1 0 67896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform 1 0 67896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform 1 0 67896 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform 1 0 67436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform 1 0 67436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform 1 0 67896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform 1 0 67896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform 1 0 67436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform 1 0 67436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform 1 0 67896 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform 1 0 67896 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform 1 0 67436 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform 1 0 67436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform 1 0 67896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform 1 0 67896 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform 1 0 67436 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform 1 0 67436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform 1 0 67896 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform 1 0 67896 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform 1 0 67436 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform 1 0 67436 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform 1 0 67896 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform -1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform -1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform -1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform -1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform -1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform -1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform -1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform 1 0 28796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform -1 0 30176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform -1 0 31004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform -1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform -1 0 32660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform -1 0 33488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform 1 0 33948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform -1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform 1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform -1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform -1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform -1 0 40756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform -1 0 41400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform -1 0 42044 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform -1 0 42872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 45356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform -1 0 46000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform -1 0 46644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform -1 0 47288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform -1 0 48116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform -1 0 49220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 50600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform -1 0 51244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform -1 0 51888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 53728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform 1 0 67436 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform 1 0 67896 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform -1 0 19228 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform -1 0 17296 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform -1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform -1 0 18952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_278
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_279
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_280
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_281
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_282
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 44914 59200 44970 60000 0 FreeSans 224 90 0 0 Sh
port 0 nsew signal tristate
flabel metal2 s 54850 59200 54906 60000 0 FreeSans 224 90 0 0 Sh_cmp
port 1 nsew signal tristate
flabel metal2 s 64786 59200 64842 60000 0 FreeSans 224 90 0 0 Sh_rst
port 2 nsew signal tristate
flabel metal2 s 25042 59200 25098 60000 0 FreeSans 224 90 0 0 Sw1
port 3 nsew signal tristate
flabel metal2 s 34978 59200 35034 60000 0 FreeSans 224 90 0 0 Sw2
port 4 nsew signal tristate
flabel metal2 s 5170 59200 5226 60000 0 FreeSans 224 90 0 0 Vd1
port 5 nsew signal tristate
flabel metal2 s 15106 59200 15162 60000 0 FreeSans 224 90 0 0 Vd2
port 6 nsew signal tristate
flabel metal3 s 69200 52368 70000 52488 0 FreeSans 480 0 0 0 clk_o
port 7 nsew signal tristate
flabel metal3 s 69200 59168 70000 59288 0 FreeSans 480 0 0 0 counter_rst
port 8 nsew signal tristate
flabel metal3 s 69200 57808 70000 57928 0 FreeSans 480 0 0 0 data_o
port 9 nsew signal tristate
flabel metal3 s 69200 55088 70000 55208 0 FreeSans 480 0 0 0 done_o
port 10 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 io_in[0]
port 11 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_in[10]
port 12 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[11]
port 13 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 io_in[12]
port 14 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 io_in[13]
port 15 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 io_in[14]
port 16 nsew signal input
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 io_in[15]
port 17 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_in[16]
port 18 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 io_in[17]
port 19 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 io_in[18]
port 20 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_in[19]
port 21 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_in[1]
port 22 nsew signal input
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 io_in[20]
port 23 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 io_in[21]
port 24 nsew signal input
flabel metal3 s 0 35096 800 35216 0 FreeSans 480 0 0 0 io_in[22]
port 25 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 io_in[23]
port 26 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_in[24]
port 27 nsew signal input
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 io_in[25]
port 28 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 io_in[26]
port 29 nsew signal input
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 io_in[27]
port 30 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 io_in[28]
port 31 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_in[29]
port 32 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_in[2]
port 33 nsew signal input
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 io_in[30]
port 34 nsew signal input
flabel metal3 s 0 48560 800 48680 0 FreeSans 480 0 0 0 io_in[31]
port 35 nsew signal input
flabel metal3 s 0 50056 800 50176 0 FreeSans 480 0 0 0 io_in[32]
port 36 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 io_in[33]
port 37 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 io_in[34]
port 38 nsew signal input
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 io_in[35]
port 39 nsew signal input
flabel metal3 s 0 56040 800 56160 0 FreeSans 480 0 0 0 io_in[36]
port 40 nsew signal input
flabel metal3 s 0 57536 800 57656 0 FreeSans 480 0 0 0 io_in[37]
port 41 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 io_in[3]
port 42 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_in[4]
port 43 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[5]
port 44 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_in[6]
port 45 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_in[7]
port 46 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_in[8]
port 47 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_in[9]
port 48 nsew signal input
flabel metal2 s 55954 0 56010 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 49 nsew signal tristate
flabel metal2 s 56874 0 56930 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 50 nsew signal tristate
flabel metal2 s 56966 0 57022 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 51 nsew signal tristate
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 52 nsew signal tristate
flabel metal2 s 57150 0 57206 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 53 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 54 nsew signal tristate
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 55 nsew signal tristate
flabel metal2 s 57426 0 57482 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 56 nsew signal tristate
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 57 nsew signal tristate
flabel metal2 s 57610 0 57666 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 58 nsew signal tristate
flabel metal2 s 57702 0 57758 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 59 nsew signal tristate
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 60 nsew signal tristate
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 61 nsew signal tristate
flabel metal2 s 57886 0 57942 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 62 nsew signal tristate
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 63 nsew signal tristate
flabel metal2 s 58070 0 58126 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 64 nsew signal tristate
flabel metal2 s 58162 0 58218 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 65 nsew signal tristate
flabel metal2 s 58254 0 58310 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 66 nsew signal tristate
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 67 nsew signal tristate
flabel metal2 s 58438 0 58494 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 68 nsew signal tristate
flabel metal2 s 58530 0 58586 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 69 nsew signal tristate
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 70 nsew signal tristate
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 71 nsew signal tristate
flabel metal2 s 58714 0 58770 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 72 nsew signal tristate
flabel metal2 s 58806 0 58862 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 73 nsew signal tristate
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 74 nsew signal tristate
flabel metal2 s 58990 0 59046 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 75 nsew signal tristate
flabel metal2 s 59082 0 59138 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 76 nsew signal tristate
flabel metal2 s 59174 0 59230 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 77 nsew signal tristate
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 78 nsew signal tristate
flabel metal2 s 59358 0 59414 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 79 nsew signal tristate
flabel metal2 s 56230 0 56286 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 80 nsew signal tristate
flabel metal2 s 56322 0 56378 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 81 nsew signal tristate
flabel metal2 s 56414 0 56470 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 82 nsew signal tristate
flabel metal2 s 56506 0 56562 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 83 nsew signal tristate
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 84 nsew signal tristate
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 85 nsew signal tristate
flabel metal2 s 56782 0 56838 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 86 nsew signal tristate
flabel metal3 s 69200 688 70000 808 0 FreeSans 480 0 0 0 io_out[0]
port 87 nsew signal tristate
flabel metal3 s 69200 14288 70000 14408 0 FreeSans 480 0 0 0 io_out[10]
port 88 nsew signal tristate
flabel metal3 s 69200 15648 70000 15768 0 FreeSans 480 0 0 0 io_out[11]
port 89 nsew signal tristate
flabel metal3 s 69200 17008 70000 17128 0 FreeSans 480 0 0 0 io_out[12]
port 90 nsew signal tristate
flabel metal3 s 69200 18368 70000 18488 0 FreeSans 480 0 0 0 io_out[13]
port 91 nsew signal tristate
flabel metal3 s 69200 19728 70000 19848 0 FreeSans 480 0 0 0 io_out[14]
port 92 nsew signal tristate
flabel metal3 s 69200 21088 70000 21208 0 FreeSans 480 0 0 0 io_out[15]
port 93 nsew signal tristate
flabel metal3 s 69200 22448 70000 22568 0 FreeSans 480 0 0 0 io_out[16]
port 94 nsew signal tristate
flabel metal3 s 69200 23808 70000 23928 0 FreeSans 480 0 0 0 io_out[17]
port 95 nsew signal tristate
flabel metal3 s 69200 25168 70000 25288 0 FreeSans 480 0 0 0 io_out[18]
port 96 nsew signal tristate
flabel metal3 s 69200 26528 70000 26648 0 FreeSans 480 0 0 0 io_out[19]
port 97 nsew signal tristate
flabel metal3 s 69200 2048 70000 2168 0 FreeSans 480 0 0 0 io_out[1]
port 98 nsew signal tristate
flabel metal3 s 69200 27888 70000 28008 0 FreeSans 480 0 0 0 io_out[20]
port 99 nsew signal tristate
flabel metal3 s 69200 29248 70000 29368 0 FreeSans 480 0 0 0 io_out[21]
port 100 nsew signal tristate
flabel metal3 s 69200 30608 70000 30728 0 FreeSans 480 0 0 0 io_out[22]
port 101 nsew signal tristate
flabel metal3 s 69200 31968 70000 32088 0 FreeSans 480 0 0 0 io_out[23]
port 102 nsew signal tristate
flabel metal3 s 69200 33328 70000 33448 0 FreeSans 480 0 0 0 io_out[24]
port 103 nsew signal tristate
flabel metal3 s 69200 34688 70000 34808 0 FreeSans 480 0 0 0 io_out[25]
port 104 nsew signal tristate
flabel metal3 s 69200 36048 70000 36168 0 FreeSans 480 0 0 0 io_out[26]
port 105 nsew signal tristate
flabel metal3 s 69200 37408 70000 37528 0 FreeSans 480 0 0 0 io_out[27]
port 106 nsew signal tristate
flabel metal3 s 69200 38768 70000 38888 0 FreeSans 480 0 0 0 io_out[28]
port 107 nsew signal tristate
flabel metal3 s 69200 40128 70000 40248 0 FreeSans 480 0 0 0 io_out[29]
port 108 nsew signal tristate
flabel metal3 s 69200 3408 70000 3528 0 FreeSans 480 0 0 0 io_out[2]
port 109 nsew signal tristate
flabel metal3 s 69200 41488 70000 41608 0 FreeSans 480 0 0 0 io_out[30]
port 110 nsew signal tristate
flabel metal3 s 69200 42848 70000 42968 0 FreeSans 480 0 0 0 io_out[31]
port 111 nsew signal tristate
flabel metal3 s 69200 44208 70000 44328 0 FreeSans 480 0 0 0 io_out[32]
port 112 nsew signal tristate
flabel metal3 s 69200 45568 70000 45688 0 FreeSans 480 0 0 0 io_out[33]
port 113 nsew signal tristate
flabel metal3 s 69200 46928 70000 47048 0 FreeSans 480 0 0 0 io_out[34]
port 114 nsew signal tristate
flabel metal3 s 69200 48288 70000 48408 0 FreeSans 480 0 0 0 io_out[35]
port 115 nsew signal tristate
flabel metal3 s 69200 49648 70000 49768 0 FreeSans 480 0 0 0 io_out[36]
port 116 nsew signal tristate
flabel metal3 s 69200 51008 70000 51128 0 FreeSans 480 0 0 0 io_out[37]
port 117 nsew signal tristate
flabel metal3 s 69200 4768 70000 4888 0 FreeSans 480 0 0 0 io_out[3]
port 118 nsew signal tristate
flabel metal3 s 69200 6128 70000 6248 0 FreeSans 480 0 0 0 io_out[4]
port 119 nsew signal tristate
flabel metal3 s 69200 7488 70000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 120 nsew signal tristate
flabel metal3 s 69200 8848 70000 8968 0 FreeSans 480 0 0 0 io_out[6]
port 121 nsew signal tristate
flabel metal3 s 69200 10208 70000 10328 0 FreeSans 480 0 0 0 io_out[7]
port 122 nsew signal tristate
flabel metal3 s 69200 11568 70000 11688 0 FreeSans 480 0 0 0 io_out[8]
port 123 nsew signal tristate
flabel metal3 s 69200 12928 70000 13048 0 FreeSans 480 0 0 0 io_out[9]
port 124 nsew signal tristate
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 irq[0]
port 125 nsew signal tristate
flabel metal2 s 55770 0 55826 800 0 FreeSans 224 90 0 0 irq[1]
port 126 nsew signal tristate
flabel metal2 s 55862 0 55918 800 0 FreeSans 224 90 0 0 irq[2]
port 127 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 128 nsew signal input
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 129 nsew signal input
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 130 nsew signal input
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 131 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 132 nsew signal input
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 133 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 134 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 135 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 136 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 137 nsew signal input
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 138 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 139 nsew signal input
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 140 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 141 nsew signal input
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 142 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 143 nsew signal input
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 144 nsew signal input
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 145 nsew signal input
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 146 nsew signal input
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 147 nsew signal input
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 148 nsew signal input
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 149 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 150 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 151 nsew signal input
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 152 nsew signal input
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 153 nsew signal input
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 154 nsew signal input
flabel metal2 s 54574 0 54630 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 155 nsew signal input
flabel metal2 s 54850 0 54906 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 156 nsew signal input
flabel metal2 s 55126 0 55182 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 157 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 158 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 159 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 160 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 161 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 162 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 163 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 164 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 165 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 166 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 167 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 168 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 169 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 170 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 171 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 172 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 173 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 174 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 175 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 176 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 177 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 178 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 179 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 180 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 181 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 182 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 183 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 184 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 185 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 186 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 187 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 188 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 189 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 190 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 191 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 192 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 193 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 194 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 195 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 196 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 197 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 198 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 199 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 200 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 201 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 202 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 203 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 204 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 205 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 206 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 207 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 208 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 209 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 210 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 211 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 212 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 213 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 214 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 215 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 216 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 217 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 218 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 219 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 220 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 221 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 222 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 223 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 224 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 225 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 226 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 227 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 228 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 229 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 230 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 231 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 232 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 233 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 234 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 235 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 236 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 237 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 238 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 239 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 240 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 241 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 242 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 243 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 244 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 245 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 246 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 247 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 248 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 249 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 250 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 251 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 252 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 253 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 254 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 255 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 256 nsew signal tristate
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 257 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 258 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 259 nsew signal tristate
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 260 nsew signal tristate
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 261 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 262 nsew signal tristate
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 263 nsew signal tristate
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 264 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 265 nsew signal tristate
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 266 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 267 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 268 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 269 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 270 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 271 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 272 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 273 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 274 nsew signal tristate
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 275 nsew signal tristate
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 276 nsew signal tristate
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 277 nsew signal tristate
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 278 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 279 nsew signal tristate
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 280 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 281 nsew signal tristate
flabel metal2 s 54390 0 54446 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 282 nsew signal tristate
flabel metal2 s 54666 0 54722 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 283 nsew signal tristate
flabel metal2 s 54942 0 54998 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 284 nsew signal tristate
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 285 nsew signal tristate
flabel metal2 s 55494 0 55550 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 286 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 287 nsew signal tristate
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 288 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 289 nsew signal tristate
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 290 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 291 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 292 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 293 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 294 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 295 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 296 nsew signal tristate
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 297 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 298 nsew signal tristate
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 299 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 300 nsew signal tristate
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 301 nsew signal tristate
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 302 nsew signal tristate
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 303 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 304 nsew signal tristate
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 305 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 306 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 307 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 308 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 309 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 310 nsew signal tristate
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 311 nsew signal tristate
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 312 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 313 nsew signal tristate
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 314 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 315 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 316 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 317 nsew signal tristate
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 318 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 319 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 320 nsew signal tristate
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 321 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 322 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 323 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 324 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 325 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 326 nsew signal tristate
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 327 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 328 nsew signal tristate
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 329 nsew signal tristate
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 330 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 331 nsew signal tristate
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 332 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 333 nsew signal tristate
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 334 nsew signal tristate
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 335 nsew signal tristate
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 336 nsew signal tristate
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 337 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 338 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 339 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 340 nsew signal tristate
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 341 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 342 nsew signal tristate
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 343 nsew signal tristate
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 344 nsew signal tristate
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 345 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 346 nsew signal tristate
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 347 nsew signal tristate
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 348 nsew signal tristate
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 349 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 350 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 351 nsew signal tristate
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 352 nsew signal tristate
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 353 nsew signal tristate
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 354 nsew signal tristate
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 355 nsew signal tristate
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 356 nsew signal tristate
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 357 nsew signal tristate
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 358 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 359 nsew signal tristate
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 360 nsew signal tristate
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 361 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 362 nsew signal tristate
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 363 nsew signal tristate
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 364 nsew signal tristate
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 365 nsew signal tristate
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 366 nsew signal tristate
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 367 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 368 nsew signal tristate
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 369 nsew signal tristate
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 370 nsew signal tristate
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 371 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 372 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 373 nsew signal tristate
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 374 nsew signal tristate
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 375 nsew signal tristate
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 376 nsew signal tristate
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 377 nsew signal tristate
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 378 nsew signal tristate
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 379 nsew signal tristate
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 380 nsew signal tristate
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 381 nsew signal tristate
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 382 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 383 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 384 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 385 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 386 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 387 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 388 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 389 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 390 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 391 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 392 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 393 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 394 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 395 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 396 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 397 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 398 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 399 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 400 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 401 nsew signal input
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 402 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 403 nsew signal input
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 404 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 405 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 406 nsew signal input
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 407 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 408 nsew signal input
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 409 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 410 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 411 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 412 nsew signal input
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 413 nsew signal input
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 414 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 415 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 416 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 417 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 418 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 419 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 420 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 421 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 422 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 423 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 424 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 425 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 426 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 427 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 428 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 429 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 430 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 431 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 432 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 433 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 434 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 435 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 436 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 437 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 438 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 439 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 440 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 441 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 442 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 443 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 444 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 445 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 446 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 447 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 448 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 449 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 450 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 451 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 452 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 453 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 454 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 455 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 456 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 457 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 458 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 459 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 460 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 461 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 462 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 463 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 464 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 465 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 466 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 467 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 468 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 469 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 470 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 471 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 472 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 473 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 474 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 475 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 476 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 477 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 478 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 479 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 480 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 481 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 482 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 483 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 484 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 485 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 486 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 487 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 488 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 489 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 490 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 491 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 492 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 493 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 494 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 495 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 496 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 497 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 498 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 499 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 500 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 501 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 502 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 503 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 504 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 505 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 506 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 507 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 508 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 509 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 510 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 511 nsew signal input
flabel metal3 s 69200 53728 70000 53848 0 FreeSans 480 0 0 0 rst_o
port 512 nsew signal tristate
flabel metal3 s 69200 56448 70000 56568 0 FreeSans 480 0 0 0 start_o
port 513 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 514 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 514 nsew power bidirectional
flabel metal4 s 65648 2128 65968 57712 0 FreeSans 1920 90 0 0 vccd1
port 514 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 515 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 515 nsew ground bidirectional
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wb_clk_i
port 516 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wb_rst_i
port 517 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 518 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 519 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 520 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 521 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 522 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 523 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 524 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 525 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 526 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 527 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 528 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 529 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 530 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 531 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 532 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 533 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 534 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 535 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 536 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 537 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 538 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 539 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 540 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 541 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 542 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 543 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 544 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 545 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 546 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 547 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 548 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 549 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 550 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 551 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 552 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 553 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 554 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 555 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 556 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 557 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 558 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 559 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 560 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 561 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 562 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 563 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 564 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 565 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 566 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 567 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 568 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 569 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 570 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 571 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 572 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 573 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 574 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 575 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 576 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 577 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 578 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 579 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 580 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 581 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 582 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 583 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 584 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 585 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 586 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 587 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 588 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 589 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 590 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 591 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 592 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 593 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 594 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 595 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 596 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 597 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 598 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 599 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 600 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 601 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 602 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 603 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 604 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 605 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 606 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 607 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 608 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 609 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 610 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 611 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 612 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 613 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 614 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 615 nsew signal tristate
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 616 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 617 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 618 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 619 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 620 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_we_i
port 621 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 60000
<< end >>
