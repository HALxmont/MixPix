magic
tech sky130A
magscale 1 2
timestamp 1668297577
<< dnwell >>
rect 30500 5100 49800 6500
rect 30500 1900 37500 5100
rect 42700 1900 49800 5100
rect 30500 500 49800 1900
<< photodiode >>
rect 39700 3300 40300 3900
<< nwell >>
rect 30300 6100 50000 6700
rect 30300 900 30900 6100
rect 37100 5000 43100 5500
rect 37100 2000 37600 5000
rect 39860 3460 40140 3740
rect 42600 2000 43100 5000
rect 37100 1500 43100 2000
rect 49400 900 50000 6100
rect 30300 300 50000 900
<< pwell >>
rect 30000 6700 50300 7000
rect 30000 300 30300 6700
rect 50000 300 50300 6700
rect 30000 0 50300 300
rect 44600 -520 44660 -440
rect 45120 -520 45180 -440
rect 45620 -520 45680 -440
rect 46140 -520 46200 -440
rect 43780 -580 46960 -520
<< psubdiff >>
rect 30100 6800 30300 6900
rect 50000 6800 50200 6900
rect 30100 6700 30200 6800
rect 50100 6700 50200 6800
rect 30100 200 30200 300
rect 50100 200 50200 300
rect 30100 100 30300 200
rect 50000 100 50200 200
<< nsubdiff >>
rect 30500 6300 30700 6500
rect 39300 6300 39500 6500
rect 40500 6300 40700 6500
rect 49600 6300 49800 6500
rect 37300 3900 37500 4300
rect 42700 3900 42900 4300
rect 39920 3640 40080 3680
rect 39920 3560 39960 3640
rect 40040 3560 40080 3640
rect 39920 3520 40080 3560
rect 37300 2900 37500 3300
rect 42700 2900 42900 3300
rect 30500 500 30700 700
rect 39300 500 39500 700
rect 40500 500 40700 700
rect 49600 500 49800 700
<< psubdiffcont >>
rect 30300 6800 50000 6900
rect 30100 300 30200 6700
rect 50100 300 50200 6700
rect 30300 100 50000 200
<< nsubdiffcont >>
rect 39500 6300 40500 6500
rect 30500 700 30700 6300
rect 37300 3300 37500 3900
rect 39960 3560 40040 3640
rect 42700 3300 42900 3900
rect 49600 700 49800 6300
rect 39500 500 40500 700
<< locali >>
rect 51700 7600 52500 8700
rect 30100 6900 53200 7600
rect 30100 6800 30300 6900
rect 50000 6800 53200 6900
rect 30100 6700 30200 6800
rect 50100 6700 50200 6800
rect 30500 6300 30700 6500
rect 39300 6300 39500 6500
rect 40500 6300 40700 6500
rect 49600 6300 49800 6500
rect 37300 3900 37500 4300
rect 42700 3900 42900 4300
rect 39900 3640 40100 3700
rect 39900 3560 39960 3640
rect 40040 3560 40100 3640
rect 39900 3500 40100 3560
rect 37300 2900 37500 3300
rect 39950 1230 40050 3500
rect 42700 2900 42900 3300
rect 39950 1130 41080 1230
rect 30500 500 30700 700
rect 39300 500 39500 700
rect 40500 500 40700 700
rect 40980 400 41080 1130
rect 49600 500 49800 700
rect 30100 200 30200 300
rect 50100 200 50200 300
rect 30100 100 30300 200
rect 50000 100 50200 200
rect 42500 0 47100 100
rect 44020 -460 44140 0
rect 44340 -180 44400 0
rect 44860 -180 44920 0
rect 45360 -180 45420 0
rect 45880 -180 45940 0
rect 46400 -180 46460 0
rect 46920 -180 46980 0
<< viali >>
rect 51700 8700 52500 9500
rect 40980 300 41080 400
<< metal1 >>
rect 51694 9506 52506 9512
rect 51688 8706 51694 9506
rect 52506 8706 52512 9506
rect 51688 8700 51700 8706
rect 52500 8700 52512 8706
rect 51688 8694 52512 8700
rect 50050 8600 50150 8606
rect 40968 400 41092 406
rect 40968 300 40980 400
rect 41080 300 41092 400
rect 40968 294 41092 300
rect 40980 -150 41080 294
rect 50050 150 50150 8500
rect 42800 50 50150 150
rect 40980 -250 42600 -150
rect 42100 -450 42200 -250
rect 42800 -350 42900 50
rect 43100 -450 43200 50
rect 43400 -400 43750 -200
rect 42100 -556 42200 -550
rect 42650 -800 42750 -500
rect 41000 -900 42750 -800
rect 43050 -800 43150 -794
rect 43250 -800 43350 -500
rect 43150 -900 43350 -800
rect 41000 -1040 41100 -900
rect 43050 -906 43150 -900
rect 43540 -960 43660 -400
rect 44600 -520 44660 -440
rect 45120 -520 45180 -440
rect 45620 -520 45680 -440
rect 46140 -520 46200 -440
rect 46660 -520 46720 -440
rect 43780 -580 46960 -520
rect 40990 -1050 41110 -1040
rect 40990 -1150 41000 -1050
rect 41100 -1150 41110 -1050
rect 43540 -1086 43660 -1080
rect 45440 -980 45560 -580
rect 45440 -1106 45560 -1100
rect 40990 -1160 41110 -1150
<< via1 >>
rect 51694 9500 52506 9506
rect 51694 8706 51700 9500
rect 51700 8706 52500 9500
rect 52500 8706 52506 9500
rect 50050 8500 50150 8600
rect 42100 -550 42200 -450
rect 43050 -900 43150 -800
rect 41000 -1150 41100 -1050
rect 43540 -1080 43660 -960
rect 45440 -1100 45560 -980
<< obsm1 >>
rect 30900 900 49400 6100
<< metal2 >>
rect 51600 9506 52600 9600
rect 51600 8706 51694 9506
rect 52506 8706 52600 9506
rect 50050 8600 50150 8609
rect 51600 8600 52600 8706
rect 50044 8500 50050 8600
rect 50150 8500 50156 8600
rect 50050 8491 50150 8500
rect 42094 -550 42100 -450
rect 42200 -550 42206 -450
rect 42100 -800 42200 -550
rect 42100 -900 43050 -800
rect 43150 -900 43156 -800
rect 40960 -1050 41160 -1030
rect 40960 -1150 41000 -1050
rect 41100 -1150 41160 -1050
rect 43534 -1080 43540 -960
rect 43660 -1080 43666 -960
rect 40960 -1200 41160 -1150
rect 43540 -1200 43660 -1080
rect 45434 -1100 45440 -980
rect 45560 -1100 45566 -980
rect 45440 -1200 45560 -1100
rect 40600 -2600 41500 -1200
rect 43200 -2600 44100 -1200
rect 45200 -2600 46100 -1200
<< via2 >>
rect 51694 8706 52506 9506
rect 50050 8500 50150 8600
<< obsm2 >>
rect 30100 100 50100 6900
<< metal3 >>
rect 51600 9511 52600 9600
rect 51600 8701 51689 9511
rect 52511 8701 52600 9511
rect 50045 8605 50155 8611
rect 51600 8600 52600 8701
rect 50045 8500 50050 8505
rect 50150 8500 50155 8505
rect 50045 8495 50155 8500
<< via3 >>
rect 51689 9506 52511 9511
rect 51689 8706 51694 9506
rect 51694 8706 52506 9506
rect 52506 8706 52511 9506
rect 51689 8701 52511 8706
rect 50045 8600 50155 8605
rect 50045 8505 50050 8600
rect 50050 8505 50150 8600
rect 50150 8505 50155 8600
<< metal4 >>
rect 49300 13400 54100 14200
rect 49300 12600 54094 13400
rect 51688 9511 52512 9512
rect 51688 9500 51689 9511
rect 49300 8701 51689 9500
rect 52511 9506 52512 9511
rect 52511 9500 55100 9506
rect 52511 8701 55300 9500
rect 49300 8700 55300 8701
rect 50050 8606 50150 8700
rect 50044 8605 50156 8606
rect 50044 8505 50045 8605
rect 50155 8505 50156 8605
rect 50044 8504 50156 8505
<< fillblock >>
rect 30200 200 50000 6800
use sky130_fd_pr__nfet_01v8_lvt_M9TU6H  sky130_fd_pr__nfet_01v8_lvt_M9TU6H_0
timestamp 1668272048
transform -1 0 42696 0 -1 -321
box -296 -379 296 379
use sky130_fd_pr__nfet_01v8_lvt_M9TU6H  sky130_fd_pr__nfet_01v8_lvt_M9TU6H_1
timestamp 1668272048
transform -1 0 43296 0 -1 -321
box -296 -379 296 379
use sky130_fd_pr__nfet_01v8_lvt_M9TU6H  sky130_fd_pr__nfet_01v8_lvt_M9TU6H_2
timestamp 1668272048
transform -1 0 43896 0 -1 -321
box -296 -379 296 379
use sky130_fd_pr__nfet_01v8_lvt_X3BG59  sky130_fd_pr__nfet_01v8_lvt_X3BG59_0
timestamp 1668272609
transform -1 0 45657 0 -1 -321
box -1457 -379 1457 379
<< labels >>
flabel metal4 54000 13400 54000 13400 0 FreeSans 1600 0 0 0 VDD
port 0 nsew power input
flabel metal4 55000 9100 55000 9100 0 FreeSans 1600 0 0 0 VSS
port 1 nsew ground input
flabel metal2 41000 -2500 41000 -2500 0 FreeSans 1600 0 0 0 RST
port 2 nsew signal input
flabel metal2 43600 -2500 43600 -2500 0 FreeSans 1600 0 0 0 OUT
port 3 nsew signal output
flabel metal2 45600 -2500 45600 -2500 0 FreeSans 1600 0 0 0 IP
port 4 nsew signal input
<< end >>
