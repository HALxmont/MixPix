magic
tech sky130B
magscale 1 2
timestamp 1667829310
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 137830 700816 137836 700868
rect 137888 700856 137894 700868
rect 157334 700856 157340 700868
rect 137888 700828 157340 700856
rect 137888 700816 137894 700828
rect 157334 700816 157340 700828
rect 157392 700816 157398 700868
rect 155954 700748 155960 700800
rect 156012 700788 156018 700800
rect 202782 700788 202788 700800
rect 156012 700760 202788 700788
rect 156012 700748 156018 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 160738 700720 160744 700732
rect 89220 700692 160744 700720
rect 89220 700680 89226 700692
rect 160738 700680 160744 700692
rect 160796 700680 160802 700732
rect 154574 700612 154580 700664
rect 154632 700652 154638 700664
rect 267642 700652 267648 700664
rect 154632 700624 267648 700652
rect 154632 700612 154638 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 24302 700544 24308 700596
rect 24360 700584 24366 700596
rect 162210 700584 162216 700596
rect 24360 700556 162216 700584
rect 24360 700544 24366 700556
rect 162210 700544 162216 700556
rect 162268 700544 162274 700596
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 162118 700516 162124 700528
rect 8168 700488 162124 700516
rect 8168 700476 8174 700488
rect 162118 700476 162124 700488
rect 162176 700476 162182 700528
rect 153286 700408 153292 700460
rect 153344 700448 153350 700460
rect 332502 700448 332508 700460
rect 153344 700420 332508 700448
rect 153344 700408 153350 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 152458 700340 152464 700392
rect 152516 700380 152522 700392
rect 413646 700380 413652 700392
rect 152516 700352 413652 700380
rect 152516 700340 152522 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 489178 700340 489184 700392
rect 489236 700380 489242 700392
rect 527174 700380 527180 700392
rect 489236 700352 527180 700380
rect 489236 700340 489242 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 527818 700340 527824 700392
rect 527876 700380 527882 700392
rect 559650 700380 559656 700392
rect 527876 700352 559656 700380
rect 527876 700340 527882 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 148318 700272 148324 700324
rect 148376 700312 148382 700324
rect 543458 700312 543464 700324
rect 148376 700284 543464 700312
rect 148376 700272 148382 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 146294 696940 146300 696992
rect 146352 696980 146358 696992
rect 580166 696980 580172 696992
rect 146352 696952 580172 696980
rect 146352 696940 146358 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 161474 683244 161480 683256
rect 3476 683216 161480 683244
rect 3476 683204 3482 683216
rect 161474 683204 161480 683216
rect 161532 683204 161538 683256
rect 146938 683136 146944 683188
rect 146996 683176 147002 683188
rect 580166 683176 580172 683188
rect 146996 683148 580172 683176
rect 146996 683136 147002 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 163498 670732 163504 670744
rect 3568 670704 163504 670732
rect 3568 670692 3574 670704
rect 163498 670692 163504 670704
rect 163556 670692 163562 670744
rect 498838 670692 498844 670744
rect 498896 670732 498902 670744
rect 580166 670732 580172 670744
rect 498896 670704 580172 670732
rect 498896 670692 498902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 163590 656928 163596 656940
rect 3476 656900 163596 656928
rect 3476 656888 3482 656900
rect 163590 656888 163596 656900
rect 163648 656888 163654 656940
rect 182818 643084 182824 643136
rect 182876 643124 182882 643136
rect 580166 643124 580172 643136
rect 182876 643096 580172 643124
rect 182876 643084 182882 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 164234 632108 164240 632120
rect 3476 632080 164240 632108
rect 3476 632068 3482 632080
rect 164234 632068 164240 632080
rect 164292 632068 164298 632120
rect 188338 630640 188344 630692
rect 188396 630680 188402 630692
rect 580166 630680 580172 630692
rect 188396 630652 580172 630680
rect 188396 630640 188402 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 164878 618304 164884 618316
rect 3200 618276 164884 618304
rect 3200 618264 3206 618276
rect 164878 618264 164884 618276
rect 164936 618264 164942 618316
rect 143626 616836 143632 616888
rect 143684 616876 143690 616888
rect 580166 616876 580172 616888
rect 143684 616848 580172 616876
rect 143684 616836 143690 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 164970 605860 164976 605872
rect 3292 605832 164976 605860
rect 3292 605820 3298 605832
rect 164970 605820 164976 605832
rect 165028 605820 165034 605872
rect 142338 590656 142344 590708
rect 142396 590696 142402 590708
rect 579798 590696 579804 590708
rect 142396 590668 579804 590696
rect 142396 590656 142402 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 165614 579680 165620 579692
rect 3384 579652 165620 579680
rect 3384 579640 3390 579652
rect 165614 579640 165620 579652
rect 165672 579640 165678 579692
rect 144178 576852 144184 576904
rect 144236 576892 144242 576904
rect 580166 576892 580172 576904
rect 144236 576864 580172 576892
rect 144236 576852 144242 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 167638 565876 167644 565888
rect 3476 565848 167644 565876
rect 3476 565836 3482 565848
rect 167638 565836 167644 565848
rect 167696 565836 167702 565888
rect 142798 563048 142804 563100
rect 142856 563088 142862 563100
rect 579798 563088 579804 563100
rect 142856 563060 579804 563088
rect 142856 563048 142862 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 166258 553432 166264 553444
rect 3476 553404 166264 553432
rect 3476 553392 3482 553404
rect 166258 553392 166264 553404
rect 166316 553392 166322 553444
rect 181438 536800 181444 536852
rect 181496 536840 181502 536852
rect 580166 536840 580172 536852
rect 181496 536812 580172 536840
rect 181496 536800 181502 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 166994 527184 167000 527196
rect 3476 527156 167000 527184
rect 3476 527144 3482 527156
rect 166994 527144 167000 527156
rect 167052 527144 167058 527196
rect 142890 524424 142896 524476
rect 142948 524464 142954 524476
rect 580166 524464 580172 524476
rect 142948 524436 580172 524464
rect 142948 524424 142954 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 7558 514808 7564 514820
rect 3476 514780 7564 514808
rect 3476 514768 3482 514780
rect 7558 514768 7564 514780
rect 7616 514768 7622 514820
rect 180058 510620 180064 510672
rect 180116 510660 180122 510672
rect 580166 510660 580172 510672
rect 180116 510632 580172 510660
rect 180116 510620 180122 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 167730 501004 167736 501016
rect 3108 500976 167736 501004
rect 3108 500964 3114 500976
rect 167730 500964 167736 500976
rect 167788 500964 167794 501016
rect 139394 484372 139400 484424
rect 139452 484412 139458 484424
rect 580166 484412 580172 484424
rect 139452 484384 580172 484412
rect 139452 484372 139458 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 140038 470568 140044 470620
rect 140096 470608 140102 470620
rect 579982 470608 579988 470620
rect 140096 470580 579988 470608
rect 140096 470568 140102 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 170398 462380 170404 462392
rect 3568 462352 170404 462380
rect 3568 462340 3574 462352
rect 170398 462340 170404 462352
rect 170456 462340 170462 462392
rect 178678 456764 178684 456816
rect 178736 456804 178742 456816
rect 580166 456804 580172 456816
rect 178736 456776 580172 456804
rect 178736 456764 178742 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 157426 450508 157432 450560
rect 157484 450548 157490 450560
rect 169754 450548 169760 450560
rect 157484 450520 169760 450548
rect 157484 450508 157490 450520
rect 169754 450508 169760 450520
rect 169812 450508 169818 450560
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 170490 448576 170496 448588
rect 3200 448548 170496 448576
rect 3200 448536 3206 448548
rect 170490 448536 170496 448548
rect 170548 448536 170554 448588
rect 138658 430584 138664 430636
rect 138716 430624 138722 430636
rect 580166 430624 580172 430636
rect 138716 430596 580172 430624
rect 138716 430584 138722 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 169754 422328 169760 422340
rect 3568 422300 169760 422328
rect 3568 422288 3574 422300
rect 169754 422288 169760 422300
rect 169812 422288 169818 422340
rect 138750 418140 138756 418192
rect 138808 418180 138814 418192
rect 580166 418180 580172 418192
rect 138808 418152 580172 418180
rect 138808 418140 138814 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 171778 409884 171784 409896
rect 2924 409856 171784 409884
rect 2924 409844 2930 409856
rect 171778 409844 171784 409856
rect 171836 409844 171842 409896
rect 185578 404336 185584 404388
rect 185636 404376 185642 404388
rect 580166 404376 580172 404388
rect 185636 404348 580172 404376
rect 185636 404336 185642 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 171870 397508 171876 397520
rect 3568 397480 171876 397508
rect 3568 397468 3574 397480
rect 171870 397468 171876 397480
rect 171928 397468 171934 397520
rect 196618 378156 196624 378208
rect 196676 378196 196682 378208
rect 580166 378196 580172 378208
rect 196676 378168 580172 378196
rect 196676 378156 196682 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 2774 371288 2780 371340
rect 2832 371328 2838 371340
rect 4798 371328 4804 371340
rect 2832 371300 4804 371328
rect 2832 371288 2838 371300
rect 4798 371288 4804 371300
rect 4856 371288 4862 371340
rect 3510 358368 3516 358420
rect 3568 358408 3574 358420
rect 8938 358408 8944 358420
rect 3568 358380 8944 358408
rect 3568 358368 3574 358380
rect 8938 358368 8944 358380
rect 8996 358368 9002 358420
rect 135254 351908 135260 351960
rect 135312 351948 135318 351960
rect 580166 351948 580172 351960
rect 135312 351920 580172 351948
rect 135312 351908 135318 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 149698 345080 149704 345092
rect 3384 345052 149704 345080
rect 3384 345040 3390 345052
rect 149698 345040 149704 345052
rect 149756 345040 149762 345092
rect 134518 324300 134524 324352
rect 134576 324340 134582 324352
rect 580166 324340 580172 324352
rect 134576 324312 580172 324340
rect 134576 324300 134582 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 173894 318832 173900 318844
rect 3384 318804 173900 318832
rect 3384 318792 3390 318804
rect 173894 318792 173900 318804
rect 173952 318792 173958 318844
rect 135898 311856 135904 311908
rect 135956 311896 135962 311908
rect 579982 311896 579988 311908
rect 135956 311868 579988 311896
rect 135956 311856 135962 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 175918 305028 175924 305040
rect 3568 305000 175924 305028
rect 3568 304988 3574 305000
rect 175918 304988 175924 305000
rect 175976 304988 175982 305040
rect 134610 298120 134616 298172
rect 134668 298160 134674 298172
rect 580166 298160 580172 298172
rect 134668 298132 580172 298160
rect 134668 298120 134674 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 174538 292584 174544 292596
rect 3568 292556 174544 292584
rect 3568 292544 3574 292556
rect 174538 292544 174544 292556
rect 174596 292544 174602 292596
rect 145558 289076 145564 289128
rect 145616 289116 145622 289128
rect 188338 289116 188344 289128
rect 145616 289088 188344 289116
rect 145616 289076 145622 289088
rect 188338 289076 188344 289088
rect 188396 289076 188402 289128
rect 149054 287648 149060 287700
rect 149112 287688 149118 287700
rect 462314 287688 462320 287700
rect 149112 287660 462320 287688
rect 149112 287648 149118 287660
rect 462314 287648 462320 287660
rect 462372 287648 462378 287700
rect 137278 286288 137284 286340
rect 137336 286328 137342 286340
rect 196618 286328 196624 286340
rect 137336 286300 196624 286328
rect 137336 286288 137342 286300
rect 196618 286288 196624 286300
rect 196676 286288 196682 286340
rect 147674 283568 147680 283620
rect 147732 283608 147738 283620
rect 489178 283608 489184 283620
rect 147732 283580 489184 283608
rect 147732 283568 147738 283580
rect 489178 283568 489184 283580
rect 489236 283568 489242 283620
rect 144914 282140 144920 282192
rect 144972 282180 144978 282192
rect 182818 282180 182824 282192
rect 144972 282152 182824 282180
rect 144972 282140 144978 282152
rect 182818 282140 182824 282152
rect 182876 282140 182882 282192
rect 140774 280780 140780 280832
rect 140832 280820 140838 280832
rect 181438 280820 181444 280832
rect 140832 280792 181444 280820
rect 140832 280780 140838 280792
rect 181438 280780 181444 280792
rect 181496 280780 181502 280832
rect 40034 279420 40040 279472
rect 40092 279460 40098 279472
rect 160094 279460 160100 279472
rect 40092 279432 160100 279460
rect 40092 279420 40098 279432
rect 160094 279420 160100 279432
rect 160152 279420 160158 279472
rect 151078 275272 151084 275324
rect 151136 275312 151142 275324
rect 428458 275312 428464 275324
rect 151136 275284 428464 275312
rect 151136 275272 151142 275284
rect 428458 275272 428464 275284
rect 428516 275272 428522 275324
rect 8938 273912 8944 273964
rect 8996 273952 9002 273964
rect 173158 273952 173164 273964
rect 8996 273924 173164 273952
rect 8996 273912 9002 273924
rect 173158 273912 173164 273924
rect 173216 273912 173222 273964
rect 186682 273912 186688 273964
rect 186740 273952 186746 273964
rect 364334 273952 364340 273964
rect 186740 273924 364340 273952
rect 186740 273912 186746 273924
rect 364334 273912 364340 273924
rect 364392 273912 364398 273964
rect 151906 273232 151912 273284
rect 151964 273272 151970 273284
rect 186682 273272 186688 273284
rect 151964 273244 186688 273272
rect 151964 273232 151970 273244
rect 186682 273232 186688 273244
rect 186740 273272 186746 273284
rect 187142 273272 187148 273284
rect 186740 273244 187148 273272
rect 186740 273232 186746 273244
rect 187142 273232 187148 273244
rect 187200 273232 187206 273284
rect 133138 271872 133144 271924
rect 133196 271912 133202 271924
rect 580166 271912 580172 271924
rect 133196 271884 580172 271912
rect 133196 271872 133202 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 7558 271192 7564 271244
rect 7616 271232 7622 271244
rect 169018 271232 169024 271244
rect 7616 271204 169024 271232
rect 7616 271192 7622 271204
rect 169018 271192 169024 271204
rect 169076 271192 169082 271244
rect 149146 271124 149152 271176
rect 149204 271164 149210 271176
rect 494054 271164 494060 271176
rect 149204 271136 494060 271164
rect 149204 271124 149210 271136
rect 494054 271124 494060 271136
rect 494112 271124 494118 271176
rect 71774 269764 71780 269816
rect 71832 269804 71838 269816
rect 119982 269804 119988 269816
rect 71832 269776 119988 269804
rect 71832 269764 71838 269776
rect 119982 269764 119988 269776
rect 120040 269764 120046 269816
rect 147766 269764 147772 269816
rect 147824 269804 147830 269816
rect 527818 269804 527824 269816
rect 147824 269776 527824 269804
rect 147824 269764 147830 269776
rect 527818 269764 527824 269776
rect 527876 269764 527882 269816
rect 119982 269084 119988 269136
rect 120040 269124 120046 269136
rect 158714 269124 158720 269136
rect 120040 269096 158720 269124
rect 120040 269084 120046 269096
rect 158714 269084 158720 269096
rect 158772 269084 158778 269136
rect 4798 268404 4804 268456
rect 4856 268444 4862 268456
rect 172698 268444 172704 268456
rect 4856 268416 172704 268444
rect 4856 268404 4862 268416
rect 172698 268404 172704 268416
rect 172756 268404 172762 268456
rect 146202 268336 146208 268388
rect 146260 268376 146266 268388
rect 498838 268376 498844 268388
rect 146260 268348 498844 268376
rect 146260 268336 146266 268348
rect 498838 268336 498844 268348
rect 498896 268336 498902 268388
rect 137830 266976 137836 267028
rect 137888 267016 137894 267028
rect 185578 267016 185584 267028
rect 137888 266988 185584 267016
rect 137888 266976 137894 266988
rect 185578 266976 185584 266988
rect 185636 266976 185642 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 175918 266404 175924 266416
rect 3108 266376 175924 266404
rect 3108 266364 3114 266376
rect 175918 266364 175924 266376
rect 175976 266364 175982 266416
rect 140958 265684 140964 265736
rect 141016 265724 141022 265736
rect 180058 265724 180064 265736
rect 141016 265696 180064 265724
rect 141016 265684 141022 265696
rect 180058 265684 180064 265696
rect 180116 265684 180122 265736
rect 3418 265616 3424 265668
rect 3476 265656 3482 265668
rect 169202 265656 169208 265668
rect 3476 265628 169208 265656
rect 3476 265616 3482 265628
rect 169202 265616 169208 265628
rect 169260 265616 169266 265668
rect 174538 265548 174544 265600
rect 174596 265588 174602 265600
rect 174596 265560 180794 265588
rect 174596 265548 174602 265560
rect 180766 265520 180794 265560
rect 193582 265520 193588 265532
rect 180766 265492 193588 265520
rect 193582 265480 193588 265492
rect 193640 265480 193646 265532
rect 173434 265412 173440 265464
rect 173492 265452 173498 265464
rect 193766 265452 193772 265464
rect 173492 265424 193772 265452
rect 173492 265412 173498 265424
rect 193766 265412 193772 265424
rect 193824 265412 193830 265464
rect 170214 265344 170220 265396
rect 170272 265384 170278 265396
rect 170490 265384 170496 265396
rect 170272 265356 170496 265384
rect 170272 265344 170278 265356
rect 170490 265344 170496 265356
rect 170548 265384 170554 265396
rect 192018 265384 192024 265396
rect 170548 265356 192024 265384
rect 170548 265344 170554 265356
rect 192018 265344 192024 265356
rect 192076 265344 192082 265396
rect 175826 265276 175832 265328
rect 175884 265316 175890 265328
rect 197814 265316 197820 265328
rect 175884 265288 197820 265316
rect 175884 265276 175890 265288
rect 197814 265276 197820 265288
rect 197872 265276 197878 265328
rect 171686 265208 171692 265260
rect 171744 265248 171750 265260
rect 171870 265248 171876 265260
rect 171744 265220 171876 265248
rect 171744 265208 171750 265220
rect 171870 265208 171876 265220
rect 171928 265248 171934 265260
rect 194962 265248 194968 265260
rect 171928 265220 194968 265248
rect 171928 265208 171934 265220
rect 194962 265208 194968 265220
rect 195020 265208 195026 265260
rect 171778 265140 171784 265192
rect 171836 265180 171842 265192
rect 195146 265180 195152 265192
rect 171836 265152 195152 265180
rect 171836 265140 171842 265152
rect 195146 265140 195152 265152
rect 195204 265140 195210 265192
rect 170398 265072 170404 265124
rect 170456 265112 170462 265124
rect 170674 265112 170680 265124
rect 170456 265084 170680 265112
rect 170456 265072 170462 265084
rect 170674 265072 170680 265084
rect 170732 265112 170738 265124
rect 196250 265112 196256 265124
rect 170732 265084 196256 265112
rect 170732 265072 170738 265084
rect 196250 265072 196256 265084
rect 196308 265072 196314 265124
rect 169110 265004 169116 265056
rect 169168 265044 169174 265056
rect 197906 265044 197912 265056
rect 169168 265016 197912 265044
rect 169168 265004 169174 265016
rect 197906 265004 197912 265016
rect 197964 265004 197970 265056
rect 163498 264936 163504 264988
rect 163556 264976 163562 264988
rect 195054 264976 195060 264988
rect 163556 264948 195060 264976
rect 163556 264936 163562 264948
rect 195054 264936 195060 264948
rect 195112 264936 195118 264988
rect 149698 264324 149704 264376
rect 149756 264364 149762 264376
rect 173250 264364 173256 264376
rect 149756 264336 173256 264364
rect 149756 264324 149762 264336
rect 173250 264324 173256 264336
rect 173308 264324 173314 264376
rect 139394 264256 139400 264308
rect 139452 264296 139458 264308
rect 178678 264296 178684 264308
rect 139452 264268 178684 264296
rect 139452 264256 139458 264268
rect 178678 264256 178684 264268
rect 178736 264256 178742 264308
rect 106918 264188 106924 264240
rect 106976 264228 106982 264240
rect 158714 264228 158720 264240
rect 106976 264200 158720 264228
rect 106976 264188 106982 264200
rect 158714 264188 158720 264200
rect 158772 264188 158778 264240
rect 116946 264052 116952 264104
rect 117004 264092 117010 264104
rect 133138 264092 133144 264104
rect 117004 264064 133144 264092
rect 117004 264052 117010 264064
rect 133138 264052 133144 264064
rect 133196 264092 133202 264104
rect 133322 264092 133328 264104
rect 133196 264064 133328 264092
rect 133196 264052 133202 264064
rect 133322 264052 133328 264064
rect 133380 264052 133386 264104
rect 118326 263984 118332 264036
rect 118384 264024 118390 264036
rect 134242 264024 134248 264036
rect 118384 263996 134248 264024
rect 118384 263984 118390 263996
rect 134242 263984 134248 263996
rect 134300 264024 134306 264036
rect 134610 264024 134616 264036
rect 134300 263996 134616 264024
rect 134300 263984 134306 263996
rect 134610 263984 134616 263996
rect 134668 263984 134674 264036
rect 119706 263916 119712 263968
rect 119764 263956 119770 263968
rect 137830 263956 137836 263968
rect 119764 263928 137836 263956
rect 119764 263916 119770 263928
rect 137830 263916 137836 263928
rect 137888 263916 137894 263968
rect 120902 263848 120908 263900
rect 120960 263888 120966 263900
rect 139394 263888 139400 263900
rect 120960 263860 139400 263888
rect 120960 263848 120966 263860
rect 139394 263848 139400 263860
rect 139452 263848 139458 263900
rect 121730 263780 121736 263832
rect 121788 263820 121794 263832
rect 142614 263820 142620 263832
rect 121788 263792 142620 263820
rect 121788 263780 121794 263792
rect 142614 263780 142620 263792
rect 142672 263780 142678 263832
rect 120994 263712 121000 263764
rect 121052 263752 121058 263764
rect 140958 263752 140964 263764
rect 121052 263724 140964 263752
rect 121052 263712 121058 263724
rect 140958 263712 140964 263724
rect 141016 263712 141022 263764
rect 172698 263712 172704 263764
rect 172756 263752 172762 263764
rect 190822 263752 190828 263764
rect 172756 263724 190828 263752
rect 172756 263712 172762 263724
rect 190822 263712 190828 263724
rect 190880 263712 190886 263764
rect 114186 263644 114192 263696
rect 114244 263684 114250 263696
rect 137186 263684 137192 263696
rect 114244 263656 137192 263684
rect 114244 263644 114250 263656
rect 137186 263644 137192 263656
rect 137244 263644 137250 263696
rect 173250 263644 173256 263696
rect 173308 263684 173314 263696
rect 190914 263684 190920 263696
rect 173308 263656 190920 263684
rect 173308 263644 173314 263656
rect 190914 263644 190920 263656
rect 190972 263644 190978 263696
rect 121086 263576 121092 263628
rect 121144 263616 121150 263628
rect 151078 263616 151084 263628
rect 121144 263588 151084 263616
rect 121144 263576 121150 263588
rect 151078 263576 151084 263588
rect 151136 263576 151142 263628
rect 158714 263576 158720 263628
rect 158772 263616 158778 263628
rect 159358 263616 159364 263628
rect 158772 263588 159364 263616
rect 158772 263576 158778 263588
rect 159358 263576 159364 263588
rect 159416 263616 159422 263628
rect 187878 263616 187884 263628
rect 159416 263588 187884 263616
rect 159416 263576 159422 263588
rect 187878 263576 187884 263588
rect 187936 263576 187942 263628
rect 137462 263508 137468 263560
rect 137520 263548 137526 263560
rect 580258 263548 580264 263560
rect 137520 263520 580264 263548
rect 137520 263508 137526 263520
rect 580258 263508 580264 263520
rect 580316 263508 580322 263560
rect 150434 263440 150440 263492
rect 150492 263480 150498 263492
rect 151354 263480 151360 263492
rect 150492 263452 151360 263480
rect 150492 263440 150498 263452
rect 151354 263440 151360 263452
rect 151412 263440 151418 263492
rect 188522 263440 188528 263492
rect 188580 263480 188586 263492
rect 347774 263480 347780 263492
rect 188580 263452 347780 263480
rect 188580 263440 188586 263452
rect 347774 263440 347780 263452
rect 347832 263440 347838 263492
rect 193122 263372 193128 263424
rect 193180 263412 193186 263424
rect 218054 263412 218060 263424
rect 193180 263384 218060 263412
rect 193180 263372 193186 263384
rect 218054 263372 218060 263384
rect 218112 263372 218118 263424
rect 3510 263032 3516 263084
rect 3568 263072 3574 263084
rect 177390 263072 177396 263084
rect 3568 263044 177396 263072
rect 3568 263032 3574 263044
rect 177390 263032 177396 263044
rect 177448 263032 177454 263084
rect 132034 262964 132040 263016
rect 132092 263004 132098 263016
rect 580350 263004 580356 263016
rect 132092 262976 580356 263004
rect 132092 262964 132098 262976
rect 580350 262964 580356 262976
rect 580408 262964 580414 263016
rect 118418 262896 118424 262948
rect 118476 262936 118482 262948
rect 125962 262936 125968 262948
rect 118476 262908 125968 262936
rect 118476 262896 118482 262908
rect 125962 262896 125968 262908
rect 126020 262896 126026 262948
rect 131114 262896 131120 262948
rect 131172 262936 131178 262948
rect 131758 262936 131764 262948
rect 131172 262908 131764 262936
rect 131172 262896 131178 262908
rect 131758 262896 131764 262908
rect 131816 262936 131822 262948
rect 580442 262936 580448 262948
rect 131816 262908 580448 262936
rect 131816 262896 131822 262908
rect 580442 262896 580448 262908
rect 580500 262896 580506 262948
rect 3418 262828 3424 262880
rect 3476 262868 3482 262880
rect 179046 262868 179052 262880
rect 3476 262840 179052 262868
rect 3476 262828 3482 262840
rect 179046 262828 179052 262840
rect 179104 262828 179110 262880
rect 179230 262828 179236 262880
rect 179288 262868 179294 262880
rect 189626 262868 189632 262880
rect 179288 262840 189632 262868
rect 179288 262828 179294 262840
rect 189626 262828 189632 262840
rect 189684 262828 189690 262880
rect 282914 262868 282920 262880
rect 200086 262840 282920 262868
rect 116854 262760 116860 262812
rect 116912 262800 116918 262812
rect 131114 262800 131120 262812
rect 116912 262772 131120 262800
rect 116912 262760 116918 262772
rect 131114 262760 131120 262772
rect 131172 262760 131178 262812
rect 167822 262760 167828 262812
rect 167880 262800 167886 262812
rect 192386 262800 192392 262812
rect 167880 262772 192392 262800
rect 167880 262760 167886 262772
rect 192386 262760 192392 262772
rect 192444 262760 192450 262812
rect 116762 262692 116768 262744
rect 116820 262732 116826 262744
rect 134518 262732 134524 262744
rect 116820 262704 134524 262732
rect 116820 262692 116826 262704
rect 134518 262692 134524 262704
rect 134576 262732 134582 262744
rect 134794 262732 134800 262744
rect 134576 262704 134800 262732
rect 134576 262692 134582 262704
rect 134794 262692 134800 262704
rect 134852 262692 134858 262744
rect 153194 262692 153200 262744
rect 153252 262732 153258 262744
rect 158714 262732 158720 262744
rect 153252 262704 158720 262732
rect 153252 262692 153258 262704
rect 158714 262692 158720 262704
rect 158772 262692 158778 262744
rect 166258 262692 166264 262744
rect 166316 262732 166322 262744
rect 192202 262732 192208 262744
rect 166316 262704 192208 262732
rect 166316 262692 166322 262704
rect 192202 262692 192208 262704
rect 192260 262692 192266 262744
rect 114002 262624 114008 262676
rect 114060 262664 114066 262676
rect 128722 262664 128728 262676
rect 114060 262636 128728 262664
rect 114060 262624 114066 262636
rect 128722 262624 128728 262636
rect 128780 262624 128786 262676
rect 153838 262624 153844 262676
rect 153896 262664 153902 262676
rect 187970 262664 187976 262676
rect 153896 262636 187976 262664
rect 153896 262624 153902 262636
rect 187970 262624 187976 262636
rect 188028 262664 188034 262676
rect 188522 262664 188528 262676
rect 188028 262636 188528 262664
rect 188028 262624 188034 262636
rect 188522 262624 188528 262636
rect 188580 262624 188586 262676
rect 119798 262556 119804 262608
rect 119856 262596 119862 262608
rect 131114 262596 131120 262608
rect 119856 262568 131120 262596
rect 119856 262556 119862 262568
rect 131114 262556 131120 262568
rect 131172 262556 131178 262608
rect 155862 262556 155868 262608
rect 155920 262596 155926 262608
rect 191006 262596 191012 262608
rect 155920 262568 191012 262596
rect 155920 262556 155926 262568
rect 191006 262556 191012 262568
rect 191064 262596 191070 262608
rect 200086 262596 200114 262840
rect 282914 262828 282920 262840
rect 282972 262828 282978 262880
rect 191064 262568 200114 262596
rect 191064 262556 191070 262568
rect 122374 262488 122380 262540
rect 122432 262528 122438 262540
rect 152182 262528 152188 262540
rect 122432 262500 152188 262528
rect 122432 262488 122438 262500
rect 152182 262488 152188 262500
rect 152240 262528 152246 262540
rect 152458 262528 152464 262540
rect 152240 262500 152464 262528
rect 152240 262488 152246 262500
rect 152458 262488 152464 262500
rect 152516 262488 152522 262540
rect 157150 262488 157156 262540
rect 157208 262528 157214 262540
rect 192294 262528 192300 262540
rect 157208 262500 192300 262528
rect 157208 262488 157214 262500
rect 192294 262488 192300 262500
rect 192352 262528 192358 262540
rect 193122 262528 193128 262540
rect 192352 262500 193128 262528
rect 192352 262488 192358 262500
rect 193122 262488 193128 262500
rect 193180 262488 193186 262540
rect 118050 262420 118056 262472
rect 118108 262460 118114 262472
rect 129274 262460 129280 262472
rect 118108 262432 129280 262460
rect 118108 262420 118114 262432
rect 129274 262420 129280 262432
rect 129332 262420 129338 262472
rect 181438 262420 181444 262472
rect 181496 262460 181502 262472
rect 192110 262460 192116 262472
rect 181496 262432 192116 262460
rect 181496 262420 181502 262432
rect 192110 262420 192116 262432
rect 192168 262420 192174 262472
rect 119614 262352 119620 262404
rect 119672 262392 119678 262404
rect 127710 262392 127716 262404
rect 119672 262364 127716 262392
rect 119672 262352 119678 262364
rect 127710 262352 127716 262364
rect 127768 262352 127774 262404
rect 184750 262352 184756 262404
rect 184808 262392 184814 262404
rect 193674 262392 193680 262404
rect 184808 262364 193680 262392
rect 184808 262352 184814 262364
rect 193674 262352 193680 262364
rect 193732 262352 193738 262404
rect 113910 262284 113916 262336
rect 113968 262324 113974 262336
rect 127066 262324 127072 262336
rect 113968 262296 127072 262324
rect 113968 262284 113974 262296
rect 127066 262284 127072 262296
rect 127124 262284 127130 262336
rect 182910 262284 182916 262336
rect 182968 262324 182974 262336
rect 190454 262324 190460 262336
rect 182968 262296 190460 262324
rect 182968 262284 182974 262296
rect 190454 262284 190460 262296
rect 190512 262284 190518 262336
rect 181162 262216 181168 262268
rect 181220 262256 181226 262268
rect 187694 262256 187700 262268
rect 181220 262228 187700 262256
rect 181220 262216 181226 262228
rect 187694 262216 187700 262228
rect 187752 262216 187758 262268
rect 129826 261400 129832 261452
rect 129884 261440 129890 261452
rect 188338 261440 188344 261452
rect 129884 261412 188344 261440
rect 129884 261400 129890 261412
rect 188338 261400 188344 261412
rect 188396 261400 188402 261452
rect 179046 261332 179052 261384
rect 179104 261372 179110 261384
rect 198090 261372 198096 261384
rect 179104 261344 198096 261372
rect 179104 261332 179110 261344
rect 198090 261332 198096 261344
rect 198148 261332 198154 261384
rect 131114 261264 131120 261316
rect 131172 261304 131178 261316
rect 471238 261304 471244 261316
rect 131172 261276 471244 261304
rect 131172 261264 131178 261276
rect 471238 261264 471244 261276
rect 471296 261264 471302 261316
rect 177942 261196 177948 261248
rect 178000 261236 178006 261248
rect 191282 261236 191288 261248
rect 178000 261208 191288 261236
rect 178000 261196 178006 261208
rect 191282 261196 191288 261208
rect 191340 261196 191346 261248
rect 180702 261128 180708 261180
rect 180760 261168 180766 261180
rect 196710 261168 196716 261180
rect 180760 261140 196716 261168
rect 180760 261128 180766 261140
rect 196710 261128 196716 261140
rect 196768 261128 196774 261180
rect 120810 261060 120816 261112
rect 120868 261100 120874 261112
rect 133230 261100 133236 261112
rect 120868 261072 133236 261100
rect 120868 261060 120874 261072
rect 133230 261060 133236 261072
rect 133288 261060 133294 261112
rect 177390 261060 177396 261112
rect 177448 261100 177454 261112
rect 196526 261100 196532 261112
rect 177448 261072 196532 261100
rect 177448 261060 177454 261072
rect 196526 261060 196532 261072
rect 196584 261060 196590 261112
rect 115290 260992 115296 261044
rect 115348 261032 115354 261044
rect 130378 261032 130384 261044
rect 115348 261004 130384 261032
rect 115348 260992 115354 261004
rect 130378 260992 130384 261004
rect 130436 260992 130442 261044
rect 181990 260992 181996 261044
rect 182048 261032 182054 261044
rect 196434 261032 196440 261044
rect 182048 261004 196440 261032
rect 182048 260992 182054 261004
rect 196434 260992 196440 261004
rect 196492 260992 196498 261044
rect 14458 260924 14464 260976
rect 14516 260964 14522 260976
rect 176194 260964 176200 260976
rect 14516 260936 176200 260964
rect 14516 260924 14522 260936
rect 176194 260924 176200 260936
rect 176252 260964 176258 260976
rect 189718 260964 189724 260976
rect 176252 260936 189724 260964
rect 176252 260924 176258 260936
rect 189718 260924 189724 260936
rect 189776 260924 189782 260976
rect 115566 260856 115572 260908
rect 115624 260896 115630 260908
rect 132034 260896 132040 260908
rect 115624 260868 132040 260896
rect 115624 260856 115630 260868
rect 132034 260856 132040 260868
rect 132092 260856 132098 260908
rect 184014 260856 184020 260908
rect 184072 260896 184078 260908
rect 197998 260896 198004 260908
rect 184072 260868 198004 260896
rect 184072 260856 184078 260868
rect 197998 260856 198004 260868
rect 198056 260856 198062 260908
rect 118234 260788 118240 260840
rect 118292 260828 118298 260840
rect 124306 260828 124312 260840
rect 118292 260800 124312 260828
rect 118292 260788 118298 260800
rect 124306 260788 124312 260800
rect 124364 260788 124370 260840
rect 181254 260516 181260 260568
rect 181312 260556 181318 260568
rect 188062 260556 188068 260568
rect 181312 260528 188068 260556
rect 181312 260516 181318 260528
rect 188062 260516 188068 260528
rect 188120 260516 188126 260568
rect 179690 260448 179696 260500
rect 179748 260488 179754 260500
rect 192294 260488 192300 260500
rect 179748 260460 192300 260488
rect 179748 260448 179754 260460
rect 192294 260448 192300 260460
rect 192352 260448 192358 260500
rect 4798 260380 4804 260432
rect 4856 260420 4862 260432
rect 177942 260420 177948 260432
rect 4856 260392 177948 260420
rect 4856 260380 4862 260392
rect 177942 260380 177948 260392
rect 178000 260380 178006 260432
rect 178678 260380 178684 260432
rect 178736 260420 178742 260432
rect 191098 260420 191104 260432
rect 178736 260392 191104 260420
rect 178736 260380 178742 260392
rect 191098 260380 191104 260392
rect 191156 260380 191162 260432
rect 133230 260312 133236 260364
rect 133288 260352 133294 260364
rect 472618 260352 472624 260364
rect 133288 260324 178816 260352
rect 133288 260312 133294 260324
rect 169202 260244 169208 260296
rect 169260 260284 169266 260296
rect 178678 260284 178684 260296
rect 169260 260256 178684 260284
rect 169260 260244 169266 260256
rect 178678 260244 178684 260256
rect 178736 260244 178742 260296
rect 178788 260284 178816 260324
rect 183526 260324 472624 260352
rect 183526 260284 183554 260324
rect 472618 260312 472624 260324
rect 472676 260312 472682 260364
rect 178788 260256 183554 260284
rect 135254 260216 135260 260228
rect 122806 260188 135260 260216
rect 122190 260108 122196 260160
rect 122248 260148 122254 260160
rect 122806 260148 122834 260188
rect 135254 260176 135260 260188
rect 135312 260216 135318 260228
rect 136220 260216 136226 260228
rect 135312 260188 136226 260216
rect 135312 260176 135318 260188
rect 136220 260176 136226 260188
rect 136278 260176 136284 260228
rect 157334 260176 157340 260228
rect 157392 260216 157398 260228
rect 158300 260216 158306 260228
rect 157392 260188 158306 260216
rect 157392 260176 157398 260188
rect 158300 260176 158306 260188
rect 158358 260176 158364 260228
rect 166994 260176 167000 260228
rect 167052 260216 167058 260228
rect 167684 260216 167690 260228
rect 167052 260188 167690 260216
rect 167052 260176 167058 260188
rect 167684 260176 167690 260188
rect 167742 260176 167748 260228
rect 169754 260176 169760 260228
rect 169812 260216 169818 260228
rect 170996 260216 171002 260228
rect 169812 260188 171002 260216
rect 169812 260176 169818 260188
rect 170996 260176 171002 260188
rect 171054 260216 171060 260228
rect 189350 260216 189356 260228
rect 171054 260188 189356 260216
rect 171054 260176 171060 260188
rect 189350 260176 189356 260188
rect 189408 260176 189414 260228
rect 122248 260120 122834 260148
rect 122248 260108 122254 260120
rect 175918 260108 175924 260160
rect 175976 260148 175982 260160
rect 189534 260148 189540 260160
rect 175976 260120 189540 260148
rect 175976 260108 175982 260120
rect 189534 260108 189540 260120
rect 189592 260108 189598 260160
rect 115474 260040 115480 260092
rect 115532 260080 115538 260092
rect 126836 260080 126842 260092
rect 115532 260052 126842 260080
rect 115532 260040 115538 260052
rect 126836 260040 126842 260052
rect 126894 260040 126900 260092
rect 167684 260040 167690 260092
rect 167742 260080 167748 260092
rect 189442 260080 189448 260092
rect 167742 260052 171134 260080
rect 167742 260040 167748 260052
rect 118142 259972 118148 260024
rect 118200 260012 118206 260024
rect 139670 260012 139676 260024
rect 118200 259984 139676 260012
rect 118200 259972 118206 259984
rect 139670 259972 139676 259984
rect 139728 259972 139734 260024
rect 171106 260012 171134 260052
rect 176626 260052 189448 260080
rect 176626 260012 176654 260052
rect 189442 260040 189448 260052
rect 189500 260040 189506 260092
rect 171106 259984 176654 260012
rect 178494 259972 178500 260024
rect 178552 260012 178558 260024
rect 181622 260012 181628 260024
rect 178552 259984 181628 260012
rect 178552 259972 178558 259984
rect 181622 259972 181628 259984
rect 181680 259972 181686 260024
rect 181714 259972 181720 260024
rect 181772 260012 181778 260024
rect 184658 260012 184664 260024
rect 181772 259984 184664 260012
rect 181772 259972 181778 259984
rect 184658 259972 184664 259984
rect 184716 259972 184722 260024
rect 187970 260012 187976 260024
rect 186286 259984 187976 260012
rect 119522 259904 119528 259956
rect 119580 259944 119586 259956
rect 140774 259944 140780 259956
rect 119580 259916 140780 259944
rect 119580 259904 119586 259916
rect 140774 259904 140780 259916
rect 140832 259944 140838 259956
rect 141418 259944 141424 259956
rect 140832 259916 141424 259944
rect 140832 259904 140838 259916
rect 141418 259904 141424 259916
rect 141476 259904 141482 259956
rect 164694 259904 164700 259956
rect 164752 259944 164758 259956
rect 186286 259944 186314 259984
rect 187970 259972 187976 259984
rect 188028 259972 188034 260024
rect 164752 259916 186314 259944
rect 164752 259904 164758 259916
rect 121914 259836 121920 259888
rect 121972 259876 121978 259888
rect 146294 259876 146300 259888
rect 121972 259848 146300 259876
rect 121972 259836 121978 259848
rect 146294 259836 146300 259848
rect 146352 259836 146358 259888
rect 166166 259836 166172 259888
rect 166224 259876 166230 259888
rect 191190 259876 191196 259888
rect 166224 259848 191196 259876
rect 166224 259836 166230 259848
rect 191190 259836 191196 259848
rect 191248 259836 191254 259888
rect 121178 259768 121184 259820
rect 121236 259808 121242 259820
rect 147674 259808 147680 259820
rect 121236 259780 147680 259808
rect 121236 259768 121242 259780
rect 147674 259768 147680 259780
rect 147732 259768 147738 259820
rect 158070 259768 158076 259820
rect 158128 259808 158134 259820
rect 181254 259808 181260 259820
rect 158128 259780 181260 259808
rect 158128 259768 158134 259780
rect 181254 259768 181260 259780
rect 181312 259768 181318 259820
rect 181622 259768 181628 259820
rect 181680 259808 181686 259820
rect 188246 259808 188252 259820
rect 181680 259780 188252 259808
rect 181680 259768 181686 259780
rect 188246 259768 188252 259780
rect 188304 259768 188310 259820
rect 119430 259700 119436 259752
rect 119488 259740 119494 259752
rect 153194 259740 153200 259752
rect 119488 259712 153200 259740
rect 119488 259700 119494 259712
rect 153194 259700 153200 259712
rect 153252 259700 153258 259752
rect 158622 259700 158628 259752
rect 158680 259740 158686 259752
rect 179690 259740 179696 259752
rect 158680 259712 179696 259740
rect 158680 259700 158686 259712
rect 179690 259700 179696 259712
rect 179748 259700 179754 259752
rect 180150 259700 180156 259752
rect 180208 259740 180214 259752
rect 180208 259712 184244 259740
rect 180208 259700 180214 259712
rect 134334 259632 134340 259684
rect 134392 259672 134398 259684
rect 134392 259644 181852 259672
rect 134392 259632 134398 259644
rect 120626 259564 120632 259616
rect 120684 259604 120690 259616
rect 178034 259604 178040 259616
rect 120684 259576 178040 259604
rect 120684 259564 120690 259576
rect 178034 259564 178040 259576
rect 178092 259564 178098 259616
rect 181714 259604 181720 259616
rect 181456 259576 181720 259604
rect 120718 259496 120724 259548
rect 120776 259536 120782 259548
rect 125594 259536 125600 259548
rect 120776 259508 125600 259536
rect 120776 259496 120782 259508
rect 125594 259496 125600 259508
rect 125652 259496 125658 259548
rect 174446 259496 174452 259548
rect 174504 259536 174510 259548
rect 181456 259536 181484 259576
rect 181714 259564 181720 259576
rect 181772 259564 181778 259616
rect 174504 259508 181484 259536
rect 174504 259496 174510 259508
rect 116670 259428 116676 259480
rect 116728 259468 116734 259480
rect 128354 259468 128360 259480
rect 116728 259440 128360 259468
rect 116728 259428 116734 259440
rect 128354 259428 128360 259440
rect 128412 259428 128418 259480
rect 181824 259468 181852 259644
rect 184216 259604 184244 259712
rect 184566 259700 184572 259752
rect 184624 259740 184630 259752
rect 190546 259740 190552 259752
rect 184624 259712 190552 259740
rect 184624 259700 184630 259712
rect 190546 259700 190552 259712
rect 190604 259700 190610 259752
rect 184658 259632 184664 259684
rect 184716 259672 184722 259684
rect 187326 259672 187332 259684
rect 184716 259644 187332 259672
rect 184716 259632 184722 259644
rect 187326 259632 187332 259644
rect 187384 259632 187390 259684
rect 187234 259604 187240 259616
rect 184216 259576 187240 259604
rect 187234 259564 187240 259576
rect 187292 259564 187298 259616
rect 183462 259496 183468 259548
rect 183520 259536 183526 259548
rect 195238 259536 195244 259548
rect 183520 259508 195244 259536
rect 183520 259496 183526 259508
rect 195238 259496 195244 259508
rect 195296 259496 195302 259548
rect 181824 259440 190454 259468
rect 190426 259400 190454 259440
rect 580166 259400 580172 259412
rect 190426 259372 580172 259400
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 472618 245556 472624 245608
rect 472676 245596 472682 245608
rect 580166 245596 580172 245608
rect 472676 245568 580172 245596
rect 472676 245556 472682 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 14458 241448 14464 241460
rect 3568 241420 14464 241448
rect 3568 241408 3574 241420
rect 14458 241408 14464 241420
rect 14516 241408 14522 241460
rect 2774 215228 2780 215280
rect 2832 215268 2838 215280
rect 4798 215268 4804 215280
rect 2832 215240 4804 215268
rect 2832 215228 2838 215240
rect 4798 215228 4804 215240
rect 4856 215228 4862 215280
rect 471238 206932 471244 206984
rect 471296 206972 471302 206984
rect 579798 206972 579804 206984
rect 471296 206944 579804 206972
rect 471296 206932 471302 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 154270 201028 179414 201056
rect 135226 200756 150434 200784
rect 111702 200608 111708 200660
rect 111760 200648 111766 200660
rect 131942 200648 131948 200660
rect 111760 200620 131948 200648
rect 111760 200608 111766 200620
rect 131942 200608 131948 200620
rect 132000 200608 132006 200660
rect 115842 200540 115848 200592
rect 115900 200580 115906 200592
rect 135226 200580 135254 200756
rect 115900 200552 135254 200580
rect 135318 200688 149882 200716
rect 115900 200540 115906 200552
rect 122742 200472 122748 200524
rect 122800 200512 122806 200524
rect 135318 200512 135346 200688
rect 122800 200484 135346 200512
rect 122800 200472 122806 200484
rect 112990 200404 112996 200456
rect 113048 200444 113054 200456
rect 132034 200444 132040 200456
rect 113048 200416 132040 200444
rect 113048 200404 113054 200416
rect 132034 200404 132040 200416
rect 132092 200404 132098 200456
rect 132144 200416 135346 200444
rect 107194 200336 107200 200388
rect 107252 200376 107258 200388
rect 132144 200376 132172 200416
rect 107252 200348 132172 200376
rect 107252 200336 107258 200348
rect 113082 200268 113088 200320
rect 113140 200308 113146 200320
rect 130930 200308 130936 200320
rect 113140 200280 130936 200308
rect 113140 200268 113146 200280
rect 130930 200268 130936 200280
rect 130988 200268 130994 200320
rect 122558 200132 122564 200184
rect 122616 200172 122622 200184
rect 135318 200172 135346 200416
rect 122616 200144 135208 200172
rect 135318 200144 136910 200172
rect 122616 200132 122622 200144
rect 125594 200064 125600 200116
rect 125652 200104 125658 200116
rect 125652 200076 134058 200104
rect 125652 200064 125658 200076
rect 125226 199928 125232 199980
rect 125284 199968 125290 199980
rect 125284 199940 133782 199968
rect 125284 199928 125290 199940
rect 133754 199912 133782 199940
rect 134030 199912 134058 200076
rect 135180 199912 135208 200144
rect 136882 199912 136910 200144
rect 136974 199940 140498 199968
rect 127526 199860 127532 199912
rect 127584 199900 127590 199912
rect 132908 199900 132914 199912
rect 127584 199872 132914 199900
rect 127584 199860 127590 199872
rect 132908 199860 132914 199872
rect 132966 199860 132972 199912
rect 133092 199860 133098 199912
rect 133150 199860 133156 199912
rect 133184 199860 133190 199912
rect 133242 199860 133248 199912
rect 133460 199860 133466 199912
rect 133518 199860 133524 199912
rect 133736 199860 133742 199912
rect 133794 199860 133800 199912
rect 134012 199860 134018 199912
rect 134070 199860 134076 199912
rect 134104 199860 134110 199912
rect 134162 199860 134168 199912
rect 134472 199900 134478 199912
rect 134444 199860 134478 199900
rect 134530 199860 134536 199912
rect 134564 199860 134570 199912
rect 134622 199860 134628 199912
rect 134656 199860 134662 199912
rect 134714 199860 134720 199912
rect 135180 199872 135214 199912
rect 135208 199860 135214 199872
rect 135266 199860 135272 199912
rect 135484 199860 135490 199912
rect 135542 199900 135548 199912
rect 135542 199860 135576 199900
rect 135668 199860 135674 199912
rect 135726 199860 135732 199912
rect 136036 199860 136042 199912
rect 136094 199860 136100 199912
rect 136312 199860 136318 199912
rect 136370 199860 136376 199912
rect 136496 199860 136502 199912
rect 136554 199860 136560 199912
rect 136680 199860 136686 199912
rect 136738 199860 136744 199912
rect 136864 199860 136870 199912
rect 136922 199860 136928 199912
rect 132862 199724 132868 199776
rect 132920 199764 132926 199776
rect 133110 199764 133138 199860
rect 132920 199736 133138 199764
rect 132920 199724 132926 199736
rect 111242 199656 111248 199708
rect 111300 199696 111306 199708
rect 128814 199696 128820 199708
rect 111300 199668 128820 199696
rect 111300 199656 111306 199668
rect 128814 199656 128820 199668
rect 128872 199656 128878 199708
rect 133202 199640 133230 199860
rect 133276 199792 133282 199844
rect 133334 199832 133340 199844
rect 133334 199792 133368 199832
rect 133340 199708 133368 199792
rect 133478 199708 133506 199860
rect 133322 199656 133328 199708
rect 133380 199656 133386 199708
rect 133414 199656 133420 199708
rect 133472 199668 133506 199708
rect 133472 199656 133478 199668
rect 134122 199640 134150 199860
rect 111518 199588 111524 199640
rect 111576 199628 111582 199640
rect 131574 199628 131580 199640
rect 111576 199600 131580 199628
rect 111576 199588 111582 199600
rect 131574 199588 131580 199600
rect 131632 199588 131638 199640
rect 133138 199588 133144 199640
rect 133196 199600 133230 199640
rect 133196 199588 133202 199600
rect 134058 199588 134064 199640
rect 134116 199600 134150 199640
rect 134444 199628 134472 199860
rect 134582 199832 134610 199860
rect 134536 199804 134610 199832
rect 134536 199776 134564 199804
rect 134674 199776 134702 199860
rect 135548 199776 135576 199860
rect 135686 199832 135714 199860
rect 135640 199804 135714 199832
rect 134518 199724 134524 199776
rect 134576 199724 134582 199776
rect 134610 199724 134616 199776
rect 134668 199736 134702 199776
rect 134668 199724 134674 199736
rect 135530 199724 135536 199776
rect 135588 199724 135594 199776
rect 135640 199708 135668 199804
rect 135622 199656 135628 199708
rect 135680 199656 135686 199708
rect 134702 199628 134708 199640
rect 134444 199600 134708 199628
rect 134116 199588 134122 199600
rect 134702 199588 134708 199600
rect 134760 199588 134766 199640
rect 135346 199588 135352 199640
rect 135404 199628 135410 199640
rect 136054 199628 136082 199860
rect 135404 199600 136082 199628
rect 135404 199588 135410 199600
rect 136174 199588 136180 199640
rect 136232 199628 136238 199640
rect 136330 199628 136358 199860
rect 136514 199696 136542 199860
rect 136698 199776 136726 199860
rect 136698 199736 136732 199776
rect 136726 199724 136732 199736
rect 136784 199724 136790 199776
rect 136818 199724 136824 199776
rect 136876 199764 136882 199776
rect 136974 199764 137002 199940
rect 140470 199912 140498 199940
rect 141298 199940 142292 199968
rect 141298 199912 141326 199940
rect 137048 199860 137054 199912
rect 137106 199860 137112 199912
rect 137416 199860 137422 199912
rect 137474 199860 137480 199912
rect 137784 199860 137790 199912
rect 137842 199860 137848 199912
rect 138244 199860 138250 199912
rect 138302 199860 138308 199912
rect 138336 199860 138342 199912
rect 138394 199860 138400 199912
rect 138520 199860 138526 199912
rect 138578 199860 138584 199912
rect 138796 199860 138802 199912
rect 138854 199860 138860 199912
rect 139072 199900 139078 199912
rect 138952 199872 139078 199900
rect 136876 199736 137002 199764
rect 136876 199724 136882 199736
rect 136468 199668 136542 199696
rect 137066 199708 137094 199860
rect 137232 199792 137238 199844
rect 137290 199792 137296 199844
rect 137250 199708 137278 199792
rect 137066 199668 137100 199708
rect 136468 199640 136496 199668
rect 137094 199656 137100 199668
rect 137152 199656 137158 199708
rect 137186 199656 137192 199708
rect 137244 199668 137278 199708
rect 137244 199656 137250 199668
rect 136232 199600 136358 199628
rect 136232 199588 136238 199600
rect 136450 199588 136456 199640
rect 136508 199588 136514 199640
rect 136542 199588 136548 199640
rect 136600 199628 136606 199640
rect 137434 199628 137462 199860
rect 137802 199776 137830 199860
rect 138262 199776 138290 199860
rect 137802 199736 137836 199776
rect 137830 199724 137836 199736
rect 137888 199724 137894 199776
rect 138198 199724 138204 199776
rect 138256 199736 138290 199776
rect 138256 199724 138262 199736
rect 136600 199600 137462 199628
rect 136600 199588 136606 199600
rect 138198 199588 138204 199640
rect 138256 199628 138262 199640
rect 138354 199628 138382 199860
rect 138538 199640 138566 199860
rect 138256 199600 138382 199628
rect 138256 199588 138262 199600
rect 138474 199588 138480 199640
rect 138532 199600 138566 199640
rect 138532 199588 138538 199600
rect 138658 199588 138664 199640
rect 138716 199628 138722 199640
rect 138814 199628 138842 199860
rect 138952 199640 138980 199872
rect 139072 199860 139078 199872
rect 139130 199860 139136 199912
rect 139164 199860 139170 199912
rect 139222 199860 139228 199912
rect 139256 199860 139262 199912
rect 139314 199860 139320 199912
rect 139348 199860 139354 199912
rect 139406 199860 139412 199912
rect 139900 199860 139906 199912
rect 139958 199860 139964 199912
rect 140084 199860 140090 199912
rect 140142 199860 140148 199912
rect 140268 199860 140274 199912
rect 140326 199860 140332 199912
rect 140452 199860 140458 199912
rect 140510 199860 140516 199912
rect 140820 199860 140826 199912
rect 140878 199860 140884 199912
rect 140912 199860 140918 199912
rect 140970 199860 140976 199912
rect 141004 199860 141010 199912
rect 141062 199860 141068 199912
rect 141096 199860 141102 199912
rect 141154 199860 141160 199912
rect 141188 199860 141194 199912
rect 141246 199860 141252 199912
rect 141280 199860 141286 199912
rect 141338 199860 141344 199912
rect 141372 199860 141378 199912
rect 141430 199860 141436 199912
rect 141556 199900 141562 199912
rect 141528 199860 141562 199900
rect 141614 199860 141620 199912
rect 141648 199860 141654 199912
rect 141706 199860 141712 199912
rect 141740 199860 141746 199912
rect 141798 199860 141804 199912
rect 141832 199860 141838 199912
rect 141890 199860 141896 199912
rect 139182 199832 139210 199860
rect 139044 199804 139210 199832
rect 138716 199600 138842 199628
rect 138716 199588 138722 199600
rect 138934 199588 138940 199640
rect 138992 199588 138998 199640
rect 139044 199628 139072 199804
rect 139118 199724 139124 199776
rect 139176 199764 139182 199776
rect 139274 199764 139302 199860
rect 139176 199736 139302 199764
rect 139176 199724 139182 199736
rect 139210 199656 139216 199708
rect 139268 199696 139274 199708
rect 139366 199696 139394 199860
rect 139268 199668 139394 199696
rect 139268 199656 139274 199668
rect 139918 199640 139946 199860
rect 139302 199628 139308 199640
rect 139044 199600 139308 199628
rect 139302 199588 139308 199600
rect 139360 199588 139366 199640
rect 139918 199600 139952 199640
rect 139946 199588 139952 199600
rect 140004 199588 140010 199640
rect 140102 199628 140130 199860
rect 140286 199708 140314 199860
rect 140360 199792 140366 199844
rect 140418 199832 140424 199844
rect 140636 199832 140642 199844
rect 140418 199792 140452 199832
rect 140424 199708 140452 199792
rect 140608 199792 140642 199832
rect 140694 199792 140700 199844
rect 140728 199792 140734 199844
rect 140786 199792 140792 199844
rect 140286 199668 140320 199708
rect 140314 199656 140320 199668
rect 140372 199656 140378 199708
rect 140406 199656 140412 199708
rect 140464 199656 140470 199708
rect 140608 199640 140636 199792
rect 140746 199696 140774 199792
rect 140700 199668 140774 199696
rect 140700 199640 140728 199668
rect 140838 199640 140866 199860
rect 140930 199776 140958 199860
rect 140912 199724 140918 199776
rect 140970 199724 140976 199776
rect 141022 199640 141050 199860
rect 141114 199708 141142 199860
rect 141206 199708 141234 199860
rect 141096 199656 141102 199708
rect 141154 199656 141160 199708
rect 141206 199668 141240 199708
rect 141234 199656 141240 199668
rect 141292 199656 141298 199708
rect 141390 199640 141418 199860
rect 140222 199628 140228 199640
rect 140102 199600 140228 199628
rect 140222 199588 140228 199600
rect 140280 199588 140286 199640
rect 140590 199588 140596 199640
rect 140648 199588 140654 199640
rect 140682 199588 140688 199640
rect 140740 199588 140746 199640
rect 140774 199588 140780 199640
rect 140832 199600 140866 199640
rect 140832 199588 140838 199600
rect 141004 199588 141010 199640
rect 141062 199588 141068 199640
rect 141390 199600 141424 199640
rect 141418 199588 141424 199600
rect 141476 199588 141482 199640
rect 141528 199628 141556 199860
rect 141666 199832 141694 199860
rect 141620 199804 141694 199832
rect 141620 199776 141648 199804
rect 141758 199776 141786 199860
rect 141602 199724 141608 199776
rect 141660 199724 141666 199776
rect 141694 199724 141700 199776
rect 141752 199736 141786 199776
rect 141752 199724 141758 199736
rect 141850 199708 141878 199860
rect 141786 199656 141792 199708
rect 141844 199668 141878 199708
rect 141844 199656 141850 199668
rect 142264 199640 142292 199940
rect 146082 199940 146294 199968
rect 146082 199912 146110 199940
rect 142384 199860 142390 199912
rect 142442 199860 142448 199912
rect 142568 199900 142574 199912
rect 142540 199860 142574 199900
rect 142626 199860 142632 199912
rect 142660 199860 142666 199912
rect 142718 199860 142724 199912
rect 142752 199860 142758 199912
rect 142810 199860 142816 199912
rect 142936 199860 142942 199912
rect 142994 199860 143000 199912
rect 143304 199860 143310 199912
rect 143362 199860 143368 199912
rect 143396 199860 143402 199912
rect 143454 199860 143460 199912
rect 143856 199860 143862 199912
rect 143914 199860 143920 199912
rect 143948 199860 143954 199912
rect 144006 199860 144012 199912
rect 144592 199860 144598 199912
rect 144650 199860 144656 199912
rect 144684 199860 144690 199912
rect 144742 199860 144748 199912
rect 144960 199860 144966 199912
rect 145018 199860 145024 199912
rect 145236 199860 145242 199912
rect 145294 199860 145300 199912
rect 145328 199860 145334 199912
rect 145386 199860 145392 199912
rect 145420 199860 145426 199912
rect 145478 199860 145484 199912
rect 145604 199860 145610 199912
rect 145662 199860 145668 199912
rect 146064 199860 146070 199912
rect 146122 199860 146128 199912
rect 146156 199860 146162 199912
rect 146214 199860 146220 199912
rect 142402 199776 142430 199860
rect 142402 199736 142436 199776
rect 142430 199724 142436 199736
rect 142488 199724 142494 199776
rect 142540 199708 142568 199860
rect 142678 199832 142706 199860
rect 142632 199804 142706 199832
rect 142632 199708 142660 199804
rect 142770 199776 142798 199860
rect 142706 199724 142712 199776
rect 142764 199736 142798 199776
rect 142764 199724 142770 199736
rect 142522 199656 142528 199708
rect 142580 199656 142586 199708
rect 142614 199656 142620 199708
rect 142672 199656 142678 199708
rect 142954 199640 142982 199860
rect 143322 199708 143350 199860
rect 143414 199764 143442 199860
rect 143414 199736 143488 199764
rect 143460 199708 143488 199736
rect 143322 199668 143356 199708
rect 143350 199656 143356 199668
rect 143408 199656 143414 199708
rect 143442 199656 143448 199708
rect 143500 199656 143506 199708
rect 141970 199628 141976 199640
rect 141528 199600 141976 199628
rect 141970 199588 141976 199600
rect 142028 199588 142034 199640
rect 142246 199588 142252 199640
rect 142304 199588 142310 199640
rect 142890 199588 142896 199640
rect 142948 199600 142982 199640
rect 143874 199640 143902 199860
rect 143966 199696 143994 199860
rect 144610 199832 144638 199860
rect 144288 199804 144638 199832
rect 143966 199668 144040 199696
rect 144012 199640 144040 199668
rect 144086 199656 144092 199708
rect 144144 199656 144150 199708
rect 143874 199600 143908 199640
rect 142948 199588 142954 199600
rect 143902 199588 143908 199600
rect 143960 199588 143966 199640
rect 143994 199588 144000 199640
rect 144052 199588 144058 199640
rect 144104 199572 144132 199656
rect 115658 199520 115664 199572
rect 115716 199560 115722 199572
rect 143626 199560 143632 199572
rect 115716 199532 143632 199560
rect 115716 199520 115722 199532
rect 143626 199520 143632 199532
rect 143684 199520 143690 199572
rect 144086 199520 144092 199572
rect 144144 199520 144150 199572
rect 144288 199560 144316 199804
rect 144702 199776 144730 199860
rect 144638 199724 144644 199776
rect 144696 199736 144730 199776
rect 144696 199724 144702 199736
rect 144978 199708 145006 199860
rect 144914 199656 144920 199708
rect 144972 199668 145006 199708
rect 145254 199708 145282 199860
rect 145346 199776 145374 199860
rect 145438 199832 145466 199860
rect 145438 199804 145512 199832
rect 145346 199736 145380 199776
rect 145374 199724 145380 199736
rect 145432 199724 145438 199776
rect 145254 199668 145288 199708
rect 144972 199656 144978 199668
rect 145282 199656 145288 199668
rect 145340 199656 145346 199708
rect 144362 199588 144368 199640
rect 144420 199628 144426 199640
rect 145484 199628 145512 199804
rect 145622 199776 145650 199860
rect 146174 199776 146202 199860
rect 145558 199724 145564 199776
rect 145616 199736 145650 199776
rect 145616 199724 145622 199736
rect 146110 199724 146116 199776
rect 146168 199736 146202 199776
rect 146168 199724 146174 199736
rect 144420 199600 145512 199628
rect 144420 199588 144426 199600
rect 146018 199588 146024 199640
rect 146076 199628 146082 199640
rect 146266 199628 146294 199940
rect 149118 199940 149514 199968
rect 149118 199912 149146 199940
rect 146432 199860 146438 199912
rect 146490 199860 146496 199912
rect 146616 199860 146622 199912
rect 146674 199860 146680 199912
rect 146892 199860 146898 199912
rect 146950 199860 146956 199912
rect 147076 199860 147082 199912
rect 147134 199860 147140 199912
rect 147168 199860 147174 199912
rect 147226 199860 147232 199912
rect 147352 199860 147358 199912
rect 147410 199860 147416 199912
rect 147628 199860 147634 199912
rect 147686 199860 147692 199912
rect 147812 199860 147818 199912
rect 147870 199860 147876 199912
rect 148088 199860 148094 199912
rect 148146 199860 148152 199912
rect 148272 199860 148278 199912
rect 148330 199860 148336 199912
rect 148456 199860 148462 199912
rect 148514 199860 148520 199912
rect 148732 199860 148738 199912
rect 148790 199860 148796 199912
rect 148824 199860 148830 199912
rect 148882 199860 148888 199912
rect 148916 199860 148922 199912
rect 148974 199860 148980 199912
rect 149100 199860 149106 199912
rect 149158 199860 149164 199912
rect 149376 199860 149382 199912
rect 149434 199860 149440 199912
rect 146076 199600 146294 199628
rect 146076 199588 146082 199600
rect 144822 199560 144828 199572
rect 144288 199532 144828 199560
rect 144822 199520 144828 199532
rect 144880 199520 144886 199572
rect 145098 199520 145104 199572
rect 145156 199560 145162 199572
rect 146450 199560 146478 199860
rect 146634 199640 146662 199860
rect 146570 199588 146576 199640
rect 146628 199600 146662 199640
rect 146910 199640 146938 199860
rect 147094 199640 147122 199860
rect 147186 199696 147214 199860
rect 147370 199764 147398 199860
rect 147370 199736 147444 199764
rect 147186 199668 147352 199696
rect 147324 199640 147352 199668
rect 146910 199600 146944 199640
rect 146628 199588 146634 199600
rect 146938 199588 146944 199600
rect 146996 199588 147002 199640
rect 147030 199588 147036 199640
rect 147088 199600 147122 199640
rect 147088 199588 147094 199600
rect 147306 199588 147312 199640
rect 147364 199588 147370 199640
rect 145156 199532 146478 199560
rect 145156 199520 145162 199532
rect 112806 199452 112812 199504
rect 112864 199492 112870 199504
rect 147416 199492 147444 199736
rect 147646 199572 147674 199860
rect 147830 199640 147858 199860
rect 148106 199776 148134 199860
rect 148042 199724 148048 199776
rect 148100 199736 148134 199776
rect 148100 199724 148106 199736
rect 148290 199640 148318 199860
rect 148474 199640 148502 199860
rect 148750 199832 148778 199860
rect 148704 199804 148778 199832
rect 148704 199776 148732 199804
rect 148842 199776 148870 199860
rect 148686 199724 148692 199776
rect 148744 199724 148750 199776
rect 148778 199724 148784 199776
rect 148836 199736 148870 199776
rect 148836 199724 148842 199736
rect 148934 199640 148962 199860
rect 149394 199696 149422 199860
rect 149486 199832 149514 199940
rect 149854 199912 149882 200688
rect 150406 199912 150434 200756
rect 150498 199940 150802 199968
rect 149560 199860 149566 199912
rect 149618 199900 149624 199912
rect 149618 199872 149790 199900
rect 149618 199860 149624 199872
rect 149486 199804 149652 199832
rect 149624 199776 149652 199804
rect 149606 199724 149612 199776
rect 149664 199724 149670 199776
rect 147766 199588 147772 199640
rect 147824 199600 147858 199640
rect 147824 199588 147830 199600
rect 148226 199588 148232 199640
rect 148284 199600 148318 199640
rect 148284 199588 148290 199600
rect 148410 199588 148416 199640
rect 148468 199600 148502 199640
rect 148468 199588 148474 199600
rect 148870 199588 148876 199640
rect 148928 199600 148962 199640
rect 149164 199668 149422 199696
rect 148928 199588 148934 199600
rect 147582 199520 147588 199572
rect 147640 199532 147674 199572
rect 147640 199520 147646 199532
rect 112864 199464 147444 199492
rect 149164 199492 149192 199668
rect 149762 199628 149790 199872
rect 149836 199860 149842 199912
rect 149894 199860 149900 199912
rect 149928 199860 149934 199912
rect 149986 199860 149992 199912
rect 150112 199860 150118 199912
rect 150170 199860 150176 199912
rect 150296 199860 150302 199912
rect 150354 199860 150360 199912
rect 150388 199860 150394 199912
rect 150446 199860 150452 199912
rect 149946 199776 149974 199860
rect 150130 199776 150158 199860
rect 149882 199724 149888 199776
rect 149940 199736 149974 199776
rect 149940 199724 149946 199736
rect 150066 199724 150072 199776
rect 150124 199736 150158 199776
rect 150124 199724 150130 199736
rect 150314 199708 150342 199860
rect 150314 199668 150348 199708
rect 150342 199656 150348 199668
rect 150400 199656 150406 199708
rect 150250 199628 150256 199640
rect 149762 199600 150256 199628
rect 150250 199588 150256 199600
rect 150308 199588 150314 199640
rect 150066 199520 150072 199572
rect 150124 199560 150130 199572
rect 150498 199560 150526 199940
rect 150774 199912 150802 199940
rect 151648 199940 152182 199968
rect 150664 199900 150670 199912
rect 150124 199532 150526 199560
rect 150636 199860 150670 199900
rect 150722 199860 150728 199912
rect 150756 199860 150762 199912
rect 150814 199860 150820 199912
rect 150848 199860 150854 199912
rect 150906 199860 150912 199912
rect 150940 199860 150946 199912
rect 150998 199860 151004 199912
rect 151216 199860 151222 199912
rect 151274 199860 151280 199912
rect 151308 199860 151314 199912
rect 151366 199860 151372 199912
rect 151400 199860 151406 199912
rect 151458 199860 151464 199912
rect 150124 199520 150130 199532
rect 149238 199492 149244 199504
rect 149164 199464 149244 199492
rect 112864 199452 112870 199464
rect 149238 199452 149244 199464
rect 149296 199452 149302 199504
rect 150636 199492 150664 199860
rect 150866 199832 150894 199860
rect 150728 199804 150894 199832
rect 150728 199776 150756 199804
rect 150710 199724 150716 199776
rect 150768 199724 150774 199776
rect 150958 199628 150986 199860
rect 151234 199708 151262 199860
rect 151170 199656 151176 199708
rect 151228 199668 151262 199708
rect 151228 199656 151234 199668
rect 151078 199628 151084 199640
rect 150958 199600 151084 199628
rect 151078 199588 151084 199600
rect 151136 199588 151142 199640
rect 151326 199572 151354 199860
rect 151418 199628 151446 199860
rect 151538 199628 151544 199640
rect 151418 199600 151544 199628
rect 151538 199588 151544 199600
rect 151596 199588 151602 199640
rect 151326 199532 151360 199572
rect 151354 199520 151360 199532
rect 151412 199520 151418 199572
rect 151262 199492 151268 199504
rect 150636 199464 151268 199492
rect 151262 199452 151268 199464
rect 151320 199452 151326 199504
rect 151648 199492 151676 199940
rect 152154 199912 152182 199940
rect 154270 199912 154298 201028
rect 162826 200892 163866 200920
rect 162826 200240 162854 200892
rect 163838 200648 163866 200892
rect 177850 200648 177856 200660
rect 163838 200620 177856 200648
rect 177850 200608 177856 200620
rect 177908 200608 177914 200660
rect 179386 200648 179414 201028
rect 180058 200648 180064 200660
rect 179386 200620 180064 200648
rect 180058 200608 180064 200620
rect 180116 200608 180122 200660
rect 183830 200540 183836 200592
rect 183888 200580 183894 200592
rect 186866 200580 186872 200592
rect 183888 200552 186872 200580
rect 183888 200540 183894 200552
rect 186866 200540 186872 200552
rect 186924 200540 186930 200592
rect 197354 200512 197360 200524
rect 161814 200212 162854 200240
rect 163930 200484 197360 200512
rect 161814 200104 161842 200212
rect 161722 200076 161842 200104
rect 162826 200144 163176 200172
rect 155374 200008 161658 200036
rect 155374 199912 155402 200008
rect 160020 199940 161474 199968
rect 151768 199860 151774 199912
rect 151826 199860 151832 199912
rect 151860 199860 151866 199912
rect 151918 199860 151924 199912
rect 151952 199860 151958 199912
rect 152010 199860 152016 199912
rect 152136 199860 152142 199912
rect 152194 199860 152200 199912
rect 153056 199860 153062 199912
rect 153114 199860 153120 199912
rect 153240 199860 153246 199912
rect 153298 199860 153304 199912
rect 153332 199860 153338 199912
rect 153390 199860 153396 199912
rect 153516 199860 153522 199912
rect 153574 199860 153580 199912
rect 153700 199860 153706 199912
rect 153758 199860 153764 199912
rect 153792 199860 153798 199912
rect 153850 199860 153856 199912
rect 154068 199860 154074 199912
rect 154126 199900 154132 199912
rect 154126 199860 154160 199900
rect 154252 199860 154258 199912
rect 154310 199860 154316 199912
rect 154528 199860 154534 199912
rect 154586 199860 154592 199912
rect 154712 199860 154718 199912
rect 154770 199900 154776 199912
rect 154770 199860 154804 199900
rect 154988 199860 154994 199912
rect 155046 199860 155052 199912
rect 155080 199860 155086 199912
rect 155138 199860 155144 199912
rect 155172 199860 155178 199912
rect 155230 199860 155236 199912
rect 155356 199860 155362 199912
rect 155414 199860 155420 199912
rect 155448 199860 155454 199912
rect 155506 199860 155512 199912
rect 155816 199860 155822 199912
rect 155874 199860 155880 199912
rect 156092 199860 156098 199912
rect 156150 199860 156156 199912
rect 156460 199900 156466 199912
rect 156432 199860 156466 199900
rect 156518 199860 156524 199912
rect 156644 199860 156650 199912
rect 156702 199860 156708 199912
rect 156736 199860 156742 199912
rect 156794 199860 156800 199912
rect 156920 199860 156926 199912
rect 156978 199860 156984 199912
rect 157104 199860 157110 199912
rect 157162 199860 157168 199912
rect 157288 199860 157294 199912
rect 157346 199860 157352 199912
rect 157380 199860 157386 199912
rect 157438 199860 157444 199912
rect 157656 199860 157662 199912
rect 157714 199860 157720 199912
rect 157932 199860 157938 199912
rect 157990 199860 157996 199912
rect 158208 199860 158214 199912
rect 158266 199860 158272 199912
rect 158484 199860 158490 199912
rect 158542 199860 158548 199912
rect 158760 199860 158766 199912
rect 158818 199860 158824 199912
rect 158944 199860 158950 199912
rect 159002 199860 159008 199912
rect 159220 199860 159226 199912
rect 159278 199860 159284 199912
rect 159312 199860 159318 199912
rect 159370 199860 159376 199912
rect 159496 199860 159502 199912
rect 159554 199860 159560 199912
rect 159864 199860 159870 199912
rect 159922 199860 159928 199912
rect 151786 199832 151814 199860
rect 151740 199804 151814 199832
rect 151740 199560 151768 199804
rect 151878 199776 151906 199860
rect 151814 199724 151820 199776
rect 151872 199736 151906 199776
rect 151872 199724 151878 199736
rect 151970 199708 151998 199860
rect 152688 199832 152694 199844
rect 151906 199656 151912 199708
rect 151964 199668 151998 199708
rect 152108 199804 152694 199832
rect 151964 199656 151970 199668
rect 151998 199588 152004 199640
rect 152056 199628 152062 199640
rect 152108 199628 152136 199804
rect 152688 199792 152694 199804
rect 152746 199792 152752 199844
rect 152780 199792 152786 199844
rect 152838 199792 152844 199844
rect 152964 199792 152970 199844
rect 153022 199792 153028 199844
rect 152056 199600 152136 199628
rect 152056 199588 152062 199600
rect 152458 199560 152464 199572
rect 151740 199532 152464 199560
rect 152458 199520 152464 199532
rect 152516 199520 152522 199572
rect 152642 199520 152648 199572
rect 152700 199560 152706 199572
rect 152798 199560 152826 199792
rect 152982 199764 153010 199792
rect 152936 199736 153010 199764
rect 152936 199640 152964 199736
rect 152918 199588 152924 199640
rect 152976 199588 152982 199640
rect 152700 199532 152826 199560
rect 152700 199520 152706 199532
rect 151648 199464 152228 199492
rect 119890 199384 119896 199436
rect 119948 199424 119954 199436
rect 145650 199424 145656 199436
rect 119948 199396 145656 199424
rect 119948 199384 119954 199396
rect 145650 199384 145656 199396
rect 145708 199384 145714 199436
rect 146846 199384 146852 199436
rect 146904 199424 146910 199436
rect 146904 199396 150434 199424
rect 146904 199384 146910 199396
rect 121178 199316 121184 199368
rect 121236 199356 121242 199368
rect 148134 199356 148140 199368
rect 121236 199328 148140 199356
rect 121236 199316 121242 199328
rect 148134 199316 148140 199328
rect 148192 199316 148198 199368
rect 117222 199248 117228 199300
rect 117280 199288 117286 199300
rect 145190 199288 145196 199300
rect 117280 199260 145196 199288
rect 117280 199248 117286 199260
rect 145190 199248 145196 199260
rect 145248 199248 145254 199300
rect 108850 199180 108856 199232
rect 108908 199220 108914 199232
rect 131482 199220 131488 199232
rect 108908 199192 131488 199220
rect 108908 199180 108914 199192
rect 131482 199180 131488 199192
rect 131540 199180 131546 199232
rect 131574 199180 131580 199232
rect 131632 199220 131638 199232
rect 136818 199220 136824 199232
rect 131632 199192 136824 199220
rect 131632 199180 131638 199192
rect 136818 199180 136824 199192
rect 136876 199180 136882 199232
rect 138842 199180 138848 199232
rect 138900 199220 138906 199232
rect 139026 199220 139032 199232
rect 138900 199192 139032 199220
rect 138900 199180 138906 199192
rect 139026 199180 139032 199192
rect 139084 199180 139090 199232
rect 145926 199220 145932 199232
rect 140746 199192 145932 199220
rect 114370 199112 114376 199164
rect 114428 199152 114434 199164
rect 140746 199152 140774 199192
rect 145926 199180 145932 199192
rect 145984 199180 145990 199232
rect 150406 199220 150434 199396
rect 151446 199384 151452 199436
rect 151504 199424 151510 199436
rect 151814 199424 151820 199436
rect 151504 199396 151820 199424
rect 151504 199384 151510 199396
rect 151814 199384 151820 199396
rect 151872 199384 151878 199436
rect 152200 199424 152228 199464
rect 152274 199452 152280 199504
rect 152332 199492 152338 199504
rect 153074 199492 153102 199860
rect 153258 199572 153286 199860
rect 153194 199520 153200 199572
rect 153252 199532 153286 199572
rect 153252 199520 153258 199532
rect 152332 199464 153102 199492
rect 153350 199492 153378 199860
rect 153534 199640 153562 199860
rect 153718 199708 153746 199860
rect 153810 199832 153838 199860
rect 153810 199804 154068 199832
rect 153718 199668 153752 199708
rect 153746 199656 153752 199668
rect 153804 199656 153810 199708
rect 153856 199668 153976 199696
rect 153470 199588 153476 199640
rect 153528 199600 153562 199640
rect 153528 199588 153534 199600
rect 153654 199588 153660 199640
rect 153712 199628 153718 199640
rect 153856 199628 153884 199668
rect 153948 199640 153976 199668
rect 153712 199600 153884 199628
rect 153712 199588 153718 199600
rect 153930 199588 153936 199640
rect 153988 199588 153994 199640
rect 153838 199520 153844 199572
rect 153896 199560 153902 199572
rect 154040 199560 154068 199804
rect 153896 199532 154068 199560
rect 153896 199520 153902 199532
rect 153930 199492 153936 199504
rect 153350 199464 153936 199492
rect 152332 199452 152338 199464
rect 153930 199452 153936 199464
rect 153988 199452 153994 199504
rect 154022 199452 154028 199504
rect 154080 199492 154086 199504
rect 154132 199492 154160 199860
rect 154298 199724 154304 199776
rect 154356 199764 154362 199776
rect 154546 199764 154574 199860
rect 154356 199736 154574 199764
rect 154356 199724 154362 199736
rect 154776 199708 154804 199860
rect 154758 199656 154764 199708
rect 154816 199656 154822 199708
rect 154666 199520 154672 199572
rect 154724 199560 154730 199572
rect 155006 199560 155034 199860
rect 154724 199532 155034 199560
rect 154724 199520 154730 199532
rect 155098 199504 155126 199860
rect 155190 199832 155218 199860
rect 155190 199804 155264 199832
rect 155236 199776 155264 199804
rect 155466 199776 155494 199860
rect 155218 199724 155224 199776
rect 155276 199724 155282 199776
rect 155402 199724 155408 199776
rect 155460 199736 155494 199776
rect 155460 199724 155466 199736
rect 155834 199640 155862 199860
rect 156110 199764 156138 199860
rect 156276 199792 156282 199844
rect 156334 199832 156340 199844
rect 156334 199792 156368 199832
rect 156110 199736 156276 199764
rect 156248 199640 156276 199736
rect 155770 199588 155776 199640
rect 155828 199600 155862 199640
rect 155828 199588 155834 199600
rect 155954 199588 155960 199640
rect 156012 199628 156018 199640
rect 156138 199628 156144 199640
rect 156012 199600 156144 199628
rect 156012 199588 156018 199600
rect 156138 199588 156144 199600
rect 156196 199588 156202 199640
rect 156230 199588 156236 199640
rect 156288 199588 156294 199640
rect 155310 199520 155316 199572
rect 155368 199520 155374 199572
rect 155862 199520 155868 199572
rect 155920 199560 155926 199572
rect 156340 199560 156368 199792
rect 156432 199708 156460 199860
rect 156414 199656 156420 199708
rect 156472 199656 156478 199708
rect 156662 199640 156690 199860
rect 156598 199588 156604 199640
rect 156656 199600 156690 199640
rect 156656 199588 156662 199600
rect 156754 199572 156782 199860
rect 156938 199776 156966 199860
rect 156874 199724 156880 199776
rect 156932 199736 156966 199776
rect 156932 199724 156938 199736
rect 157122 199572 157150 199860
rect 157306 199708 157334 199860
rect 157398 199764 157426 199860
rect 157398 199736 157472 199764
rect 157306 199668 157340 199708
rect 157334 199656 157340 199668
rect 157392 199656 157398 199708
rect 157242 199588 157248 199640
rect 157300 199628 157306 199640
rect 157444 199628 157472 199736
rect 157300 199600 157472 199628
rect 157300 199588 157306 199600
rect 155920 199532 156368 199560
rect 155920 199520 155926 199532
rect 156690 199520 156696 199572
rect 156748 199532 156782 199572
rect 156748 199520 156754 199532
rect 157058 199520 157064 199572
rect 157116 199532 157150 199572
rect 157116 199520 157122 199532
rect 154080 199464 154160 199492
rect 154080 199452 154086 199464
rect 155034 199452 155040 199504
rect 155092 199464 155126 199504
rect 155328 199492 155356 199520
rect 155586 199492 155592 199504
rect 155328 199464 155592 199492
rect 155092 199452 155098 199464
rect 155586 199452 155592 199464
rect 155644 199452 155650 199504
rect 157674 199492 157702 199860
rect 157950 199560 157978 199860
rect 158226 199640 158254 199860
rect 158502 199640 158530 199860
rect 158226 199600 158260 199640
rect 158254 199588 158260 199600
rect 158312 199588 158318 199640
rect 158438 199588 158444 199640
rect 158496 199600 158530 199640
rect 158496 199588 158502 199600
rect 158622 199560 158628 199572
rect 157950 199532 158628 199560
rect 158622 199520 158628 199532
rect 158680 199520 158686 199572
rect 155696 199464 157702 199492
rect 158778 199504 158806 199860
rect 158962 199776 158990 199860
rect 159238 199832 159266 199860
rect 159192 199804 159266 199832
rect 158962 199736 158996 199776
rect 158990 199724 158996 199736
rect 159048 199724 159054 199776
rect 159192 199640 159220 199804
rect 159330 199776 159358 199860
rect 159266 199724 159272 199776
rect 159324 199736 159358 199776
rect 159324 199724 159330 199736
rect 159514 199640 159542 199860
rect 159882 199696 159910 199860
rect 159744 199668 159910 199696
rect 159174 199588 159180 199640
rect 159232 199588 159238 199640
rect 159514 199600 159548 199640
rect 159542 199588 159548 199600
rect 159600 199588 159606 199640
rect 158778 199464 158812 199504
rect 153010 199424 153016 199436
rect 152200 199396 153016 199424
rect 153010 199384 153016 199396
rect 153068 199384 153074 199436
rect 153286 199384 153292 199436
rect 153344 199424 153350 199436
rect 155696 199424 155724 199464
rect 158806 199452 158812 199464
rect 158864 199452 158870 199504
rect 159744 199492 159772 199668
rect 159818 199588 159824 199640
rect 159876 199628 159882 199640
rect 160020 199628 160048 199940
rect 161446 199912 161474 199940
rect 160140 199860 160146 199912
rect 160198 199860 160204 199912
rect 160324 199860 160330 199912
rect 160382 199860 160388 199912
rect 160508 199860 160514 199912
rect 160566 199860 160572 199912
rect 160692 199860 160698 199912
rect 160750 199860 160756 199912
rect 160784 199860 160790 199912
rect 160842 199860 160848 199912
rect 161152 199860 161158 199912
rect 161210 199860 161216 199912
rect 161428 199860 161434 199912
rect 161486 199860 161492 199912
rect 159876 199600 160048 199628
rect 160158 199640 160186 199860
rect 160342 199640 160370 199860
rect 160526 199640 160554 199860
rect 160710 199764 160738 199860
rect 160158 199600 160192 199640
rect 159876 199588 159882 199600
rect 160186 199588 160192 199600
rect 160244 199588 160250 199640
rect 160342 199600 160376 199640
rect 160370 199588 160376 199600
rect 160428 199588 160434 199640
rect 160462 199588 160468 199640
rect 160520 199600 160554 199640
rect 160664 199736 160738 199764
rect 160664 199628 160692 199736
rect 160802 199708 160830 199860
rect 160738 199656 160744 199708
rect 160796 199668 160830 199708
rect 160796 199656 160802 199668
rect 160922 199628 160928 199640
rect 160664 199600 160928 199628
rect 160520 199588 160526 199600
rect 160922 199588 160928 199600
rect 160980 199588 160986 199640
rect 161170 199628 161198 199860
rect 161630 199832 161658 200008
rect 161722 199912 161750 200076
rect 162826 200036 162854 200144
rect 161814 200008 162854 200036
rect 161704 199860 161710 199912
rect 161762 199860 161768 199912
rect 161814 199832 161842 200008
rect 162182 199940 163084 199968
rect 162182 199912 162210 199940
rect 161888 199860 161894 199912
rect 161946 199860 161952 199912
rect 162164 199860 162170 199912
rect 162222 199860 162228 199912
rect 162256 199860 162262 199912
rect 162314 199860 162320 199912
rect 162348 199860 162354 199912
rect 162406 199860 162412 199912
rect 162440 199860 162446 199912
rect 162498 199900 162504 199912
rect 162624 199900 162630 199912
rect 162498 199860 162532 199900
rect 161630 199804 161842 199832
rect 161566 199628 161572 199640
rect 161170 199600 161572 199628
rect 161566 199588 161572 199600
rect 161624 199588 161630 199640
rect 160646 199520 160652 199572
rect 160704 199560 160710 199572
rect 161658 199560 161664 199572
rect 160704 199532 161664 199560
rect 160704 199520 160710 199532
rect 161658 199520 161664 199532
rect 161716 199520 161722 199572
rect 159910 199492 159916 199504
rect 159744 199464 159916 199492
rect 159910 199452 159916 199464
rect 159968 199452 159974 199504
rect 153344 199396 155724 199424
rect 153344 199384 153350 199396
rect 156138 199384 156144 199436
rect 156196 199424 156202 199436
rect 161198 199424 161204 199436
rect 156196 199396 161204 199424
rect 156196 199384 156202 199396
rect 161198 199384 161204 199396
rect 161256 199384 161262 199436
rect 150802 199316 150808 199368
rect 150860 199356 150866 199368
rect 155954 199356 155960 199368
rect 150860 199328 155960 199356
rect 150860 199316 150866 199328
rect 155954 199316 155960 199328
rect 156012 199316 156018 199368
rect 159358 199316 159364 199368
rect 159416 199356 159422 199368
rect 161906 199356 161934 199860
rect 162274 199832 162302 199860
rect 162228 199804 162302 199832
rect 162072 199764 162078 199776
rect 162044 199724 162078 199764
rect 162130 199724 162136 199776
rect 162044 199572 162072 199724
rect 162026 199520 162032 199572
rect 162084 199520 162090 199572
rect 162228 199504 162256 199804
rect 162366 199776 162394 199860
rect 162302 199724 162308 199776
rect 162360 199736 162394 199776
rect 162360 199724 162366 199736
rect 162504 199572 162532 199860
rect 162596 199860 162630 199900
rect 162682 199860 162688 199912
rect 162596 199640 162624 199860
rect 163056 199640 163084 199940
rect 162578 199588 162584 199640
rect 162636 199588 162642 199640
rect 163038 199588 163044 199640
rect 163096 199588 163102 199640
rect 163148 199628 163176 200144
rect 163930 199912 163958 200484
rect 197354 200472 197360 200484
rect 197412 200472 197418 200524
rect 198826 200444 198832 200456
rect 165310 200416 198832 200444
rect 165310 199912 165338 200416
rect 198826 200404 198832 200416
rect 198884 200404 198890 200456
rect 178862 200376 178868 200388
rect 167242 200348 178868 200376
rect 167242 199912 167270 200348
rect 178862 200336 178868 200348
rect 178920 200336 178926 200388
rect 193306 200308 193312 200320
rect 168024 200280 193312 200308
rect 168024 199968 168052 200280
rect 193306 200268 193312 200280
rect 193364 200268 193370 200320
rect 178034 200200 178040 200252
rect 178092 200240 178098 200252
rect 193490 200240 193496 200252
rect 178092 200212 193496 200240
rect 178092 200200 178098 200212
rect 193490 200200 193496 200212
rect 193548 200200 193554 200252
rect 186774 200172 186780 200184
rect 171014 200144 186780 200172
rect 167656 199940 168052 199968
rect 168806 200008 169524 200036
rect 163912 199860 163918 199912
rect 163970 199860 163976 199912
rect 164556 199860 164562 199912
rect 164614 199860 164620 199912
rect 164648 199860 164654 199912
rect 164706 199860 164712 199912
rect 164740 199860 164746 199912
rect 164798 199900 164804 199912
rect 164924 199900 164930 199912
rect 164798 199860 164832 199900
rect 164574 199640 164602 199860
rect 163774 199628 163780 199640
rect 163148 199600 163780 199628
rect 163774 199588 163780 199600
rect 163832 199588 163838 199640
rect 164510 199588 164516 199640
rect 164568 199600 164602 199640
rect 164666 199640 164694 199860
rect 164804 199708 164832 199860
rect 164896 199860 164930 199900
rect 164982 199860 164988 199912
rect 165016 199860 165022 199912
rect 165074 199860 165080 199912
rect 165108 199860 165114 199912
rect 165166 199860 165172 199912
rect 165292 199860 165298 199912
rect 165350 199860 165356 199912
rect 165384 199860 165390 199912
rect 165442 199860 165448 199912
rect 165476 199860 165482 199912
rect 165534 199860 165540 199912
rect 165568 199860 165574 199912
rect 165626 199860 165632 199912
rect 165660 199860 165666 199912
rect 165718 199860 165724 199912
rect 165752 199860 165758 199912
rect 165810 199900 165816 199912
rect 165810 199872 166166 199900
rect 165810 199860 165816 199872
rect 164786 199656 164792 199708
rect 164844 199656 164850 199708
rect 164666 199600 164700 199640
rect 164568 199588 164574 199600
rect 164694 199588 164700 199600
rect 164752 199588 164758 199640
rect 164896 199628 164924 199860
rect 165034 199832 165062 199860
rect 164988 199804 165062 199832
rect 164988 199708 165016 199804
rect 165126 199708 165154 199860
rect 165402 199832 165430 199860
rect 165356 199804 165430 199832
rect 165356 199708 165384 199804
rect 165494 199776 165522 199860
rect 165430 199724 165436 199776
rect 165488 199736 165522 199776
rect 165488 199724 165494 199736
rect 165586 199708 165614 199860
rect 165678 199764 165706 199860
rect 166028 199792 166034 199844
rect 166086 199792 166092 199844
rect 165678 199736 165752 199764
rect 165724 199708 165752 199736
rect 164970 199656 164976 199708
rect 165028 199656 165034 199708
rect 165062 199656 165068 199708
rect 165120 199668 165154 199708
rect 165120 199656 165126 199668
rect 165338 199656 165344 199708
rect 165396 199656 165402 199708
rect 165522 199656 165528 199708
rect 165580 199668 165614 199708
rect 165580 199656 165586 199668
rect 165706 199656 165712 199708
rect 165764 199656 165770 199708
rect 166046 199640 166074 199792
rect 165154 199628 165160 199640
rect 164896 199600 165160 199628
rect 165154 199588 165160 199600
rect 165212 199588 165218 199640
rect 165982 199588 165988 199640
rect 166040 199600 166074 199640
rect 166040 199588 166046 199600
rect 162486 199520 162492 199572
rect 162544 199520 162550 199572
rect 166138 199560 166166 199872
rect 166212 199860 166218 199912
rect 166270 199860 166276 199912
rect 166764 199900 166770 199912
rect 166736 199860 166770 199900
rect 166822 199860 166828 199912
rect 166856 199860 166862 199912
rect 166914 199860 166920 199912
rect 167040 199860 167046 199912
rect 167098 199860 167104 199912
rect 167132 199860 167138 199912
rect 167190 199860 167196 199912
rect 167224 199860 167230 199912
rect 167282 199860 167288 199912
rect 167408 199860 167414 199912
rect 167466 199860 167472 199912
rect 166230 199628 166258 199860
rect 166304 199792 166310 199844
rect 166362 199792 166368 199844
rect 166322 199696 166350 199792
rect 166736 199776 166764 199860
rect 166874 199776 166902 199860
rect 166718 199724 166724 199776
rect 166776 199724 166782 199776
rect 166874 199736 166908 199776
rect 166902 199724 166908 199736
rect 166960 199724 166966 199776
rect 166810 199696 166816 199708
rect 166322 199668 166816 199696
rect 166810 199656 166816 199668
rect 166868 199656 166874 199708
rect 166230 199600 166948 199628
rect 166810 199560 166816 199572
rect 166138 199532 166816 199560
rect 166810 199520 166816 199532
rect 166868 199520 166874 199572
rect 162210 199452 162216 199504
rect 162268 199452 162274 199504
rect 162762 199452 162768 199504
rect 162820 199492 162826 199504
rect 164234 199492 164240 199504
rect 162820 199464 164240 199492
rect 162820 199452 162826 199464
rect 164234 199452 164240 199464
rect 164292 199452 164298 199504
rect 166166 199452 166172 199504
rect 166224 199492 166230 199504
rect 166920 199492 166948 199600
rect 167058 199572 167086 199860
rect 167150 199708 167178 199860
rect 167150 199668 167184 199708
rect 167178 199656 167184 199668
rect 167236 199656 167242 199708
rect 167426 199640 167454 199860
rect 167362 199588 167368 199640
rect 167420 199600 167454 199640
rect 167420 199588 167426 199600
rect 166994 199520 167000 199572
rect 167052 199532 167086 199572
rect 167052 199520 167058 199532
rect 166224 199464 166948 199492
rect 166224 199452 166230 199464
rect 165246 199384 165252 199436
rect 165304 199424 165310 199436
rect 165614 199424 165620 199436
rect 165304 199396 165620 199424
rect 165304 199384 165310 199396
rect 165614 199384 165620 199396
rect 165672 199384 165678 199436
rect 159416 199328 161934 199356
rect 159416 199316 159422 199328
rect 162762 199316 162768 199368
rect 162820 199356 162826 199368
rect 167656 199356 167684 199940
rect 168806 199912 168834 200008
rect 168990 199940 169386 199968
rect 168990 199912 169018 199940
rect 167868 199860 167874 199912
rect 167926 199860 167932 199912
rect 167960 199860 167966 199912
rect 168018 199860 168024 199912
rect 168052 199860 168058 199912
rect 168110 199860 168116 199912
rect 168420 199860 168426 199912
rect 168478 199860 168484 199912
rect 168788 199860 168794 199912
rect 168846 199860 168852 199912
rect 168880 199860 168886 199912
rect 168938 199860 168944 199912
rect 168972 199860 168978 199912
rect 169030 199860 169036 199912
rect 169248 199860 169254 199912
rect 169306 199860 169312 199912
rect 167886 199832 167914 199860
rect 167840 199804 167914 199832
rect 167840 199492 167868 199804
rect 167978 199776 168006 199860
rect 167914 199724 167920 199776
rect 167972 199736 168006 199776
rect 167972 199724 167978 199736
rect 168070 199708 168098 199860
rect 168006 199656 168012 199708
rect 168064 199668 168098 199708
rect 168064 199656 168070 199668
rect 168438 199640 168466 199860
rect 168898 199832 168926 199860
rect 168760 199804 168926 199832
rect 168438 199600 168472 199640
rect 168466 199588 168472 199600
rect 168524 199588 168530 199640
rect 168760 199628 168788 199804
rect 169266 199764 169294 199860
rect 168852 199736 169294 199764
rect 168852 199708 168880 199736
rect 168834 199656 168840 199708
rect 168892 199656 168898 199708
rect 168926 199656 168932 199708
rect 168984 199696 168990 199708
rect 169358 199696 169386 199940
rect 168984 199668 169386 199696
rect 168984 199656 168990 199668
rect 169386 199628 169392 199640
rect 168760 199600 169392 199628
rect 169386 199588 169392 199600
rect 169444 199588 169450 199640
rect 169202 199520 169208 199572
rect 169260 199560 169266 199572
rect 169496 199560 169524 200008
rect 169616 199900 169622 199912
rect 169588 199860 169622 199900
rect 169674 199860 169680 199912
rect 169708 199860 169714 199912
rect 169766 199860 169772 199912
rect 169800 199860 169806 199912
rect 169858 199860 169864 199912
rect 169892 199860 169898 199912
rect 169950 199860 169956 199912
rect 170076 199860 170082 199912
rect 170134 199860 170140 199912
rect 170168 199860 170174 199912
rect 170226 199860 170232 199912
rect 170536 199860 170542 199912
rect 170594 199860 170600 199912
rect 170628 199860 170634 199912
rect 170686 199860 170692 199912
rect 170720 199860 170726 199912
rect 170778 199860 170784 199912
rect 170812 199860 170818 199912
rect 170870 199900 170876 199912
rect 170870 199860 170904 199900
rect 169588 199708 169616 199860
rect 169726 199832 169754 199860
rect 169680 199804 169754 199832
rect 169680 199708 169708 199804
rect 169818 199764 169846 199860
rect 169772 199736 169846 199764
rect 169570 199656 169576 199708
rect 169628 199656 169634 199708
rect 169662 199656 169668 199708
rect 169720 199656 169726 199708
rect 169260 199532 169524 199560
rect 169260 199520 169266 199532
rect 169570 199520 169576 199572
rect 169628 199520 169634 199572
rect 168650 199492 168656 199504
rect 167840 199464 168656 199492
rect 168650 199452 168656 199464
rect 168708 199452 168714 199504
rect 162820 199328 167684 199356
rect 162820 199316 162826 199328
rect 167730 199316 167736 199368
rect 167788 199356 167794 199368
rect 169588 199356 169616 199520
rect 169772 199504 169800 199736
rect 169910 199708 169938 199860
rect 170094 199776 170122 199860
rect 170030 199724 170036 199776
rect 170088 199736 170122 199776
rect 170088 199724 170094 199736
rect 169846 199656 169852 199708
rect 169904 199668 169938 199708
rect 169904 199656 169910 199668
rect 170186 199640 170214 199860
rect 170554 199776 170582 199860
rect 170490 199724 170496 199776
rect 170548 199736 170582 199776
rect 170548 199724 170554 199736
rect 170646 199708 170674 199860
rect 170582 199656 170588 199708
rect 170640 199668 170674 199708
rect 170738 199696 170766 199860
rect 170738 199668 170812 199696
rect 170640 199656 170646 199668
rect 170122 199588 170128 199640
rect 170180 199600 170214 199640
rect 170180 199588 170186 199600
rect 170784 199504 170812 199668
rect 170876 199572 170904 199860
rect 171014 199776 171042 200144
rect 186774 200132 186780 200144
rect 186832 200132 186838 200184
rect 186866 200132 186872 200184
rect 186924 200172 186930 200184
rect 190546 200172 190552 200184
rect 186924 200144 190552 200172
rect 186924 200132 186930 200144
rect 190546 200132 190552 200144
rect 190604 200132 190610 200184
rect 181898 200104 181904 200116
rect 171934 200076 181904 200104
rect 171934 199912 171962 200076
rect 181898 200064 181904 200076
rect 181956 200064 181962 200116
rect 187510 200036 187516 200048
rect 172210 200008 175366 200036
rect 172210 199912 172238 200008
rect 172762 199940 173388 199968
rect 172762 199912 172790 199940
rect 171088 199860 171094 199912
rect 171146 199900 171152 199912
rect 171146 199872 171226 199900
rect 171146 199860 171152 199872
rect 171014 199736 171048 199776
rect 171042 199724 171048 199736
rect 171100 199724 171106 199776
rect 170858 199520 170864 199572
rect 170916 199520 170922 199572
rect 171198 199560 171226 199872
rect 171272 199860 171278 199912
rect 171330 199860 171336 199912
rect 171824 199860 171830 199912
rect 171882 199860 171888 199912
rect 171916 199860 171922 199912
rect 171974 199860 171980 199912
rect 172192 199860 172198 199912
rect 172250 199860 172256 199912
rect 172560 199860 172566 199912
rect 172618 199860 172624 199912
rect 172744 199860 172750 199912
rect 172802 199860 172808 199912
rect 173112 199860 173118 199912
rect 173170 199860 173176 199912
rect 171290 199696 171318 199860
rect 171842 199708 171870 199860
rect 171290 199668 171364 199696
rect 171842 199668 171876 199708
rect 171336 199640 171364 199668
rect 171870 199656 171876 199668
rect 171928 199656 171934 199708
rect 171318 199588 171324 199640
rect 171376 199588 171382 199640
rect 172054 199588 172060 199640
rect 172112 199628 172118 199640
rect 172238 199628 172244 199640
rect 172112 199600 172244 199628
rect 172112 199588 172118 199600
rect 172238 199588 172244 199600
rect 172296 199588 172302 199640
rect 172578 199628 172606 199860
rect 173130 199696 173158 199860
rect 172348 199600 172606 199628
rect 172670 199668 173158 199696
rect 172348 199572 172376 199600
rect 172146 199560 172152 199572
rect 171198 199532 172152 199560
rect 172146 199520 172152 199532
rect 172204 199520 172210 199572
rect 172330 199520 172336 199572
rect 172388 199520 172394 199572
rect 172422 199520 172428 199572
rect 172480 199560 172486 199572
rect 172670 199560 172698 199668
rect 172480 199532 172698 199560
rect 172480 199520 172486 199532
rect 172790 199520 172796 199572
rect 172848 199520 172854 199572
rect 169754 199452 169760 199504
rect 169812 199452 169818 199504
rect 170766 199452 170772 199504
rect 170824 199452 170830 199504
rect 171594 199452 171600 199504
rect 171652 199492 171658 199504
rect 171962 199492 171968 199504
rect 171652 199464 171968 199492
rect 171652 199452 171658 199464
rect 171962 199452 171968 199464
rect 172020 199452 172026 199504
rect 169754 199356 169760 199368
rect 167788 199328 169064 199356
rect 169588 199328 169760 199356
rect 167788 199316 167794 199328
rect 151078 199248 151084 199300
rect 151136 199288 151142 199300
rect 157150 199288 157156 199300
rect 151136 199260 157156 199288
rect 151136 199248 151142 199260
rect 157150 199248 157156 199260
rect 157208 199248 157214 199300
rect 160554 199248 160560 199300
rect 160612 199288 160618 199300
rect 161842 199288 161848 199300
rect 160612 199260 161848 199288
rect 160612 199248 160618 199260
rect 161842 199248 161848 199260
rect 161900 199248 161906 199300
rect 164878 199248 164884 199300
rect 164936 199288 164942 199300
rect 169036 199288 169064 199328
rect 169754 199316 169760 199328
rect 169812 199316 169818 199368
rect 171962 199316 171968 199368
rect 172020 199356 172026 199368
rect 172808 199356 172836 199520
rect 173360 199504 173388 199940
rect 173590 199940 173894 199968
rect 173590 199912 173618 199940
rect 173572 199860 173578 199912
rect 173630 199860 173636 199912
rect 173526 199520 173532 199572
rect 173584 199560 173590 199572
rect 173866 199560 173894 199940
rect 174602 199940 174814 199968
rect 174032 199860 174038 199912
rect 174090 199860 174096 199912
rect 174124 199860 174130 199912
rect 174182 199860 174188 199912
rect 174216 199860 174222 199912
rect 174274 199900 174280 199912
rect 174274 199860 174308 199900
rect 174400 199860 174406 199912
rect 174458 199860 174464 199912
rect 174492 199860 174498 199912
rect 174550 199860 174556 199912
rect 174050 199776 174078 199860
rect 174142 199832 174170 199860
rect 174142 199804 174216 199832
rect 174050 199736 174084 199776
rect 174078 199724 174084 199736
rect 174136 199724 174142 199776
rect 173584 199532 173894 199560
rect 173584 199520 173590 199532
rect 174188 199504 174216 199804
rect 174280 199572 174308 199860
rect 174418 199764 174446 199860
rect 174372 199736 174446 199764
rect 174262 199520 174268 199572
rect 174320 199520 174326 199572
rect 173342 199452 173348 199504
rect 173400 199452 173406 199504
rect 174170 199452 174176 199504
rect 174228 199452 174234 199504
rect 174372 199492 174400 199736
rect 174510 199708 174538 199860
rect 174446 199656 174452 199708
rect 174504 199668 174538 199708
rect 174504 199656 174510 199668
rect 174602 199560 174630 199940
rect 174786 199912 174814 199940
rect 174676 199860 174682 199912
rect 174734 199860 174740 199912
rect 174768 199860 174774 199912
rect 174826 199860 174832 199912
rect 174952 199860 174958 199912
rect 175010 199860 175016 199912
rect 174694 199628 174722 199860
rect 174970 199640 174998 199860
rect 174814 199628 174820 199640
rect 174694 199600 174820 199628
rect 174814 199588 174820 199600
rect 174872 199588 174878 199640
rect 174970 199600 175004 199640
rect 174998 199588 175004 199600
rect 175056 199588 175062 199640
rect 174722 199560 174728 199572
rect 174602 199532 174728 199560
rect 174722 199520 174728 199532
rect 174780 199520 174786 199572
rect 175338 199560 175366 200008
rect 176074 200008 187516 200036
rect 176074 199912 176102 200008
rect 187510 199996 187516 200008
rect 187568 199996 187574 200048
rect 176718 199940 198734 199968
rect 176718 199912 176746 199940
rect 175504 199860 175510 199912
rect 175562 199860 175568 199912
rect 175596 199860 175602 199912
rect 175654 199860 175660 199912
rect 175964 199860 175970 199912
rect 176022 199860 176028 199912
rect 176056 199860 176062 199912
rect 176114 199860 176120 199912
rect 176148 199860 176154 199912
rect 176206 199860 176212 199912
rect 176240 199860 176246 199912
rect 176298 199860 176304 199912
rect 176700 199860 176706 199912
rect 176758 199860 176764 199912
rect 176792 199860 176798 199912
rect 176850 199860 176856 199912
rect 176976 199860 176982 199912
rect 177034 199860 177040 199912
rect 177252 199860 177258 199912
rect 177310 199900 177316 199912
rect 177666 199900 177672 199912
rect 177310 199872 177672 199900
rect 177310 199860 177316 199872
rect 177666 199860 177672 199872
rect 177724 199860 177730 199912
rect 175522 199764 175550 199860
rect 175476 199736 175550 199764
rect 175476 199628 175504 199736
rect 175614 199708 175642 199860
rect 175982 199776 176010 199860
rect 176166 199776 176194 199860
rect 175918 199724 175924 199776
rect 175976 199736 176010 199776
rect 175976 199724 175982 199736
rect 176102 199724 176108 199776
rect 176160 199736 176194 199776
rect 176160 199724 176166 199736
rect 175550 199656 175556 199708
rect 175608 199668 175642 199708
rect 175608 199656 175614 199668
rect 176258 199640 176286 199860
rect 176810 199776 176838 199860
rect 176994 199776 177022 199860
rect 195514 199832 195520 199844
rect 177178 199804 195520 199832
rect 177178 199776 177206 199804
rect 195514 199792 195520 199804
rect 195572 199792 195578 199844
rect 176810 199736 176844 199776
rect 176838 199724 176844 199736
rect 176896 199724 176902 199776
rect 176930 199724 176936 199776
rect 176988 199736 177022 199776
rect 176988 199724 176994 199736
rect 177160 199724 177166 199776
rect 177218 199724 177224 199776
rect 198706 199764 198734 199940
rect 199562 199764 199568 199776
rect 198706 199736 199568 199764
rect 199562 199724 199568 199736
rect 199620 199724 199626 199776
rect 176010 199628 176016 199640
rect 175476 199600 176016 199628
rect 176010 199588 176016 199600
rect 176068 199588 176074 199640
rect 176194 199588 176200 199640
rect 176252 199600 176286 199640
rect 176252 199588 176258 199600
rect 177390 199560 177396 199572
rect 175338 199532 177396 199560
rect 177390 199520 177396 199532
rect 177448 199520 177454 199572
rect 177666 199520 177672 199572
rect 177724 199560 177730 199572
rect 177942 199560 177948 199572
rect 177724 199532 177948 199560
rect 177724 199520 177730 199532
rect 177942 199520 177948 199532
rect 178000 199520 178006 199572
rect 178218 199520 178224 199572
rect 178276 199560 178282 199572
rect 186590 199560 186596 199572
rect 178276 199532 186596 199560
rect 178276 199520 178282 199532
rect 186590 199520 186596 199532
rect 186648 199520 186654 199572
rect 175182 199492 175188 199504
rect 174372 199464 175188 199492
rect 175182 199452 175188 199464
rect 175240 199452 175246 199504
rect 175918 199452 175924 199504
rect 175976 199492 175982 199504
rect 176378 199492 176384 199504
rect 175976 199464 176384 199492
rect 175976 199452 175982 199464
rect 176378 199452 176384 199464
rect 176436 199452 176442 199504
rect 177574 199452 177580 199504
rect 177632 199492 177638 199504
rect 178126 199492 178132 199504
rect 177632 199464 178132 199492
rect 177632 199452 177638 199464
rect 178126 199452 178132 199464
rect 178184 199452 178190 199504
rect 173802 199384 173808 199436
rect 173860 199424 173866 199436
rect 180334 199424 180340 199436
rect 173860 199396 180340 199424
rect 173860 199384 173866 199396
rect 180334 199384 180340 199396
rect 180392 199384 180398 199436
rect 182818 199384 182824 199436
rect 182876 199424 182882 199436
rect 190454 199424 190460 199436
rect 182876 199396 190460 199424
rect 182876 199384 182882 199396
rect 190454 199384 190460 199396
rect 190512 199384 190518 199436
rect 203058 199356 203064 199368
rect 172020 199328 172836 199356
rect 191806 199328 203064 199356
rect 172020 199316 172026 199328
rect 178034 199288 178040 199300
rect 164936 199260 168972 199288
rect 169036 199260 178040 199288
rect 164936 199248 164942 199260
rect 156138 199220 156144 199232
rect 150406 199192 156144 199220
rect 156138 199180 156144 199192
rect 156196 199180 156202 199232
rect 159726 199180 159732 199232
rect 159784 199220 159790 199232
rect 159784 199192 167500 199220
rect 159784 199180 159790 199192
rect 114428 199124 140774 199152
rect 114428 199112 114434 199124
rect 143626 199112 143632 199164
rect 143684 199152 143690 199164
rect 148410 199152 148416 199164
rect 143684 199124 148416 199152
rect 143684 199112 143690 199124
rect 148410 199112 148416 199124
rect 148468 199112 148474 199164
rect 152826 199112 152832 199164
rect 152884 199152 152890 199164
rect 152884 199124 160140 199152
rect 152884 199112 152890 199124
rect 115750 199044 115756 199096
rect 115808 199084 115814 199096
rect 147582 199084 147588 199096
rect 115808 199056 147588 199084
rect 115808 199044 115814 199056
rect 147582 199044 147588 199056
rect 147640 199044 147646 199096
rect 159450 199044 159456 199096
rect 159508 199084 159514 199096
rect 160002 199084 160008 199096
rect 159508 199056 160008 199084
rect 159508 199044 159514 199056
rect 160002 199044 160008 199056
rect 160060 199044 160066 199096
rect 160112 199084 160140 199124
rect 162394 199112 162400 199164
rect 162452 199152 162458 199164
rect 165706 199152 165712 199164
rect 162452 199124 165712 199152
rect 162452 199112 162458 199124
rect 165706 199112 165712 199124
rect 165764 199112 165770 199164
rect 164878 199084 164884 199096
rect 160112 199056 164884 199084
rect 164878 199044 164884 199056
rect 164936 199044 164942 199096
rect 167472 199084 167500 199192
rect 168944 199152 168972 199260
rect 178034 199248 178040 199260
rect 178092 199248 178098 199300
rect 169386 199180 169392 199232
rect 169444 199220 169450 199232
rect 169444 199192 172284 199220
rect 169444 199180 169450 199192
rect 171134 199152 171140 199164
rect 168944 199124 171140 199152
rect 171134 199112 171140 199124
rect 171192 199112 171198 199164
rect 172256 199152 172284 199192
rect 172330 199180 172336 199232
rect 172388 199220 172394 199232
rect 173710 199220 173716 199232
rect 172388 199192 173716 199220
rect 172388 199180 172394 199192
rect 173710 199180 173716 199192
rect 173768 199180 173774 199232
rect 191806 199220 191834 199328
rect 203058 199316 203064 199328
rect 203116 199316 203122 199368
rect 175108 199192 191834 199220
rect 175108 199152 175136 199192
rect 172256 199124 175136 199152
rect 175182 199112 175188 199164
rect 175240 199152 175246 199164
rect 201034 199152 201040 199164
rect 175240 199124 201040 199152
rect 175240 199112 175246 199124
rect 201034 199112 201040 199124
rect 201092 199112 201098 199164
rect 169386 199084 169392 199096
rect 167472 199056 169392 199084
rect 169386 199044 169392 199056
rect 169444 199044 169450 199096
rect 169938 199044 169944 199096
rect 169996 199084 170002 199096
rect 170766 199084 170772 199096
rect 169996 199056 170772 199084
rect 169996 199044 170002 199056
rect 170766 199044 170772 199056
rect 170824 199044 170830 199096
rect 175734 199044 175740 199096
rect 175792 199084 175798 199096
rect 186406 199084 186412 199096
rect 175792 199056 186412 199084
rect 175792 199044 175798 199056
rect 186406 199044 186412 199056
rect 186464 199044 186470 199096
rect 187510 199044 187516 199096
rect 187568 199084 187574 199096
rect 198734 199084 198740 199096
rect 187568 199056 198740 199084
rect 187568 199044 187574 199056
rect 198734 199044 198740 199056
rect 198792 199044 198798 199096
rect 133138 198976 133144 199028
rect 133196 199016 133202 199028
rect 159818 199016 159824 199028
rect 133196 198988 159824 199016
rect 133196 198976 133202 198988
rect 159818 198976 159824 198988
rect 159876 198976 159882 199028
rect 166350 198976 166356 199028
rect 166408 199016 166414 199028
rect 200206 199016 200212 199028
rect 166408 198988 200212 199016
rect 166408 198976 166414 198988
rect 200206 198976 200212 198988
rect 200264 198976 200270 199028
rect 114462 198908 114468 198960
rect 114520 198948 114526 198960
rect 147030 198948 147036 198960
rect 114520 198920 147036 198948
rect 114520 198908 114526 198920
rect 147030 198908 147036 198920
rect 147088 198908 147094 198960
rect 159634 198908 159640 198960
rect 159692 198948 159698 198960
rect 160002 198948 160008 198960
rect 159692 198920 160008 198948
rect 159692 198908 159698 198920
rect 160002 198908 160008 198920
rect 160060 198908 160066 198960
rect 169386 198908 169392 198960
rect 169444 198948 169450 198960
rect 170766 198948 170772 198960
rect 169444 198920 170772 198948
rect 169444 198908 169450 198920
rect 170766 198908 170772 198920
rect 170824 198908 170830 198960
rect 174262 198908 174268 198960
rect 174320 198948 174326 198960
rect 178770 198948 178776 198960
rect 174320 198920 178776 198948
rect 174320 198908 174326 198920
rect 178770 198908 178776 198920
rect 178828 198908 178834 198960
rect 181070 198908 181076 198960
rect 181128 198948 181134 198960
rect 187694 198948 187700 198960
rect 181128 198920 187700 198948
rect 181128 198908 181134 198920
rect 187694 198908 187700 198920
rect 187752 198908 187758 198960
rect 121362 198840 121368 198892
rect 121420 198880 121426 198892
rect 140314 198880 140320 198892
rect 121420 198852 140320 198880
rect 121420 198840 121426 198852
rect 140314 198840 140320 198852
rect 140372 198840 140378 198892
rect 159174 198840 159180 198892
rect 159232 198880 159238 198892
rect 162762 198880 162768 198892
rect 159232 198852 162768 198880
rect 159232 198840 159238 198852
rect 162762 198840 162768 198852
rect 162820 198840 162826 198892
rect 167454 198840 167460 198892
rect 167512 198880 167518 198892
rect 201862 198880 201868 198892
rect 167512 198852 201868 198880
rect 167512 198840 167518 198852
rect 201862 198840 201868 198852
rect 201920 198840 201926 198892
rect 126330 198772 126336 198824
rect 126388 198812 126394 198824
rect 147674 198812 147680 198824
rect 126388 198784 147680 198812
rect 126388 198772 126394 198784
rect 147674 198772 147680 198784
rect 147732 198772 147738 198824
rect 150250 198772 150256 198824
rect 150308 198812 150314 198824
rect 157426 198812 157432 198824
rect 150308 198784 157432 198812
rect 150308 198772 150314 198784
rect 157426 198772 157432 198784
rect 157484 198772 157490 198824
rect 158990 198772 158996 198824
rect 159048 198812 159054 198824
rect 167730 198812 167736 198824
rect 159048 198784 167736 198812
rect 159048 198772 159054 198784
rect 167730 198772 167736 198784
rect 167788 198772 167794 198824
rect 167822 198772 167828 198824
rect 167880 198812 167886 198824
rect 170122 198812 170128 198824
rect 167880 198784 170128 198812
rect 167880 198772 167886 198784
rect 170122 198772 170128 198784
rect 170180 198772 170186 198824
rect 171134 198772 171140 198824
rect 171192 198812 171198 198824
rect 174262 198812 174268 198824
rect 171192 198784 174268 198812
rect 171192 198772 171198 198784
rect 174262 198772 174268 198784
rect 174320 198772 174326 198824
rect 180150 198812 180156 198824
rect 174372 198784 180156 198812
rect 118602 198704 118608 198756
rect 118660 198744 118666 198756
rect 144362 198744 144368 198756
rect 118660 198716 144368 198744
rect 118660 198704 118666 198716
rect 144362 198704 144368 198716
rect 144420 198704 144426 198756
rect 170766 198704 170772 198756
rect 170824 198744 170830 198756
rect 174372 198744 174400 198784
rect 180150 198772 180156 198784
rect 180208 198772 180214 198824
rect 186406 198772 186412 198824
rect 186464 198812 186470 198824
rect 200942 198812 200948 198824
rect 186464 198784 200948 198812
rect 186464 198772 186470 198784
rect 200942 198772 200948 198784
rect 201000 198772 201006 198824
rect 170824 198716 174400 198744
rect 170824 198704 170830 198716
rect 174814 198704 174820 198756
rect 174872 198744 174878 198756
rect 200574 198744 200580 198756
rect 174872 198716 200580 198744
rect 174872 198704 174878 198716
rect 200574 198704 200580 198716
rect 200632 198704 200638 198756
rect 130930 198636 130936 198688
rect 130988 198676 130994 198688
rect 144822 198676 144828 198688
rect 130988 198648 144828 198676
rect 130988 198636 130994 198648
rect 144822 198636 144828 198648
rect 144880 198636 144886 198688
rect 173066 198636 173072 198688
rect 173124 198676 173130 198688
rect 195974 198676 195980 198688
rect 173124 198648 195980 198676
rect 173124 198636 173130 198648
rect 195974 198636 195980 198648
rect 196032 198636 196038 198688
rect 126698 198568 126704 198620
rect 126756 198608 126762 198620
rect 146662 198608 146668 198620
rect 126756 198580 146668 198608
rect 126756 198568 126762 198580
rect 146662 198568 146668 198580
rect 146720 198568 146726 198620
rect 167086 198568 167092 198620
rect 167144 198608 167150 198620
rect 178678 198608 178684 198620
rect 167144 198580 178684 198608
rect 167144 198568 167150 198580
rect 178678 198568 178684 198580
rect 178736 198568 178742 198620
rect 181898 198568 181904 198620
rect 181956 198608 181962 198620
rect 194042 198608 194048 198620
rect 181956 198580 194048 198608
rect 181956 198568 181962 198580
rect 194042 198568 194048 198580
rect 194100 198568 194106 198620
rect 108666 198500 108672 198552
rect 108724 198540 108730 198552
rect 133322 198540 133328 198552
rect 108724 198512 133328 198540
rect 108724 198500 108730 198512
rect 133322 198500 133328 198512
rect 133380 198500 133386 198552
rect 157886 198500 157892 198552
rect 157944 198540 157950 198552
rect 171778 198540 171784 198552
rect 157944 198512 171784 198540
rect 157944 198500 157950 198512
rect 171778 198500 171784 198512
rect 171836 198500 171842 198552
rect 123294 198432 123300 198484
rect 123352 198472 123358 198484
rect 143718 198472 143724 198484
rect 123352 198444 143724 198472
rect 123352 198432 123358 198444
rect 143718 198432 143724 198444
rect 143776 198432 143782 198484
rect 156690 198432 156696 198484
rect 156748 198472 156754 198484
rect 171502 198472 171508 198484
rect 156748 198444 171508 198472
rect 156748 198432 156754 198444
rect 171502 198432 171508 198444
rect 171560 198432 171566 198484
rect 173250 198432 173256 198484
rect 173308 198472 173314 198484
rect 199102 198472 199108 198484
rect 173308 198444 199108 198472
rect 173308 198432 173314 198444
rect 199102 198432 199108 198444
rect 199160 198432 199166 198484
rect 108390 198364 108396 198416
rect 108448 198404 108454 198416
rect 132494 198404 132500 198416
rect 108448 198376 132500 198404
rect 108448 198364 108454 198376
rect 132494 198364 132500 198376
rect 132552 198364 132558 198416
rect 159818 198364 159824 198416
rect 159876 198404 159882 198416
rect 171318 198404 171324 198416
rect 159876 198376 171324 198404
rect 159876 198364 159882 198376
rect 171318 198364 171324 198376
rect 171376 198364 171382 198416
rect 177390 198364 177396 198416
rect 177448 198404 177454 198416
rect 197722 198404 197728 198416
rect 177448 198376 197728 198404
rect 177448 198364 177454 198376
rect 197722 198364 197728 198376
rect 197780 198364 197786 198416
rect 122466 198296 122472 198348
rect 122524 198336 122530 198348
rect 148226 198336 148232 198348
rect 122524 198308 148232 198336
rect 122524 198296 122530 198308
rect 148226 198296 148232 198308
rect 148284 198296 148290 198348
rect 169938 198296 169944 198348
rect 169996 198336 170002 198348
rect 196618 198336 196624 198348
rect 169996 198308 196624 198336
rect 169996 198296 170002 198308
rect 196618 198296 196624 198308
rect 196676 198296 196682 198348
rect 106918 198228 106924 198280
rect 106976 198268 106982 198280
rect 127526 198268 127532 198280
rect 106976 198240 127532 198268
rect 106976 198228 106982 198240
rect 127526 198228 127532 198240
rect 127584 198228 127590 198280
rect 136542 198228 136548 198280
rect 136600 198268 136606 198280
rect 138014 198268 138020 198280
rect 136600 198240 138020 198268
rect 136600 198228 136606 198240
rect 138014 198228 138020 198240
rect 138072 198228 138078 198280
rect 172514 198228 172520 198280
rect 172572 198268 172578 198280
rect 198182 198268 198188 198280
rect 172572 198240 198188 198268
rect 172572 198228 172578 198240
rect 198182 198228 198188 198240
rect 198240 198228 198246 198280
rect 122282 198160 122288 198212
rect 122340 198200 122346 198212
rect 149146 198200 149152 198212
rect 122340 198172 149152 198200
rect 122340 198160 122346 198172
rect 149146 198160 149152 198172
rect 149204 198160 149210 198212
rect 156414 198160 156420 198212
rect 156472 198200 156478 198212
rect 171318 198200 171324 198212
rect 156472 198172 171324 198200
rect 156472 198160 156478 198172
rect 171318 198160 171324 198172
rect 171376 198160 171382 198212
rect 172146 198160 172152 198212
rect 172204 198200 172210 198212
rect 181438 198200 181444 198212
rect 172204 198172 181444 198200
rect 172204 198160 172210 198172
rect 181438 198160 181444 198172
rect 181496 198160 181502 198212
rect 199562 198160 199568 198212
rect 199620 198200 199626 198212
rect 204714 198200 204720 198212
rect 199620 198172 204720 198200
rect 199620 198160 199626 198172
rect 204714 198160 204720 198172
rect 204772 198160 204778 198212
rect 103330 198092 103336 198144
rect 103388 198132 103394 198144
rect 134886 198132 134892 198144
rect 103388 198104 134892 198132
rect 103388 198092 103394 198104
rect 134886 198092 134892 198104
rect 134944 198092 134950 198144
rect 153378 198092 153384 198144
rect 153436 198132 153442 198144
rect 171134 198132 171140 198144
rect 153436 198104 171140 198132
rect 153436 198092 153442 198104
rect 171134 198092 171140 198104
rect 171192 198092 171198 198144
rect 173894 198092 173900 198144
rect 173952 198132 173958 198144
rect 200390 198132 200396 198144
rect 173952 198104 200396 198132
rect 173952 198092 173958 198104
rect 200390 198092 200396 198104
rect 200448 198092 200454 198144
rect 103422 198024 103428 198076
rect 103480 198064 103486 198076
rect 133598 198064 133604 198076
rect 103480 198036 133604 198064
rect 103480 198024 103486 198036
rect 133598 198024 133604 198036
rect 133656 198024 133662 198076
rect 173342 198024 173348 198076
rect 173400 198064 173406 198076
rect 200666 198064 200672 198076
rect 173400 198036 200672 198064
rect 173400 198024 173406 198036
rect 200666 198024 200672 198036
rect 200724 198024 200730 198076
rect 102870 197956 102876 198008
rect 102928 197996 102934 198008
rect 125594 197996 125600 198008
rect 102928 197968 125600 197996
rect 102928 197956 102934 197968
rect 125594 197956 125600 197968
rect 125652 197956 125658 198008
rect 157610 197956 157616 198008
rect 157668 197996 157674 198008
rect 169754 197996 169760 198008
rect 157668 197968 169760 197996
rect 157668 197956 157674 197968
rect 169754 197956 169760 197968
rect 169812 197956 169818 198008
rect 172238 197956 172244 198008
rect 172296 197996 172302 198008
rect 199378 197996 199384 198008
rect 172296 197968 199384 197996
rect 172296 197956 172302 197968
rect 199378 197956 199384 197968
rect 199436 197956 199442 198008
rect 151170 197928 151176 197940
rect 134168 197900 151176 197928
rect 132218 197820 132224 197872
rect 132276 197860 132282 197872
rect 134168 197860 134196 197900
rect 151170 197888 151176 197900
rect 151228 197888 151234 197940
rect 163314 197888 163320 197940
rect 163372 197928 163378 197940
rect 163498 197928 163504 197940
rect 163372 197900 163504 197928
rect 163372 197888 163378 197900
rect 163498 197888 163504 197900
rect 163556 197888 163562 197940
rect 171870 197928 171876 197940
rect 166966 197900 171876 197928
rect 132276 197832 134196 197860
rect 132276 197820 132282 197832
rect 138290 197820 138296 197872
rect 138348 197860 138354 197872
rect 149422 197860 149428 197872
rect 138348 197832 149428 197860
rect 138348 197820 138354 197832
rect 149422 197820 149428 197832
rect 149480 197820 149486 197872
rect 155034 197820 155040 197872
rect 155092 197860 155098 197872
rect 166966 197860 166994 197900
rect 171870 197888 171876 197900
rect 171928 197888 171934 197940
rect 173526 197888 173532 197940
rect 173584 197928 173590 197940
rect 193858 197928 193864 197940
rect 173584 197900 193864 197928
rect 173584 197888 173590 197900
rect 193858 197888 193864 197900
rect 193916 197888 193922 197940
rect 155092 197832 166994 197860
rect 155092 197820 155098 197832
rect 170490 197820 170496 197872
rect 170548 197860 170554 197872
rect 187694 197860 187700 197872
rect 170548 197832 187700 197860
rect 170548 197820 170554 197832
rect 187694 197820 187700 197832
rect 187752 197820 187758 197872
rect 126146 197752 126152 197804
rect 126204 197792 126210 197804
rect 144822 197792 144828 197804
rect 126204 197764 131114 197792
rect 126204 197752 126210 197764
rect 131086 197724 131114 197764
rect 137848 197764 144828 197792
rect 137848 197724 137876 197764
rect 144822 197752 144828 197764
rect 144880 197752 144886 197804
rect 170214 197752 170220 197804
rect 170272 197792 170278 197804
rect 186682 197792 186688 197804
rect 170272 197764 186688 197792
rect 170272 197752 170278 197764
rect 186682 197752 186688 197764
rect 186740 197752 186746 197804
rect 131086 197696 137876 197724
rect 163774 197684 163780 197736
rect 163832 197724 163838 197736
rect 189074 197724 189080 197736
rect 163832 197696 189080 197724
rect 163832 197684 163838 197696
rect 189074 197684 189080 197696
rect 189132 197684 189138 197736
rect 131022 197616 131028 197668
rect 131080 197656 131086 197668
rect 138290 197656 138296 197668
rect 131080 197628 138296 197656
rect 131080 197616 131086 197628
rect 138290 197616 138296 197628
rect 138348 197616 138354 197668
rect 171778 197616 171784 197668
rect 171836 197656 171842 197668
rect 180426 197656 180432 197668
rect 171836 197628 180432 197656
rect 171836 197616 171842 197628
rect 180426 197616 180432 197628
rect 180484 197616 180490 197668
rect 165614 197548 165620 197600
rect 165672 197588 165678 197600
rect 181622 197588 181628 197600
rect 165672 197560 181628 197588
rect 165672 197548 165678 197560
rect 181622 197548 181628 197560
rect 181680 197548 181686 197600
rect 145466 197480 145472 197532
rect 145524 197520 145530 197532
rect 147674 197520 147680 197532
rect 145524 197492 147680 197520
rect 145524 197480 145530 197492
rect 147674 197480 147680 197492
rect 147732 197480 147738 197532
rect 171318 197480 171324 197532
rect 171376 197520 171382 197532
rect 172422 197520 172428 197532
rect 171376 197492 172428 197520
rect 171376 197480 171382 197492
rect 172422 197480 172428 197492
rect 172480 197480 172486 197532
rect 120442 197412 120448 197464
rect 120500 197452 120506 197464
rect 144178 197452 144184 197464
rect 120500 197424 144184 197452
rect 120500 197412 120506 197424
rect 144178 197412 144184 197424
rect 144236 197412 144242 197464
rect 171502 197412 171508 197464
rect 171560 197452 171566 197464
rect 172146 197452 172152 197464
rect 171560 197424 172152 197452
rect 171560 197412 171566 197424
rect 172146 197412 172152 197424
rect 172204 197412 172210 197464
rect 117314 197344 117320 197396
rect 117372 197384 117378 197396
rect 138934 197384 138940 197396
rect 117372 197356 138940 197384
rect 117372 197344 117378 197356
rect 138934 197344 138940 197356
rect 138992 197344 138998 197396
rect 174078 197344 174084 197396
rect 174136 197384 174142 197396
rect 174446 197384 174452 197396
rect 174136 197356 174452 197384
rect 174136 197344 174142 197356
rect 174446 197344 174452 197356
rect 174504 197344 174510 197396
rect 130562 197276 130568 197328
rect 130620 197316 130626 197328
rect 150526 197316 150532 197328
rect 130620 197288 150532 197316
rect 130620 197276 130626 197288
rect 150526 197276 150532 197288
rect 150584 197276 150590 197328
rect 164786 197276 164792 197328
rect 164844 197316 164850 197328
rect 199010 197316 199016 197328
rect 164844 197288 199016 197316
rect 164844 197276 164850 197288
rect 199010 197276 199016 197288
rect 199068 197276 199074 197328
rect 112898 197208 112904 197260
rect 112956 197248 112962 197260
rect 112956 197220 140314 197248
rect 112956 197208 112962 197220
rect 117130 197140 117136 197192
rect 117188 197180 117194 197192
rect 120442 197180 120448 197192
rect 117188 197152 120448 197180
rect 117188 197140 117194 197152
rect 120442 197140 120448 197152
rect 120500 197140 120506 197192
rect 132954 197140 132960 197192
rect 133012 197180 133018 197192
rect 140038 197180 140044 197192
rect 133012 197152 140044 197180
rect 133012 197140 133018 197152
rect 140038 197140 140044 197152
rect 140096 197140 140102 197192
rect 140286 197180 140314 197220
rect 164142 197208 164148 197260
rect 164200 197248 164206 197260
rect 193214 197248 193220 197260
rect 164200 197220 193220 197248
rect 164200 197208 164206 197220
rect 193214 197208 193220 197220
rect 193272 197208 193278 197260
rect 142890 197180 142896 197192
rect 140286 197152 142896 197180
rect 142890 197140 142896 197152
rect 142948 197140 142954 197192
rect 164418 197140 164424 197192
rect 164476 197180 164482 197192
rect 199654 197180 199660 197192
rect 164476 197152 199660 197180
rect 164476 197140 164482 197152
rect 199654 197140 199660 197152
rect 199712 197140 199718 197192
rect 111610 197072 111616 197124
rect 111668 197112 111674 197124
rect 143258 197112 143264 197124
rect 111668 197084 143264 197112
rect 111668 197072 111674 197084
rect 143258 197072 143264 197084
rect 143316 197072 143322 197124
rect 147582 197072 147588 197124
rect 147640 197112 147646 197124
rect 154850 197112 154856 197124
rect 147640 197084 154856 197112
rect 147640 197072 147646 197084
rect 154850 197072 154856 197084
rect 154908 197072 154914 197124
rect 163498 197072 163504 197124
rect 163556 197112 163562 197124
rect 197446 197112 197452 197124
rect 163556 197084 197452 197112
rect 163556 197072 163562 197084
rect 197446 197072 197452 197084
rect 197504 197072 197510 197124
rect 117038 197004 117044 197056
rect 117096 197044 117102 197056
rect 148594 197044 148600 197056
rect 117096 197016 148600 197044
rect 117096 197004 117102 197016
rect 148594 197004 148600 197016
rect 148652 197004 148658 197056
rect 160830 197004 160836 197056
rect 160888 197044 160894 197056
rect 194686 197044 194692 197056
rect 160888 197016 194692 197044
rect 160888 197004 160894 197016
rect 194686 197004 194692 197016
rect 194744 197004 194750 197056
rect 112714 196936 112720 196988
rect 112772 196976 112778 196988
rect 132770 196976 132776 196988
rect 112772 196948 132776 196976
rect 112772 196936 112778 196948
rect 132770 196936 132776 196948
rect 132828 196936 132834 196988
rect 133138 196936 133144 196988
rect 133196 196976 133202 196988
rect 142522 196976 142528 196988
rect 133196 196948 142528 196976
rect 133196 196936 133202 196948
rect 142522 196936 142528 196948
rect 142580 196936 142586 196988
rect 163682 196936 163688 196988
rect 163740 196976 163746 196988
rect 197538 196976 197544 196988
rect 163740 196948 197544 196976
rect 163740 196936 163746 196948
rect 197538 196936 197544 196948
rect 197596 196936 197602 196988
rect 110322 196868 110328 196920
rect 110380 196908 110386 196920
rect 142798 196908 142804 196920
rect 110380 196880 142804 196908
rect 110380 196868 110386 196880
rect 142798 196868 142804 196880
rect 142856 196868 142862 196920
rect 160370 196868 160376 196920
rect 160428 196908 160434 196920
rect 194870 196908 194876 196920
rect 160428 196880 194876 196908
rect 160428 196868 160434 196880
rect 194870 196868 194876 196880
rect 194928 196868 194934 196920
rect 111334 196800 111340 196852
rect 111392 196840 111398 196852
rect 132954 196840 132960 196852
rect 111392 196812 132960 196840
rect 111392 196800 111398 196812
rect 132954 196800 132960 196812
rect 133012 196800 133018 196852
rect 140130 196840 140136 196852
rect 133064 196812 140136 196840
rect 106826 196732 106832 196784
rect 106884 196772 106890 196784
rect 133064 196772 133092 196812
rect 140130 196800 140136 196812
rect 140188 196800 140194 196852
rect 177850 196800 177856 196852
rect 177908 196840 177914 196852
rect 196342 196840 196348 196852
rect 177908 196812 196348 196840
rect 177908 196800 177914 196812
rect 196342 196800 196348 196812
rect 196400 196800 196406 196852
rect 106884 196744 133092 196772
rect 106884 196732 106890 196744
rect 140038 196732 140044 196784
rect 140096 196772 140102 196784
rect 143718 196772 143724 196784
rect 140096 196744 143724 196772
rect 140096 196732 140102 196744
rect 143718 196732 143724 196744
rect 143776 196732 143782 196784
rect 158990 196732 158996 196784
rect 159048 196772 159054 196784
rect 187786 196772 187792 196784
rect 159048 196744 187792 196772
rect 159048 196732 159054 196744
rect 187786 196732 187792 196744
rect 187844 196732 187850 196784
rect 109770 196664 109776 196716
rect 109828 196704 109834 196716
rect 133138 196704 133144 196716
rect 109828 196676 133144 196704
rect 109828 196664 109834 196676
rect 133138 196664 133144 196676
rect 133196 196664 133202 196716
rect 171778 196664 171784 196716
rect 171836 196704 171842 196716
rect 197630 196704 197636 196716
rect 171836 196676 197636 196704
rect 171836 196664 171842 196676
rect 197630 196664 197636 196676
rect 197688 196664 197694 196716
rect 106090 196596 106096 196648
rect 106148 196636 106154 196648
rect 139578 196636 139584 196648
rect 106148 196608 139584 196636
rect 106148 196596 106154 196608
rect 139578 196596 139584 196608
rect 139636 196596 139642 196648
rect 159542 196596 159548 196648
rect 159600 196636 159606 196648
rect 193398 196636 193404 196648
rect 159600 196608 193404 196636
rect 159600 196596 159606 196608
rect 193398 196596 193404 196608
rect 193456 196596 193462 196648
rect 180242 196568 180248 196580
rect 166920 196540 180248 196568
rect 123386 196460 123392 196512
rect 123444 196500 123450 196512
rect 123444 196472 124214 196500
rect 123444 196460 123450 196472
rect 124186 196432 124214 196472
rect 133322 196460 133328 196512
rect 133380 196500 133386 196512
rect 144086 196500 144092 196512
rect 133380 196472 144092 196500
rect 133380 196460 133386 196472
rect 144086 196460 144092 196472
rect 144144 196460 144150 196512
rect 162302 196460 162308 196512
rect 162360 196500 162366 196512
rect 166920 196500 166948 196540
rect 180242 196528 180248 196540
rect 180300 196528 180306 196580
rect 162360 196472 166948 196500
rect 162360 196460 162366 196472
rect 143442 196432 143448 196444
rect 124186 196404 143448 196432
rect 143442 196392 143448 196404
rect 143500 196392 143506 196444
rect 132770 196256 132776 196308
rect 132828 196296 132834 196308
rect 133322 196296 133328 196308
rect 132828 196268 133328 196296
rect 132828 196256 132834 196268
rect 133322 196256 133328 196268
rect 133380 196256 133386 196308
rect 147950 196188 147956 196240
rect 148008 196228 148014 196240
rect 157886 196228 157892 196240
rect 148008 196200 157892 196228
rect 148008 196188 148014 196200
rect 157886 196188 157892 196200
rect 157944 196188 157950 196240
rect 165614 196188 165620 196240
rect 165672 196228 165678 196240
rect 166166 196228 166172 196240
rect 165672 196200 166172 196228
rect 165672 196188 165678 196200
rect 166166 196188 166172 196200
rect 166224 196188 166230 196240
rect 134150 196052 134156 196104
rect 134208 196092 134214 196104
rect 134702 196092 134708 196104
rect 134208 196064 134708 196092
rect 134208 196052 134214 196064
rect 134702 196052 134708 196064
rect 134760 196052 134766 196104
rect 133690 195984 133696 196036
rect 133748 196024 133754 196036
rect 135990 196024 135996 196036
rect 133748 195996 135996 196024
rect 133748 195984 133754 195996
rect 135990 195984 135996 195996
rect 136048 195984 136054 196036
rect 122650 195916 122656 195968
rect 122708 195956 122714 195968
rect 154298 195956 154304 195968
rect 122708 195928 154304 195956
rect 122708 195916 122714 195928
rect 154298 195916 154304 195928
rect 154356 195916 154362 195968
rect 172146 195916 172152 195968
rect 172204 195956 172210 195968
rect 190638 195956 190644 195968
rect 172204 195928 190644 195956
rect 172204 195916 172210 195928
rect 190638 195916 190644 195928
rect 190696 195916 190702 195968
rect 111426 195848 111432 195900
rect 111484 195888 111490 195900
rect 133690 195888 133696 195900
rect 111484 195860 133696 195888
rect 111484 195848 111490 195860
rect 133690 195848 133696 195860
rect 133748 195848 133754 195900
rect 133984 195860 134196 195888
rect 114094 195780 114100 195832
rect 114152 195820 114158 195832
rect 133984 195820 134012 195860
rect 114152 195792 134012 195820
rect 134168 195820 134196 195860
rect 151998 195848 152004 195900
rect 152056 195888 152062 195900
rect 152642 195888 152648 195900
rect 152056 195860 152648 195888
rect 152056 195848 152062 195860
rect 152642 195848 152648 195860
rect 152700 195848 152706 195900
rect 172422 195848 172428 195900
rect 172480 195888 172486 195900
rect 190730 195888 190736 195900
rect 172480 195860 190736 195888
rect 172480 195848 172486 195860
rect 190730 195848 190736 195860
rect 190788 195848 190794 195900
rect 145006 195820 145012 195832
rect 134168 195792 145012 195820
rect 114152 195780 114158 195792
rect 145006 195780 145012 195792
rect 145064 195780 145070 195832
rect 156966 195780 156972 195832
rect 157024 195820 157030 195832
rect 166258 195820 166264 195832
rect 157024 195792 166264 195820
rect 157024 195780 157030 195792
rect 166258 195780 166264 195792
rect 166316 195780 166322 195832
rect 169754 195780 169760 195832
rect 169812 195820 169818 195832
rect 192570 195820 192576 195832
rect 169812 195792 192576 195820
rect 169812 195780 169818 195792
rect 192570 195780 192576 195792
rect 192628 195780 192634 195832
rect 103054 195712 103060 195764
rect 103112 195752 103118 195764
rect 134334 195752 134340 195764
rect 103112 195724 134340 195752
rect 103112 195712 103118 195724
rect 134334 195712 134340 195724
rect 134392 195712 134398 195764
rect 135990 195712 135996 195764
rect 136048 195752 136054 195764
rect 142430 195752 142436 195764
rect 136048 195724 142436 195752
rect 136048 195712 136054 195724
rect 142430 195712 142436 195724
rect 142488 195712 142494 195764
rect 158070 195712 158076 195764
rect 158128 195752 158134 195764
rect 191834 195752 191840 195764
rect 158128 195724 191840 195752
rect 158128 195712 158134 195724
rect 191834 195712 191840 195724
rect 191892 195712 191898 195764
rect 107010 195644 107016 195696
rect 107068 195684 107074 195696
rect 137922 195684 137928 195696
rect 107068 195656 137928 195684
rect 107068 195644 107074 195656
rect 137922 195644 137928 195656
rect 137980 195644 137986 195696
rect 165706 195644 165712 195696
rect 165764 195684 165770 195696
rect 196066 195684 196072 195696
rect 165764 195656 196072 195684
rect 165764 195644 165770 195656
rect 196066 195644 196072 195656
rect 196124 195644 196130 195696
rect 110230 195576 110236 195628
rect 110288 195616 110294 195628
rect 143074 195616 143080 195628
rect 110288 195588 143080 195616
rect 110288 195576 110294 195588
rect 143074 195576 143080 195588
rect 143132 195576 143138 195628
rect 161566 195576 161572 195628
rect 161624 195616 161630 195628
rect 194594 195616 194600 195628
rect 161624 195588 194600 195616
rect 161624 195576 161630 195588
rect 194594 195576 194600 195588
rect 194652 195576 194658 195628
rect 114278 195508 114284 195560
rect 114336 195548 114342 195560
rect 147122 195548 147128 195560
rect 114336 195520 147128 195548
rect 114336 195508 114342 195520
rect 147122 195508 147128 195520
rect 147180 195508 147186 195560
rect 166258 195508 166264 195560
rect 166316 195548 166322 195560
rect 190454 195548 190460 195560
rect 166316 195520 190460 195548
rect 166316 195508 166322 195520
rect 190454 195508 190460 195520
rect 190512 195508 190518 195560
rect 118878 195440 118884 195492
rect 118936 195480 118942 195492
rect 153102 195480 153108 195492
rect 118936 195452 153108 195480
rect 118936 195440 118942 195452
rect 153102 195440 153108 195452
rect 153160 195440 153166 195492
rect 162210 195440 162216 195492
rect 162268 195480 162274 195492
rect 196158 195480 196164 195492
rect 162268 195452 196164 195480
rect 162268 195440 162274 195452
rect 196158 195440 196164 195452
rect 196216 195440 196222 195492
rect 105630 195372 105636 195424
rect 105688 195412 105694 195424
rect 117314 195412 117320 195424
rect 105688 195384 117320 195412
rect 105688 195372 105694 195384
rect 117314 195372 117320 195384
rect 117372 195372 117378 195424
rect 138658 195372 138664 195424
rect 138716 195412 138722 195424
rect 140774 195412 140780 195424
rect 138716 195384 140780 195412
rect 138716 195372 138722 195384
rect 140774 195372 140780 195384
rect 140832 195372 140838 195424
rect 157334 195372 157340 195424
rect 157392 195412 157398 195424
rect 190546 195412 190552 195424
rect 157392 195384 190552 195412
rect 157392 195372 157398 195384
rect 190546 195372 190552 195384
rect 190604 195372 190610 195424
rect 105814 195304 105820 195356
rect 105872 195344 105878 195356
rect 139854 195344 139860 195356
rect 105872 195316 139860 195344
rect 105872 195304 105878 195316
rect 139854 195304 139860 195316
rect 139912 195304 139918 195356
rect 158714 195304 158720 195356
rect 158772 195344 158778 195356
rect 191926 195344 191932 195356
rect 158772 195316 191932 195344
rect 158772 195304 158778 195316
rect 191926 195304 191932 195316
rect 191984 195304 191990 195356
rect 112622 195236 112628 195288
rect 112680 195276 112686 195288
rect 145098 195276 145104 195288
rect 112680 195248 145104 195276
rect 112680 195236 112686 195248
rect 145098 195236 145104 195248
rect 145156 195236 145162 195288
rect 157242 195236 157248 195288
rect 157300 195276 157306 195288
rect 157794 195276 157800 195288
rect 157300 195248 157800 195276
rect 157300 195236 157306 195248
rect 157794 195236 157800 195248
rect 157852 195236 157858 195288
rect 161842 195236 161848 195288
rect 161900 195276 161906 195288
rect 194778 195276 194784 195288
rect 161900 195248 194784 195276
rect 161900 195236 161906 195248
rect 194778 195236 194784 195248
rect 194836 195236 194842 195288
rect 118510 195168 118516 195220
rect 118568 195208 118574 195220
rect 148962 195208 148968 195220
rect 118568 195180 148968 195208
rect 118568 195168 118574 195180
rect 148962 195168 148968 195180
rect 149020 195168 149026 195220
rect 164970 195168 164976 195220
rect 165028 195208 165034 195220
rect 165154 195208 165160 195220
rect 165028 195180 165160 195208
rect 165028 195168 165034 195180
rect 165154 195168 165160 195180
rect 165212 195168 165218 195220
rect 169018 195168 169024 195220
rect 169076 195208 169082 195220
rect 169570 195208 169576 195220
rect 169076 195180 169576 195208
rect 169076 195168 169082 195180
rect 169570 195168 169576 195180
rect 169628 195168 169634 195220
rect 189166 195208 189172 195220
rect 177776 195180 189172 195208
rect 148226 195100 148232 195152
rect 148284 195140 148290 195152
rect 148778 195140 148784 195152
rect 148284 195112 148784 195140
rect 148284 195100 148290 195112
rect 148778 195100 148784 195112
rect 148836 195100 148842 195152
rect 168742 195100 168748 195152
rect 168800 195140 168806 195152
rect 169202 195140 169208 195152
rect 168800 195112 169208 195140
rect 168800 195100 168806 195112
rect 169202 195100 169208 195112
rect 169260 195100 169266 195152
rect 171870 194896 171876 194948
rect 171928 194936 171934 194948
rect 177776 194936 177804 195180
rect 189166 195168 189172 195180
rect 189224 195168 189230 195220
rect 188154 195140 188160 195152
rect 171928 194908 177804 194936
rect 177868 195112 188160 195140
rect 171928 194896 171934 194908
rect 171134 194828 171140 194880
rect 171192 194868 171198 194880
rect 177868 194868 177896 195112
rect 188154 195100 188160 195112
rect 188212 195100 188218 195152
rect 171192 194840 177896 194868
rect 171192 194828 171198 194840
rect 124858 194760 124864 194812
rect 124916 194800 124922 194812
rect 137646 194800 137652 194812
rect 124916 194772 137652 194800
rect 124916 194760 124922 194772
rect 137646 194760 137652 194772
rect 137704 194760 137710 194812
rect 166994 194624 167000 194676
rect 167052 194664 167058 194676
rect 184198 194664 184204 194676
rect 167052 194636 184204 194664
rect 167052 194624 167058 194636
rect 184198 194624 184204 194636
rect 184256 194624 184262 194676
rect 122098 194488 122104 194540
rect 122156 194528 122162 194540
rect 149422 194528 149428 194540
rect 122156 194500 149428 194528
rect 122156 194488 122162 194500
rect 149422 194488 149428 194500
rect 149480 194488 149486 194540
rect 166994 194488 167000 194540
rect 167052 194528 167058 194540
rect 168650 194528 168656 194540
rect 167052 194500 168656 194528
rect 167052 194488 167058 194500
rect 168650 194488 168656 194500
rect 168708 194488 168714 194540
rect 104158 194420 104164 194472
rect 104216 194460 104222 194472
rect 132586 194460 132592 194472
rect 104216 194432 132592 194460
rect 104216 194420 104222 194432
rect 132586 194420 132592 194432
rect 132644 194420 132650 194472
rect 111058 194352 111064 194404
rect 111116 194392 111122 194404
rect 141786 194392 141792 194404
rect 111116 194364 141792 194392
rect 111116 194352 111122 194364
rect 141786 194352 141792 194364
rect 141844 194352 141850 194404
rect 166074 194352 166080 194404
rect 166132 194392 166138 194404
rect 182910 194392 182916 194404
rect 166132 194364 182916 194392
rect 166132 194352 166138 194364
rect 182910 194352 182916 194364
rect 182968 194352 182974 194404
rect 108758 194284 108764 194336
rect 108816 194324 108822 194336
rect 136910 194324 136916 194336
rect 108816 194296 136916 194324
rect 108816 194284 108822 194296
rect 136910 194284 136916 194296
rect 136968 194284 136974 194336
rect 138750 194284 138756 194336
rect 138808 194324 138814 194336
rect 138934 194324 138940 194336
rect 138808 194296 138940 194324
rect 138808 194284 138814 194296
rect 138934 194284 138940 194296
rect 138992 194284 138998 194336
rect 104710 194216 104716 194268
rect 104768 194256 104774 194268
rect 136358 194256 136364 194268
rect 104768 194228 136364 194256
rect 104768 194216 104774 194228
rect 136358 194216 136364 194228
rect 136416 194216 136422 194268
rect 161474 194216 161480 194268
rect 161532 194256 161538 194268
rect 161750 194256 161756 194268
rect 161532 194228 161756 194256
rect 161532 194216 161538 194228
rect 161750 194216 161756 194228
rect 161808 194216 161814 194268
rect 168006 194216 168012 194268
rect 168064 194256 168070 194268
rect 201586 194256 201592 194268
rect 168064 194228 201592 194256
rect 168064 194216 168070 194228
rect 201586 194216 201592 194228
rect 201644 194216 201650 194268
rect 104342 194148 104348 194200
rect 104400 194188 104406 194200
rect 135714 194188 135720 194200
rect 104400 194160 135720 194188
rect 104400 194148 104406 194160
rect 135714 194148 135720 194160
rect 135772 194148 135778 194200
rect 168558 194148 168564 194200
rect 168616 194188 168622 194200
rect 203334 194188 203340 194200
rect 168616 194160 203340 194188
rect 168616 194148 168622 194160
rect 203334 194148 203340 194160
rect 203392 194148 203398 194200
rect 104526 194080 104532 194132
rect 104584 194120 104590 194132
rect 136082 194120 136088 194132
rect 104584 194092 136088 194120
rect 104584 194080 104590 194092
rect 136082 194080 136088 194092
rect 136140 194080 136146 194132
rect 169110 194080 169116 194132
rect 169168 194120 169174 194132
rect 203242 194120 203248 194132
rect 169168 194092 203248 194120
rect 169168 194080 169174 194092
rect 203242 194080 203248 194092
rect 203300 194080 203306 194132
rect 100570 194012 100576 194064
rect 100628 194052 100634 194064
rect 125226 194052 125232 194064
rect 100628 194024 125232 194052
rect 100628 194012 100634 194024
rect 125226 194012 125232 194024
rect 125284 194012 125290 194064
rect 167178 194012 167184 194064
rect 167236 194052 167242 194064
rect 202046 194052 202052 194064
rect 167236 194024 202052 194052
rect 167236 194012 167242 194024
rect 202046 194012 202052 194024
rect 202104 194012 202110 194064
rect 101674 193944 101680 193996
rect 101732 193984 101738 193996
rect 134058 193984 134064 193996
rect 101732 193956 134064 193984
rect 101732 193944 101738 193956
rect 134058 193944 134064 193956
rect 134116 193944 134122 193996
rect 153930 193944 153936 193996
rect 153988 193984 153994 193996
rect 205818 193984 205824 193996
rect 153988 193956 205824 193984
rect 153988 193944 153994 193956
rect 205818 193944 205824 193956
rect 205876 193944 205882 193996
rect 103146 193876 103152 193928
rect 103204 193916 103210 193928
rect 135530 193916 135536 193928
rect 103204 193888 135536 193916
rect 103204 193876 103210 193888
rect 135530 193876 135536 193888
rect 135588 193876 135594 193928
rect 161842 193876 161848 193928
rect 161900 193916 161906 193928
rect 205726 193916 205732 193928
rect 161900 193888 205732 193916
rect 161900 193876 161906 193888
rect 205726 193876 205732 193888
rect 205784 193876 205790 193928
rect 105906 193808 105912 193860
rect 105964 193848 105970 193860
rect 140498 193848 140504 193860
rect 105964 193820 140504 193848
rect 105964 193808 105970 193820
rect 140498 193808 140504 193820
rect 140556 193808 140562 193860
rect 151262 193808 151268 193860
rect 151320 193848 151326 193860
rect 206094 193848 206100 193860
rect 151320 193820 206100 193848
rect 151320 193808 151326 193820
rect 206094 193808 206100 193820
rect 206152 193808 206158 193860
rect 112530 193740 112536 193792
rect 112588 193780 112594 193792
rect 117682 193780 117688 193792
rect 112588 193752 117688 193780
rect 112588 193740 112594 193752
rect 117682 193740 117688 193752
rect 117740 193740 117746 193792
rect 122006 193672 122012 193724
rect 122064 193712 122070 193724
rect 147950 193712 147956 193724
rect 122064 193684 147956 193712
rect 122064 193672 122070 193684
rect 147950 193672 147956 193684
rect 148008 193672 148014 193724
rect 123202 193604 123208 193656
rect 123260 193644 123266 193656
rect 146018 193644 146024 193656
rect 123260 193616 146024 193644
rect 123260 193604 123266 193616
rect 146018 193604 146024 193616
rect 146076 193604 146082 193656
rect 176010 193536 176016 193588
rect 176068 193576 176074 193588
rect 188706 193576 188712 193588
rect 176068 193548 188712 193576
rect 176068 193536 176074 193548
rect 188706 193536 188712 193548
rect 188764 193536 188770 193588
rect 105722 193128 105728 193180
rect 105780 193168 105786 193180
rect 137002 193168 137008 193180
rect 105780 193140 137008 193168
rect 105780 193128 105786 193140
rect 137002 193128 137008 193140
rect 137060 193128 137066 193180
rect 156322 193128 156328 193180
rect 156380 193168 156386 193180
rect 183094 193168 183100 193180
rect 156380 193140 183100 193168
rect 156380 193128 156386 193140
rect 183094 193128 183100 193140
rect 183152 193128 183158 193180
rect 188338 193128 188344 193180
rect 188396 193168 188402 193180
rect 580166 193168 580172 193180
rect 188396 193140 580172 193168
rect 188396 193128 188402 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 108298 193060 108304 193112
rect 108356 193100 108362 193112
rect 140682 193100 140688 193112
rect 108356 193072 140688 193100
rect 108356 193060 108362 193072
rect 140682 193060 140688 193072
rect 140740 193060 140746 193112
rect 176838 193060 176844 193112
rect 176896 193100 176902 193112
rect 204346 193100 204352 193112
rect 176896 193072 204352 193100
rect 176896 193060 176902 193072
rect 204346 193060 204352 193072
rect 204404 193060 204410 193112
rect 110138 192992 110144 193044
rect 110196 193032 110202 193044
rect 144730 193032 144736 193044
rect 110196 193004 144736 193032
rect 110196 192992 110202 193004
rect 144730 192992 144736 193004
rect 144788 192992 144794 193044
rect 165522 192992 165528 193044
rect 165580 193032 165586 193044
rect 192478 193032 192484 193044
rect 165580 193004 192484 193032
rect 165580 192992 165586 193004
rect 192478 192992 192484 193004
rect 192536 192992 192542 193044
rect 111150 192924 111156 192976
rect 111208 192964 111214 192976
rect 144362 192964 144368 192976
rect 111208 192936 144368 192964
rect 111208 192924 111214 192936
rect 144362 192924 144368 192936
rect 144420 192924 144426 192976
rect 153378 192924 153384 192976
rect 153436 192964 153442 192976
rect 154022 192964 154028 192976
rect 153436 192936 154028 192964
rect 153436 192924 153442 192936
rect 154022 192924 154028 192936
rect 154080 192924 154086 192976
rect 170122 192924 170128 192976
rect 170180 192964 170186 192976
rect 201770 192964 201776 192976
rect 170180 192936 201776 192964
rect 170180 192924 170186 192936
rect 201770 192924 201776 192936
rect 201828 192924 201834 192976
rect 110046 192856 110052 192908
rect 110104 192896 110110 192908
rect 143994 192896 144000 192908
rect 110104 192868 144000 192896
rect 110104 192856 110110 192868
rect 143994 192856 144000 192868
rect 144052 192856 144058 192908
rect 167270 192856 167276 192908
rect 167328 192896 167334 192908
rect 168282 192896 168288 192908
rect 167328 192868 168288 192896
rect 167328 192856 167334 192868
rect 168282 192856 168288 192868
rect 168340 192856 168346 192908
rect 174446 192856 174452 192908
rect 174504 192896 174510 192908
rect 205910 192896 205916 192908
rect 174504 192868 205916 192896
rect 174504 192856 174510 192868
rect 205910 192856 205916 192868
rect 205968 192856 205974 192908
rect 105998 192788 106004 192840
rect 106056 192828 106062 192840
rect 131574 192828 131580 192840
rect 106056 192800 131580 192828
rect 106056 192788 106062 192800
rect 131574 192788 131580 192800
rect 131632 192788 131638 192840
rect 163038 192788 163044 192840
rect 163096 192828 163102 192840
rect 163406 192828 163412 192840
rect 163096 192800 163412 192828
rect 163096 192788 163102 192800
rect 163406 192788 163412 192800
rect 163464 192788 163470 192840
rect 172698 192788 172704 192840
rect 172756 192828 172762 192840
rect 206002 192828 206008 192840
rect 172756 192800 206008 192828
rect 172756 192788 172762 192800
rect 206002 192788 206008 192800
rect 206060 192788 206066 192840
rect 115382 192720 115388 192772
rect 115440 192760 115446 192772
rect 149790 192760 149796 192772
rect 115440 192732 149796 192760
rect 115440 192720 115446 192732
rect 149790 192720 149796 192732
rect 149848 192720 149854 192772
rect 164234 192720 164240 192772
rect 164292 192760 164298 192772
rect 195974 192760 195980 192772
rect 164292 192732 195980 192760
rect 164292 192720 164298 192732
rect 195974 192720 195980 192732
rect 196032 192720 196038 192772
rect 104250 192652 104256 192704
rect 104308 192692 104314 192704
rect 136542 192692 136548 192704
rect 104308 192664 136548 192692
rect 104308 192652 104314 192664
rect 136542 192652 136548 192664
rect 136600 192652 136606 192704
rect 169478 192652 169484 192704
rect 169536 192692 169542 192704
rect 202874 192692 202880 192704
rect 169536 192664 202880 192692
rect 169536 192652 169542 192664
rect 202874 192652 202880 192664
rect 202932 192652 202938 192704
rect 109862 192584 109868 192636
rect 109920 192624 109926 192636
rect 144546 192624 144552 192636
rect 109920 192596 144552 192624
rect 109920 192584 109926 192596
rect 144546 192584 144552 192596
rect 144604 192584 144610 192636
rect 168190 192584 168196 192636
rect 168248 192624 168254 192636
rect 201678 192624 201684 192636
rect 168248 192596 201684 192624
rect 168248 192584 168254 192596
rect 201678 192584 201684 192596
rect 201736 192584 201742 192636
rect 102778 192516 102784 192568
rect 102836 192556 102842 192568
rect 136818 192556 136824 192568
rect 102836 192528 136824 192556
rect 102836 192516 102842 192528
rect 136818 192516 136824 192528
rect 136876 192516 136882 192568
rect 178678 192516 178684 192568
rect 178736 192556 178742 192568
rect 200298 192556 200304 192568
rect 178736 192528 200304 192556
rect 178736 192516 178742 192528
rect 200298 192516 200304 192528
rect 200356 192516 200362 192568
rect 108574 192448 108580 192500
rect 108632 192488 108638 192500
rect 141970 192488 141976 192500
rect 108632 192460 141976 192488
rect 108632 192448 108638 192460
rect 141970 192448 141976 192460
rect 142028 192448 142034 192500
rect 166810 192448 166816 192500
rect 166868 192488 166874 192500
rect 200758 192488 200764 192500
rect 166868 192460 200764 192488
rect 166868 192448 166874 192460
rect 200758 192448 200764 192460
rect 200816 192448 200822 192500
rect 107470 192380 107476 192432
rect 107528 192420 107534 192432
rect 137738 192420 137744 192432
rect 107528 192392 137744 192420
rect 107528 192380 107534 192392
rect 137738 192380 137744 192392
rect 137796 192380 137802 192432
rect 156230 192380 156236 192432
rect 156288 192420 156294 192432
rect 181530 192420 181536 192432
rect 156288 192392 181536 192420
rect 156288 192380 156294 192392
rect 181530 192380 181536 192392
rect 181588 192380 181594 192432
rect 157518 192312 157524 192364
rect 157576 192352 157582 192364
rect 181438 192352 181444 192364
rect 157576 192324 181444 192352
rect 157576 192312 157582 192324
rect 181438 192312 181444 192324
rect 181496 192312 181502 192364
rect 157426 192244 157432 192296
rect 157484 192284 157490 192296
rect 158254 192284 158260 192296
rect 157484 192256 158260 192284
rect 157484 192244 157490 192256
rect 158254 192244 158260 192256
rect 158312 192244 158318 192296
rect 165798 192244 165804 192296
rect 165856 192284 165862 192296
rect 166718 192284 166724 192296
rect 165856 192256 166724 192284
rect 165856 192244 165862 192256
rect 166718 192244 166724 192256
rect 166776 192244 166782 192296
rect 158990 191224 158996 191276
rect 159048 191264 159054 191276
rect 159910 191264 159916 191276
rect 159048 191236 159916 191264
rect 159048 191224 159054 191236
rect 159910 191224 159916 191236
rect 159968 191224 159974 191276
rect 164326 191224 164332 191276
rect 164384 191264 164390 191276
rect 164602 191264 164608 191276
rect 164384 191236 164608 191264
rect 164384 191224 164390 191236
rect 164602 191224 164608 191236
rect 164660 191224 164666 191276
rect 167086 191224 167092 191276
rect 167144 191264 167150 191276
rect 168098 191264 168104 191276
rect 167144 191236 168104 191264
rect 167144 191224 167150 191236
rect 168098 191224 168104 191236
rect 168156 191224 168162 191276
rect 150526 191156 150532 191208
rect 150584 191196 150590 191208
rect 151814 191196 151820 191208
rect 150584 191168 151820 191196
rect 150584 191156 150590 191168
rect 151814 191156 151820 191168
rect 151872 191156 151878 191208
rect 173986 191156 173992 191208
rect 174044 191196 174050 191208
rect 174998 191196 175004 191208
rect 174044 191168 175004 191196
rect 174044 191156 174050 191168
rect 174998 191156 175004 191168
rect 175056 191156 175062 191208
rect 146754 191088 146760 191140
rect 146812 191128 146818 191140
rect 147306 191128 147312 191140
rect 146812 191100 147312 191128
rect 146812 191088 146818 191100
rect 147306 191088 147312 191100
rect 147364 191088 147370 191140
rect 151722 191088 151728 191140
rect 151780 191128 151786 191140
rect 152182 191128 152188 191140
rect 151780 191100 152188 191128
rect 151780 191088 151786 191100
rect 152182 191088 152188 191100
rect 152240 191088 152246 191140
rect 157610 191088 157616 191140
rect 157668 191128 157674 191140
rect 158438 191128 158444 191140
rect 157668 191100 158444 191128
rect 157668 191088 157674 191100
rect 158438 191088 158444 191100
rect 158496 191088 158502 191140
rect 160370 191088 160376 191140
rect 160428 191128 160434 191140
rect 161290 191128 161296 191140
rect 160428 191100 161296 191128
rect 160428 191088 160434 191100
rect 161290 191088 161296 191100
rect 161348 191088 161354 191140
rect 161658 191088 161664 191140
rect 161716 191128 161722 191140
rect 162578 191128 162584 191140
rect 161716 191100 162584 191128
rect 161716 191088 161722 191100
rect 162578 191088 162584 191100
rect 162636 191088 162642 191140
rect 170674 191088 170680 191140
rect 170732 191128 170738 191140
rect 171502 191128 171508 191140
rect 170732 191100 171508 191128
rect 170732 191088 170738 191100
rect 171502 191088 171508 191100
rect 171560 191088 171566 191140
rect 174262 191088 174268 191140
rect 174320 191128 174326 191140
rect 174722 191128 174728 191140
rect 174320 191100 174728 191128
rect 174320 191088 174326 191100
rect 174722 191088 174728 191100
rect 174780 191088 174786 191140
rect 160186 191020 160192 191072
rect 160244 191060 160250 191072
rect 160922 191060 160928 191072
rect 160244 191032 160928 191060
rect 160244 191020 160250 191032
rect 160922 191020 160928 191032
rect 160980 191020 160986 191072
rect 171962 191020 171968 191072
rect 172020 191060 172026 191072
rect 172698 191060 172704 191072
rect 172020 191032 172704 191060
rect 172020 191020 172026 191032
rect 172698 191020 172704 191032
rect 172756 191020 172762 191072
rect 160094 190952 160100 191004
rect 160152 190992 160158 191004
rect 161014 190992 161020 191004
rect 160152 190964 161020 190992
rect 160152 190952 160158 190964
rect 161014 190952 161020 190964
rect 161072 190952 161078 191004
rect 145650 190816 145656 190868
rect 145708 190856 145714 190868
rect 151906 190856 151912 190868
rect 145708 190828 151912 190856
rect 145708 190816 145714 190828
rect 151906 190816 151912 190828
rect 151964 190816 151970 190868
rect 151906 190680 151912 190732
rect 151964 190720 151970 190732
rect 152642 190720 152648 190732
rect 151964 190692 152648 190720
rect 151964 190680 151970 190692
rect 152642 190680 152648 190692
rect 152700 190680 152706 190732
rect 141418 190544 141424 190596
rect 141476 190584 141482 190596
rect 143810 190584 143816 190596
rect 141476 190556 143816 190584
rect 141476 190544 141482 190556
rect 143810 190544 143816 190556
rect 143868 190544 143874 190596
rect 173894 190544 173900 190596
rect 173952 190584 173958 190596
rect 174170 190584 174176 190596
rect 173952 190556 174176 190584
rect 173952 190544 173958 190556
rect 174170 190544 174176 190556
rect 174228 190544 174234 190596
rect 113818 190408 113824 190460
rect 113876 190448 113882 190460
rect 141878 190448 141884 190460
rect 113876 190420 141884 190448
rect 113876 190408 113882 190420
rect 141878 190408 141884 190420
rect 141936 190408 141942 190460
rect 174170 190408 174176 190460
rect 174228 190448 174234 190460
rect 174538 190448 174544 190460
rect 174228 190420 174544 190448
rect 174228 190408 174234 190420
rect 174538 190408 174544 190420
rect 174596 190408 174602 190460
rect 110966 190340 110972 190392
rect 111024 190380 111030 190392
rect 138658 190380 138664 190392
rect 111024 190352 138664 190380
rect 111024 190340 111030 190352
rect 138658 190340 138664 190352
rect 138716 190340 138722 190392
rect 109954 190272 109960 190324
rect 110012 190312 110018 190324
rect 139946 190312 139952 190324
rect 110012 190284 139952 190312
rect 110012 190272 110018 190284
rect 139946 190272 139952 190284
rect 140004 190272 140010 190324
rect 112346 190204 112352 190256
rect 112404 190244 112410 190256
rect 141234 190244 141240 190256
rect 112404 190216 141240 190244
rect 112404 190204 112410 190216
rect 141234 190204 141240 190216
rect 141292 190204 141298 190256
rect 157242 190204 157248 190256
rect 157300 190244 157306 190256
rect 158806 190244 158812 190256
rect 157300 190216 158812 190244
rect 157300 190204 157306 190216
rect 158806 190204 158812 190216
rect 158864 190204 158870 190256
rect 107562 190136 107568 190188
rect 107620 190176 107626 190188
rect 140222 190176 140228 190188
rect 107620 190148 140228 190176
rect 107620 190136 107626 190148
rect 140222 190136 140228 190148
rect 140280 190136 140286 190188
rect 101766 190068 101772 190120
rect 101824 190108 101830 190120
rect 134058 190108 134064 190120
rect 101824 190080 134064 190108
rect 101824 190068 101830 190080
rect 134058 190068 134064 190080
rect 134116 190068 134122 190120
rect 101858 190000 101864 190052
rect 101916 190040 101922 190052
rect 134794 190040 134800 190052
rect 101916 190012 134800 190040
rect 101916 190000 101922 190012
rect 134794 190000 134800 190012
rect 134852 190000 134858 190052
rect 102962 189932 102968 189984
rect 103020 189972 103026 189984
rect 136174 189972 136180 189984
rect 103020 189944 136180 189972
rect 103020 189932 103026 189944
rect 136174 189932 136180 189944
rect 136232 189932 136238 189984
rect 101582 189864 101588 189916
rect 101640 189904 101646 189916
rect 134978 189904 134984 189916
rect 101640 189876 134984 189904
rect 101640 189864 101646 189876
rect 134978 189864 134984 189876
rect 135036 189864 135042 189916
rect 150986 189864 150992 189916
rect 151044 189904 151050 189916
rect 151630 189904 151636 189916
rect 151044 189876 151636 189904
rect 151044 189864 151050 189876
rect 151630 189864 151636 189876
rect 151688 189864 151694 189916
rect 102042 189796 102048 189848
rect 102100 189836 102106 189848
rect 135898 189836 135904 189848
rect 102100 189808 135904 189836
rect 102100 189796 102106 189808
rect 135898 189796 135904 189808
rect 135956 189796 135962 189848
rect 101950 189728 101956 189780
rect 102008 189768 102014 189780
rect 135254 189768 135260 189780
rect 102008 189740 135260 189768
rect 102008 189728 102014 189740
rect 135254 189728 135260 189740
rect 135312 189728 135318 189780
rect 134150 189660 134156 189712
rect 134208 189700 134214 189712
rect 134426 189700 134432 189712
rect 134208 189672 134432 189700
rect 134208 189660 134214 189672
rect 134426 189660 134432 189672
rect 134484 189660 134490 189712
rect 162854 189660 162860 189712
rect 162912 189700 162918 189712
rect 163222 189700 163228 189712
rect 162912 189672 163228 189700
rect 162912 189660 162918 189672
rect 163222 189660 163228 189672
rect 163280 189660 163286 189712
rect 126422 189456 126428 189508
rect 126480 189496 126486 189508
rect 149698 189496 149704 189508
rect 126480 189468 149704 189496
rect 126480 189456 126486 189468
rect 149698 189456 149704 189468
rect 149756 189456 149762 189508
rect 149698 189320 149704 189372
rect 149756 189360 149762 189372
rect 153194 189360 153200 189372
rect 149756 189332 153200 189360
rect 149756 189320 149762 189332
rect 153194 189320 153200 189332
rect 153252 189320 153258 189372
rect 162854 189320 162860 189372
rect 162912 189360 162918 189372
rect 163958 189360 163964 189372
rect 162912 189332 163964 189360
rect 162912 189320 162918 189332
rect 163958 189320 163964 189332
rect 164016 189320 164022 189372
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 120626 189020 120632 189032
rect 3476 188992 120632 189020
rect 3476 188980 3482 188992
rect 120626 188980 120632 188992
rect 120684 188980 120690 189032
rect 169754 188980 169760 189032
rect 169812 189020 169818 189032
rect 170950 189020 170956 189032
rect 169812 188992 170956 189020
rect 169812 188980 169818 188992
rect 170950 188980 170956 188992
rect 171008 188980 171014 189032
rect 132862 188912 132868 188964
rect 132920 188952 132926 188964
rect 133414 188952 133420 188964
rect 132920 188924 133420 188952
rect 132920 188912 132926 188924
rect 133414 188912 133420 188924
rect 133472 188912 133478 188964
rect 171410 188912 171416 188964
rect 171468 188952 171474 188964
rect 171594 188952 171600 188964
rect 171468 188924 171600 188952
rect 171468 188912 171474 188924
rect 171594 188912 171600 188924
rect 171652 188912 171658 188964
rect 154758 188776 154764 188828
rect 154816 188816 154822 188828
rect 155494 188816 155500 188828
rect 154816 188788 155500 188816
rect 154816 188776 154822 188788
rect 155494 188776 155500 188788
rect 155552 188776 155558 188828
rect 169938 188640 169944 188692
rect 169996 188680 170002 188692
rect 170582 188680 170588 188692
rect 169996 188652 170588 188680
rect 169996 188640 170002 188652
rect 170582 188640 170588 188652
rect 170640 188640 170646 188692
rect 131758 188436 131764 188488
rect 131816 188476 131822 188488
rect 139394 188476 139400 188488
rect 131816 188448 139400 188476
rect 131816 188436 131822 188448
rect 139394 188436 139400 188448
rect 139452 188436 139458 188488
rect 125502 188368 125508 188420
rect 125560 188408 125566 188420
rect 143534 188408 143540 188420
rect 125560 188380 143540 188408
rect 125560 188368 125566 188380
rect 143534 188368 143540 188380
rect 143592 188368 143598 188420
rect 176838 188368 176844 188420
rect 176896 188408 176902 188420
rect 177942 188408 177948 188420
rect 176896 188380 177948 188408
rect 176896 188368 176902 188380
rect 177942 188368 177948 188380
rect 178000 188368 178006 188420
rect 130378 188300 130384 188352
rect 130436 188340 130442 188352
rect 139302 188340 139308 188352
rect 130436 188312 139308 188340
rect 130436 188300 130442 188312
rect 139302 188300 139308 188312
rect 139360 188300 139366 188352
rect 176746 188300 176752 188352
rect 176804 188340 176810 188352
rect 177758 188340 177764 188352
rect 176804 188312 177764 188340
rect 176804 188300 176810 188312
rect 177758 188300 177764 188312
rect 177816 188300 177822 188352
rect 135622 188232 135628 188284
rect 135680 188272 135686 188284
rect 136266 188272 136272 188284
rect 135680 188244 136272 188272
rect 135680 188232 135686 188244
rect 136266 188232 136272 188244
rect 136324 188232 136330 188284
rect 176654 187892 176660 187944
rect 176712 187932 176718 187944
rect 178126 187932 178132 187944
rect 176712 187904 178132 187932
rect 176712 187892 176718 187904
rect 178126 187892 178132 187904
rect 178184 187892 178190 187944
rect 132678 187484 132684 187536
rect 132736 187524 132742 187536
rect 133874 187524 133880 187536
rect 132736 187496 133880 187524
rect 132736 187484 132742 187496
rect 133874 187484 133880 187496
rect 133932 187484 133938 187536
rect 126238 187416 126244 187468
rect 126296 187456 126302 187468
rect 150066 187456 150072 187468
rect 126296 187428 150072 187456
rect 126296 187416 126302 187428
rect 150066 187416 150072 187428
rect 150124 187416 150130 187468
rect 149514 186328 149520 186380
rect 149572 186368 149578 186380
rect 150158 186368 150164 186380
rect 149572 186340 150164 186368
rect 149572 186328 149578 186340
rect 150158 186328 150164 186340
rect 150216 186328 150222 186380
rect 148686 185784 148692 185836
rect 148744 185824 148750 185836
rect 154574 185824 154580 185836
rect 148744 185796 154580 185824
rect 148744 185784 148750 185796
rect 154574 185784 154580 185796
rect 154632 185784 154638 185836
rect 141142 185444 141148 185496
rect 141200 185484 141206 185496
rect 142062 185484 142068 185496
rect 141200 185456 142068 185484
rect 141200 185444 141206 185456
rect 142062 185444 142068 185456
rect 142120 185444 142126 185496
rect 161474 185104 161480 185156
rect 161532 185144 161538 185156
rect 162118 185144 162124 185156
rect 161532 185116 162124 185144
rect 161532 185104 161538 185116
rect 162118 185104 162124 185116
rect 162176 185104 162182 185156
rect 145742 184968 145748 185020
rect 145800 185008 145806 185020
rect 156506 185008 156512 185020
rect 145800 184980 156512 185008
rect 145800 184968 145806 184980
rect 156506 184968 156512 184980
rect 156564 184968 156570 185020
rect 175274 184968 175280 185020
rect 175332 185008 175338 185020
rect 176102 185008 176108 185020
rect 175332 184980 176108 185008
rect 175332 184968 175338 184980
rect 176102 184968 176108 184980
rect 176160 184968 176166 185020
rect 153470 184696 153476 184748
rect 153528 184736 153534 184748
rect 154298 184736 154304 184748
rect 153528 184708 154304 184736
rect 153528 184696 153534 184708
rect 154298 184696 154304 184708
rect 154356 184696 154362 184748
rect 175550 184696 175556 184748
rect 175608 184736 175614 184748
rect 175918 184736 175924 184748
rect 175608 184708 175924 184736
rect 175608 184696 175614 184708
rect 175918 184696 175924 184708
rect 175976 184696 175982 184748
rect 159266 184016 159272 184068
rect 159324 184056 159330 184068
rect 160002 184056 160008 184068
rect 159324 184028 160008 184056
rect 159324 184016 159330 184028
rect 160002 184016 160008 184028
rect 160060 184016 160066 184068
rect 172606 183472 172612 183524
rect 172664 183512 172670 183524
rect 172882 183512 172888 183524
rect 172664 183484 172888 183512
rect 172664 183472 172670 183484
rect 172882 183472 172888 183484
rect 172940 183472 172946 183524
rect 164326 183336 164332 183388
rect 164384 183376 164390 183388
rect 165338 183376 165344 183388
rect 164384 183348 165344 183376
rect 164384 183336 164390 183348
rect 165338 183336 165344 183348
rect 165396 183336 165402 183388
rect 129090 183064 129096 183116
rect 129148 183104 129154 183116
rect 137370 183104 137376 183116
rect 129148 183076 137376 183104
rect 129148 183064 129154 183076
rect 137370 183064 137376 183076
rect 137428 183064 137434 183116
rect 127618 181976 127624 182028
rect 127676 182016 127682 182028
rect 141602 182016 141608 182028
rect 127676 181988 141608 182016
rect 127676 181976 127682 181988
rect 141602 181976 141608 181988
rect 141660 181976 141666 182028
rect 171134 181432 171140 181484
rect 171192 181472 171198 181484
rect 171318 181472 171324 181484
rect 171192 181444 171324 181472
rect 171192 181432 171198 181444
rect 171318 181432 171324 181444
rect 171376 181432 171382 181484
rect 129274 180276 129280 180328
rect 129332 180316 129338 180328
rect 149882 180316 149888 180328
rect 129332 180288 149888 180316
rect 129332 180276 129338 180288
rect 149882 180276 149888 180288
rect 149940 180276 149946 180328
rect 145834 179120 145840 179172
rect 145892 179160 145898 179172
rect 146570 179160 146576 179172
rect 145892 179132 146576 179160
rect 145892 179120 145898 179132
rect 146570 179120 146576 179132
rect 146628 179120 146634 179172
rect 188614 178032 188620 178084
rect 188672 178072 188678 178084
rect 580166 178072 580172 178084
rect 188672 178044 580172 178072
rect 188672 178032 188678 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 189810 165588 189816 165640
rect 189868 165628 189874 165640
rect 580166 165628 580172 165640
rect 189868 165600 580172 165628
rect 189868 165588 189874 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 168650 155320 168656 155372
rect 168708 155360 168714 155372
rect 203426 155360 203432 155372
rect 168708 155332 203432 155360
rect 168708 155320 168714 155332
rect 203426 155320 203432 155332
rect 203484 155320 203490 155372
rect 169570 155252 169576 155304
rect 169628 155292 169634 155304
rect 203518 155292 203524 155304
rect 169628 155264 203524 155292
rect 169628 155252 169634 155264
rect 203518 155252 203524 155264
rect 203576 155252 203582 155304
rect 167270 155184 167276 155236
rect 167328 155224 167334 155236
rect 202322 155224 202328 155236
rect 167328 155196 202328 155224
rect 167328 155184 167334 155196
rect 202322 155184 202328 155196
rect 202380 155184 202386 155236
rect 163130 153144 163136 153196
rect 163188 153184 163194 153196
rect 185946 153184 185952 153196
rect 163188 153156 185952 153184
rect 163188 153144 163194 153156
rect 185946 153144 185952 153156
rect 186004 153144 186010 153196
rect 161750 153076 161756 153128
rect 161808 153116 161814 153128
rect 185578 153116 185584 153128
rect 161808 153088 185584 153116
rect 161808 153076 161814 153088
rect 185578 153076 185584 153088
rect 185636 153076 185642 153128
rect 160278 153008 160284 153060
rect 160336 153048 160342 153060
rect 184290 153048 184296 153060
rect 160336 153020 184296 153048
rect 160336 153008 160342 153020
rect 184290 153008 184296 153020
rect 184348 153008 184354 153060
rect 161842 152940 161848 152992
rect 161900 152980 161906 152992
rect 186038 152980 186044 152992
rect 161900 152952 186044 152980
rect 161900 152940 161906 152952
rect 186038 152940 186044 152952
rect 186096 152940 186102 152992
rect 160462 152872 160468 152924
rect 160520 152912 160526 152924
rect 185670 152912 185676 152924
rect 160520 152884 185676 152912
rect 160520 152872 160526 152884
rect 185670 152872 185676 152884
rect 185728 152872 185734 152924
rect 158990 152804 158996 152856
rect 159048 152844 159054 152856
rect 184382 152844 184388 152856
rect 159048 152816 184388 152844
rect 159048 152804 159054 152816
rect 184382 152804 184388 152816
rect 184440 152804 184446 152856
rect 160370 152736 160376 152788
rect 160428 152776 160434 152788
rect 186130 152776 186136 152788
rect 160428 152748 186136 152776
rect 160428 152736 160434 152748
rect 186130 152736 186136 152748
rect 186188 152736 186194 152788
rect 160002 152668 160008 152720
rect 160060 152708 160066 152720
rect 184750 152708 184756 152720
rect 160060 152680 184756 152708
rect 160060 152668 160066 152680
rect 184750 152668 184756 152680
rect 184808 152668 184814 152720
rect 167086 152600 167092 152652
rect 167144 152640 167150 152652
rect 199194 152640 199200 152652
rect 167144 152612 199200 152640
rect 167144 152600 167150 152612
rect 199194 152600 199200 152612
rect 199252 152600 199258 152652
rect 164602 152532 164608 152584
rect 164660 152572 164666 152584
rect 199286 152572 199292 152584
rect 164660 152544 199292 152572
rect 164660 152532 164666 152544
rect 199286 152532 199292 152544
rect 199344 152532 199350 152584
rect 165706 152464 165712 152516
rect 165764 152504 165770 152516
rect 200850 152504 200856 152516
rect 165764 152476 200856 152504
rect 165764 152464 165770 152476
rect 200850 152464 200856 152476
rect 200908 152464 200914 152516
rect 163222 152396 163228 152448
rect 163280 152436 163286 152448
rect 185854 152436 185860 152448
rect 163280 152408 185860 152436
rect 163280 152396 163286 152408
rect 185854 152396 185860 152408
rect 185912 152396 185918 152448
rect 165798 152328 165804 152380
rect 165856 152368 165862 152380
rect 184566 152368 184572 152380
rect 165856 152340 184572 152368
rect 165856 152328 165862 152340
rect 184566 152328 184572 152340
rect 184624 152328 184630 152380
rect 168374 152260 168380 152312
rect 168432 152300 168438 152312
rect 183186 152300 183192 152312
rect 168432 152272 183192 152300
rect 168432 152260 168438 152272
rect 183186 152260 183192 152272
rect 183244 152260 183250 152312
rect 100202 151172 100208 151224
rect 100260 151212 100266 151224
rect 132678 151212 132684 151224
rect 100260 151184 132684 151212
rect 100260 151172 100266 151184
rect 132678 151172 132684 151184
rect 132736 151172 132742 151224
rect 100294 151104 100300 151156
rect 100352 151144 100358 151156
rect 134242 151144 134248 151156
rect 100352 151116 134248 151144
rect 100352 151104 100358 151116
rect 134242 151104 134248 151116
rect 134300 151104 134306 151156
rect 100386 151036 100392 151088
rect 100444 151076 100450 151088
rect 134426 151076 134432 151088
rect 100444 151048 134432 151076
rect 100444 151036 100450 151048
rect 134426 151036 134432 151048
rect 134484 151036 134490 151088
rect 176930 150356 176936 150408
rect 176988 150396 176994 150408
rect 202782 150396 202788 150408
rect 176988 150368 202788 150396
rect 176988 150356 176994 150368
rect 202782 150356 202788 150368
rect 202840 150356 202846 150408
rect 176838 150288 176844 150340
rect 176896 150328 176902 150340
rect 201402 150328 201408 150340
rect 176896 150300 201408 150328
rect 176896 150288 176902 150300
rect 201402 150288 201408 150300
rect 201460 150288 201466 150340
rect 184198 150220 184204 150272
rect 184256 150260 184262 150272
rect 202230 150260 202236 150272
rect 184256 150232 202236 150260
rect 184256 150220 184262 150232
rect 202230 150220 202236 150232
rect 202288 150220 202294 150272
rect 175550 150152 175556 150204
rect 175608 150192 175614 150204
rect 204530 150192 204536 150204
rect 175608 150164 204536 150192
rect 175608 150152 175614 150164
rect 204530 150152 204536 150164
rect 204588 150152 204594 150204
rect 175458 150084 175464 150136
rect 175516 150124 175522 150136
rect 204622 150124 204628 150136
rect 175516 150096 204628 150124
rect 175516 150084 175522 150096
rect 204622 150084 204628 150096
rect 204680 150084 204686 150136
rect 174354 150016 174360 150068
rect 174412 150056 174418 150068
rect 203702 150056 203708 150068
rect 174412 150028 203708 150056
rect 174412 150016 174418 150028
rect 203702 150016 203708 150028
rect 203760 150016 203766 150068
rect 174170 149948 174176 150000
rect 174228 149988 174234 150000
rect 203610 149988 203616 150000
rect 174228 149960 203616 149988
rect 174228 149948 174234 149960
rect 203610 149948 203616 149960
rect 203668 149948 203674 150000
rect 175642 149880 175648 149932
rect 175700 149920 175706 149932
rect 206186 149920 206192 149932
rect 175700 149892 206192 149920
rect 175700 149880 175706 149892
rect 206186 149880 206192 149892
rect 206244 149880 206250 149932
rect 175274 149812 175280 149864
rect 175332 149852 175338 149864
rect 206278 149852 206284 149864
rect 175332 149824 206284 149852
rect 175332 149812 175338 149824
rect 206278 149812 206284 149824
rect 206336 149812 206342 149864
rect 175366 149744 175372 149796
rect 175424 149784 175430 149796
rect 206370 149784 206376 149796
rect 175424 149756 206376 149784
rect 175424 149744 175430 149756
rect 206370 149744 206376 149756
rect 206428 149744 206434 149796
rect 148962 149676 148968 149728
rect 149020 149716 149026 149728
rect 184658 149716 184664 149728
rect 149020 149688 184664 149716
rect 149020 149676 149026 149688
rect 184658 149676 184664 149688
rect 184716 149676 184722 149728
rect 3418 149064 3424 149116
rect 3476 149104 3482 149116
rect 9582 149104 9588 149116
rect 3476 149076 9588 149104
rect 3476 149064 3482 149076
rect 9582 149064 9588 149076
rect 9640 149064 9646 149116
rect 126606 148996 126612 149048
rect 126664 149036 126670 149048
rect 154850 149036 154856 149048
rect 126664 149008 154856 149036
rect 126664 148996 126670 149008
rect 154850 148996 154856 149008
rect 154908 148996 154914 149048
rect 113358 148928 113364 148980
rect 113416 148968 113422 148980
rect 142614 148968 142620 148980
rect 113416 148940 142620 148968
rect 113416 148928 113422 148940
rect 142614 148928 142620 148940
rect 142672 148928 142678 148980
rect 125042 148860 125048 148912
rect 125100 148900 125106 148912
rect 153470 148900 153476 148912
rect 125100 148872 153476 148900
rect 125100 148860 125106 148872
rect 153470 148860 153476 148872
rect 153528 148860 153534 148912
rect 123110 148792 123116 148844
rect 123168 148832 123174 148844
rect 152090 148832 152096 148844
rect 123168 148804 152096 148832
rect 123168 148792 123174 148804
rect 152090 148792 152096 148804
rect 152148 148792 152154 148844
rect 102686 148724 102692 148776
rect 102744 148764 102750 148776
rect 131850 148764 131856 148776
rect 102744 148736 131856 148764
rect 102744 148724 102750 148736
rect 131850 148724 131856 148736
rect 131908 148724 131914 148776
rect 178678 148724 178684 148776
rect 178736 148764 178742 148776
rect 195514 148764 195520 148776
rect 178736 148736 195520 148764
rect 178736 148724 178742 148736
rect 195514 148724 195520 148736
rect 195572 148724 195578 148776
rect 124490 148656 124496 148708
rect 124548 148696 124554 148708
rect 156138 148696 156144 148708
rect 124548 148668 156144 148696
rect 124548 148656 124554 148668
rect 156138 148656 156144 148668
rect 156196 148656 156202 148708
rect 164418 148656 164424 148708
rect 164476 148696 164482 148708
rect 186958 148696 186964 148708
rect 164476 148668 186964 148696
rect 164476 148656 164482 148668
rect 186958 148656 186964 148668
rect 187016 148656 187022 148708
rect 104066 148588 104072 148640
rect 104124 148628 104130 148640
rect 135622 148628 135628 148640
rect 104124 148600 135628 148628
rect 104124 148588 104130 148600
rect 135622 148588 135628 148600
rect 135680 148588 135686 148640
rect 160186 148588 160192 148640
rect 160244 148628 160250 148640
rect 184106 148628 184112 148640
rect 160244 148600 184112 148628
rect 160244 148588 160250 148600
rect 184106 148588 184112 148600
rect 184164 148588 184170 148640
rect 120442 148520 120448 148572
rect 120500 148560 120506 148572
rect 153286 148560 153292 148572
rect 120500 148532 153292 148560
rect 120500 148520 120506 148532
rect 153286 148520 153292 148532
rect 153344 148520 153350 148572
rect 166994 148520 167000 148572
rect 167052 148560 167058 148572
rect 198274 148560 198280 148572
rect 167052 148532 198280 148560
rect 167052 148520 167058 148532
rect 198274 148520 198280 148532
rect 198332 148520 198338 148572
rect 117590 148452 117596 148504
rect 117648 148492 117654 148504
rect 152182 148492 152188 148504
rect 117648 148464 152188 148492
rect 117648 148452 117654 148464
rect 152182 148452 152188 148464
rect 152240 148452 152246 148504
rect 163038 148452 163044 148504
rect 163096 148492 163102 148504
rect 196986 148492 196992 148504
rect 163096 148464 196992 148492
rect 163096 148452 163102 148464
rect 196986 148452 196992 148464
rect 197044 148452 197050 148504
rect 116210 148384 116216 148436
rect 116268 148424 116274 148436
rect 151722 148424 151728 148436
rect 116268 148396 151728 148424
rect 116268 148384 116274 148396
rect 151722 148384 151728 148396
rect 151780 148384 151786 148436
rect 164510 148384 164516 148436
rect 164568 148424 164574 148436
rect 199470 148424 199476 148436
rect 164568 148396 199476 148424
rect 164568 148384 164574 148396
rect 199470 148384 199476 148396
rect 199528 148384 199534 148436
rect 9582 148316 9588 148368
rect 9640 148356 9646 148368
rect 180886 148356 180892 148368
rect 9640 148328 180892 148356
rect 9640 148316 9646 148328
rect 180886 148316 180892 148328
rect 180944 148356 180950 148368
rect 196710 148356 196716 148368
rect 180944 148328 196716 148356
rect 180944 148316 180950 148328
rect 196710 148316 196716 148328
rect 196768 148316 196774 148368
rect 113542 148248 113548 148300
rect 113600 148288 113606 148300
rect 142982 148288 142988 148300
rect 113600 148260 142988 148288
rect 113600 148248 113606 148260
rect 142982 148248 142988 148260
rect 143040 148248 143046 148300
rect 116118 148180 116124 148232
rect 116176 148220 116182 148232
rect 142522 148220 142528 148232
rect 116176 148192 142528 148220
rect 116176 148180 116182 148192
rect 142522 148180 142528 148192
rect 142580 148180 142586 148232
rect 126514 148112 126520 148164
rect 126572 148152 126578 148164
rect 148318 148152 148324 148164
rect 126572 148124 148324 148152
rect 126572 148112 126578 148124
rect 148318 148112 148324 148124
rect 148376 148112 148382 148164
rect 178218 147568 178224 147620
rect 178276 147608 178282 147620
rect 196526 147608 196532 147620
rect 178276 147580 196532 147608
rect 178276 147568 178282 147580
rect 196526 147568 196532 147580
rect 196584 147568 196590 147620
rect 178034 147500 178040 147552
rect 178092 147540 178098 147552
rect 198090 147540 198096 147552
rect 178092 147512 198096 147540
rect 178092 147500 178098 147512
rect 198090 147500 198096 147512
rect 198148 147500 198154 147552
rect 171226 147432 171232 147484
rect 171284 147472 171290 147484
rect 194318 147472 194324 147484
rect 171284 147444 194324 147472
rect 171284 147432 171290 147444
rect 194318 147432 194324 147444
rect 194376 147432 194382 147484
rect 172790 147364 172796 147416
rect 172848 147404 172854 147416
rect 195330 147404 195336 147416
rect 172848 147376 195336 147404
rect 172848 147364 172854 147376
rect 195330 147364 195336 147376
rect 195388 147364 195394 147416
rect 172882 147296 172888 147348
rect 172940 147336 172946 147348
rect 196526 147336 196532 147348
rect 172940 147308 196532 147336
rect 172940 147296 172946 147308
rect 196526 147296 196532 147308
rect 196584 147296 196590 147348
rect 113910 147228 113916 147280
rect 113968 147268 113974 147280
rect 126974 147268 126980 147280
rect 113968 147240 126980 147268
rect 113968 147228 113974 147240
rect 126974 147228 126980 147240
rect 127032 147228 127038 147280
rect 170030 147228 170036 147280
rect 170088 147268 170094 147280
rect 193950 147268 193956 147280
rect 170088 147240 193956 147268
rect 170088 147228 170094 147240
rect 193950 147228 193956 147240
rect 194008 147228 194014 147280
rect 115014 147160 115020 147212
rect 115072 147200 115078 147212
rect 137278 147200 137284 147212
rect 115072 147172 137284 147200
rect 115072 147160 115078 147172
rect 137278 147160 137284 147172
rect 137336 147160 137342 147212
rect 171318 147160 171324 147212
rect 171376 147200 171382 147212
rect 195422 147200 195428 147212
rect 171376 147172 195428 147200
rect 171376 147160 171382 147172
rect 195422 147160 195428 147172
rect 195480 147160 195486 147212
rect 114922 147092 114928 147144
rect 114980 147132 114986 147144
rect 140958 147132 140964 147144
rect 114980 147104 140964 147132
rect 114980 147092 114986 147104
rect 140958 147092 140964 147104
rect 141016 147092 141022 147144
rect 172698 147092 172704 147144
rect 172756 147132 172762 147144
rect 198366 147132 198372 147144
rect 172756 147104 198372 147132
rect 172756 147092 172762 147104
rect 198366 147092 198372 147104
rect 198424 147092 198430 147144
rect 112254 147024 112260 147076
rect 112312 147064 112318 147076
rect 138474 147064 138480 147076
rect 112312 147036 138480 147064
rect 112312 147024 112318 147036
rect 138474 147024 138480 147036
rect 138532 147024 138538 147076
rect 171410 147024 171416 147076
rect 171468 147064 171474 147076
rect 196710 147064 196716 147076
rect 171468 147036 196716 147064
rect 171468 147024 171474 147036
rect 196710 147024 196716 147036
rect 196768 147024 196774 147076
rect 117498 146956 117504 147008
rect 117556 146996 117562 147008
rect 145650 146996 145656 147008
rect 117556 146968 145656 146996
rect 117556 146956 117562 146968
rect 145650 146956 145656 146968
rect 145708 146956 145714 147008
rect 171502 146956 171508 147008
rect 171560 146996 171566 147008
rect 198090 146996 198096 147008
rect 171560 146968 198096 146996
rect 171560 146956 171566 146968
rect 198090 146956 198096 146968
rect 198148 146956 198154 147008
rect 110874 146888 110880 146940
rect 110932 146928 110938 146940
rect 139762 146928 139768 146940
rect 110932 146900 139768 146928
rect 110932 146888 110938 146900
rect 139762 146888 139768 146900
rect 139820 146888 139826 146940
rect 173986 146888 173992 146940
rect 174044 146928 174050 146940
rect 206462 146928 206468 146940
rect 174044 146900 206468 146928
rect 174044 146888 174050 146900
rect 206462 146888 206468 146900
rect 206520 146888 206526 146940
rect 179598 146820 179604 146872
rect 179656 146860 179662 146872
rect 197906 146860 197912 146872
rect 179656 146832 197912 146860
rect 179656 146820 179662 146832
rect 197906 146820 197912 146832
rect 197964 146820 197970 146872
rect 178402 146752 178408 146804
rect 178460 146792 178466 146804
rect 195146 146792 195152 146804
rect 178460 146764 195152 146792
rect 178460 146752 178466 146764
rect 195146 146752 195152 146764
rect 195204 146752 195210 146804
rect 179690 146684 179696 146736
rect 179748 146724 179754 146736
rect 193766 146724 193772 146736
rect 179748 146696 193772 146724
rect 179748 146684 179754 146696
rect 193766 146684 193772 146696
rect 193824 146684 193830 146736
rect 116854 146208 116860 146260
rect 116912 146248 116918 146260
rect 131298 146248 131304 146260
rect 116912 146220 131304 146248
rect 116912 146208 116918 146220
rect 131298 146208 131304 146220
rect 131356 146208 131362 146260
rect 178310 146208 178316 146260
rect 178368 146248 178374 146260
rect 188246 146248 188252 146260
rect 178368 146220 188252 146248
rect 178368 146208 178374 146220
rect 188246 146208 188252 146220
rect 188304 146208 188310 146260
rect 116762 146140 116768 146192
rect 116820 146180 116826 146192
rect 131206 146180 131212 146192
rect 116820 146152 131212 146180
rect 116820 146140 116826 146152
rect 131206 146140 131212 146152
rect 131264 146140 131270 146192
rect 178126 146140 178132 146192
rect 178184 146180 178190 146192
rect 191282 146180 191288 146192
rect 178184 146152 191288 146180
rect 178184 146140 178190 146152
rect 191282 146140 191288 146152
rect 191340 146140 191346 146192
rect 121914 146072 121920 146124
rect 121972 146112 121978 146124
rect 146662 146112 146668 146124
rect 121972 146084 146668 146112
rect 121972 146072 121978 146084
rect 146662 146072 146668 146084
rect 146720 146072 146726 146124
rect 175550 146072 175556 146124
rect 175608 146112 175614 146124
rect 197814 146112 197820 146124
rect 175608 146084 197820 146112
rect 175608 146072 175614 146084
rect 197814 146072 197820 146084
rect 197872 146072 197878 146124
rect 121822 146004 121828 146056
rect 121880 146044 121886 146056
rect 149514 146044 149520 146056
rect 121880 146016 149520 146044
rect 121880 146004 121886 146016
rect 149514 146004 149520 146016
rect 149572 146004 149578 146056
rect 161566 146004 161572 146056
rect 161624 146044 161630 146056
rect 188338 146044 188344 146056
rect 161624 146016 188344 146044
rect 161624 146004 161630 146016
rect 188338 146004 188344 146016
rect 188396 146004 188402 146056
rect 118786 145936 118792 145988
rect 118844 145976 118850 145988
rect 146570 145976 146576 145988
rect 118844 145948 146576 145976
rect 118844 145936 118850 145948
rect 146570 145936 146576 145948
rect 146628 145936 146634 145988
rect 165614 145936 165620 145988
rect 165672 145976 165678 145988
rect 194134 145976 194140 145988
rect 165672 145948 194140 145976
rect 165672 145936 165678 145948
rect 194134 145936 194140 145948
rect 194192 145936 194198 145988
rect 118970 145868 118976 145920
rect 119028 145908 119034 145920
rect 146478 145908 146484 145920
rect 119028 145880 146484 145908
rect 119028 145868 119034 145880
rect 146478 145868 146484 145880
rect 146536 145868 146542 145920
rect 161474 145868 161480 145920
rect 161532 145908 161538 145920
rect 190086 145908 190092 145920
rect 161532 145880 190092 145908
rect 161532 145868 161538 145880
rect 190086 145868 190092 145880
rect 190144 145868 190150 145920
rect 119062 145800 119068 145852
rect 119120 145840 119126 145852
rect 147674 145840 147680 145852
rect 119120 145812 147680 145840
rect 119120 145800 119126 145812
rect 147674 145800 147680 145812
rect 147732 145800 147738 145852
rect 162946 145800 162952 145852
rect 163004 145840 163010 145852
rect 194226 145840 194232 145852
rect 163004 145812 194232 145840
rect 163004 145800 163010 145812
rect 194226 145800 194232 145812
rect 194284 145800 194290 145852
rect 120350 145732 120356 145784
rect 120408 145772 120414 145784
rect 153102 145772 153108 145784
rect 120408 145744 153108 145772
rect 120408 145732 120414 145744
rect 153102 145732 153108 145744
rect 153160 145732 153166 145784
rect 160094 145732 160100 145784
rect 160152 145772 160158 145784
rect 195146 145772 195152 145784
rect 160152 145744 195152 145772
rect 160152 145732 160158 145744
rect 195146 145732 195152 145744
rect 195204 145732 195210 145784
rect 116394 145664 116400 145716
rect 116452 145704 116458 145716
rect 150618 145704 150624 145716
rect 116452 145676 150624 145704
rect 116452 145664 116458 145676
rect 150618 145664 150624 145676
rect 150676 145664 150682 145716
rect 159910 145664 159916 145716
rect 159968 145704 159974 145716
rect 191374 145704 191380 145716
rect 159968 145676 191380 145704
rect 159968 145664 159974 145676
rect 191374 145664 191380 145676
rect 191432 145664 191438 145716
rect 119982 145596 119988 145648
rect 120040 145636 120046 145648
rect 160094 145636 160100 145648
rect 120040 145608 160100 145636
rect 120040 145596 120046 145608
rect 160094 145596 160100 145608
rect 160152 145596 160158 145648
rect 161658 145596 161664 145648
rect 161716 145636 161722 145648
rect 192938 145636 192944 145648
rect 161716 145608 192944 145636
rect 161716 145596 161722 145608
rect 192938 145596 192944 145608
rect 192996 145596 193002 145648
rect 3510 145528 3516 145580
rect 3568 145568 3574 145580
rect 179782 145568 179788 145580
rect 3568 145540 179788 145568
rect 3568 145528 3574 145540
rect 179782 145528 179788 145540
rect 179840 145568 179846 145580
rect 189626 145568 189632 145580
rect 179840 145540 189632 145568
rect 179840 145528 179846 145540
rect 189626 145528 189632 145540
rect 189684 145528 189690 145580
rect 116762 145460 116768 145512
rect 116820 145500 116826 145512
rect 130562 145500 130568 145512
rect 116820 145472 130568 145500
rect 116820 145460 116826 145472
rect 130562 145460 130568 145472
rect 130620 145460 130626 145512
rect 180426 145460 180432 145512
rect 180484 145500 180490 145512
rect 190178 145500 190184 145512
rect 180484 145472 190184 145500
rect 180484 145460 180490 145472
rect 190178 145460 190184 145472
rect 190236 145460 190242 145512
rect 116946 145392 116952 145444
rect 117004 145432 117010 145444
rect 129734 145432 129740 145444
rect 117004 145404 129740 145432
rect 117004 145392 117010 145404
rect 129734 145392 129740 145404
rect 129792 145392 129798 145444
rect 180334 145392 180340 145444
rect 180392 145432 180398 145444
rect 189994 145432 190000 145444
rect 180392 145404 190000 145432
rect 180392 145392 180398 145404
rect 189994 145392 190000 145404
rect 190052 145392 190058 145444
rect 179414 145324 179420 145376
rect 179472 145364 179478 145376
rect 189718 145364 189724 145376
rect 179472 145336 189724 145364
rect 179472 145324 179478 145336
rect 189718 145324 189724 145336
rect 189776 145324 189782 145376
rect 183002 144848 183008 144900
rect 183060 144888 183066 144900
rect 192754 144888 192760 144900
rect 183060 144860 192760 144888
rect 183060 144848 183066 144860
rect 192754 144848 192760 144860
rect 192812 144848 192818 144900
rect 179506 144780 179512 144832
rect 179564 144820 179570 144832
rect 193582 144820 193588 144832
rect 179564 144792 193588 144820
rect 179564 144780 179570 144792
rect 193582 144780 193588 144792
rect 193640 144780 193646 144832
rect 118050 144712 118056 144764
rect 118108 144752 118114 144764
rect 130010 144752 130016 144764
rect 118108 144724 130016 144752
rect 118108 144712 118114 144724
rect 130010 144712 130016 144724
rect 130068 144712 130074 144764
rect 173802 144712 173808 144764
rect 173860 144752 173866 144764
rect 190914 144752 190920 144764
rect 173860 144724 190920 144752
rect 173860 144712 173866 144724
rect 190914 144712 190920 144724
rect 190972 144712 190978 144764
rect 119706 144644 119712 144696
rect 119764 144684 119770 144696
rect 138106 144684 138112 144696
rect 119764 144656 138112 144684
rect 119764 144644 119770 144656
rect 138106 144644 138112 144656
rect 138164 144644 138170 144696
rect 170766 144644 170772 144696
rect 170824 144684 170830 144696
rect 192018 144684 192024 144696
rect 170824 144656 192024 144684
rect 170824 144644 170830 144656
rect 192018 144644 192024 144656
rect 192076 144644 192082 144696
rect 116486 144576 116492 144628
rect 116544 144616 116550 144628
rect 143810 144616 143816 144628
rect 116544 144588 143816 144616
rect 116544 144576 116550 144588
rect 143810 144576 143816 144588
rect 143868 144576 143874 144628
rect 172422 144576 172428 144628
rect 172480 144616 172486 144628
rect 194962 144616 194968 144628
rect 172480 144588 194968 144616
rect 172480 144576 172486 144588
rect 194962 144576 194968 144588
rect 195020 144576 195026 144628
rect 122374 144508 122380 144560
rect 122432 144548 122438 144560
rect 152642 144548 152648 144560
rect 122432 144520 152648 144548
rect 122432 144508 122438 144520
rect 152642 144508 152648 144520
rect 152700 144508 152706 144560
rect 169110 144508 169116 144560
rect 169168 144548 169174 144560
rect 192386 144548 192392 144560
rect 169168 144520 192392 144548
rect 169168 144508 169174 144520
rect 192386 144508 192392 144520
rect 192444 144508 192450 144560
rect 122558 144440 122564 144492
rect 122616 144480 122622 144492
rect 153838 144480 153844 144492
rect 122616 144452 153844 144480
rect 122616 144440 122622 144452
rect 153838 144440 153844 144452
rect 153896 144440 153902 144492
rect 158162 144440 158168 144492
rect 158220 144480 158226 144492
rect 192846 144480 192852 144492
rect 158220 144452 192852 144480
rect 158220 144440 158226 144452
rect 192846 144440 192852 144452
rect 192904 144440 192910 144492
rect 119706 144372 119712 144424
rect 119764 144412 119770 144424
rect 150526 144412 150532 144424
rect 119764 144384 150532 144412
rect 119764 144372 119770 144384
rect 150526 144372 150532 144384
rect 150584 144372 150590 144424
rect 152550 144372 152556 144424
rect 152608 144412 152614 144424
rect 186406 144412 186412 144424
rect 152608 144384 186412 144412
rect 152608 144372 152614 144384
rect 186406 144372 186412 144384
rect 186464 144372 186470 144424
rect 116854 144304 116860 144356
rect 116912 144344 116918 144356
rect 148594 144344 148600 144356
rect 116912 144316 148600 144344
rect 116912 144304 116918 144316
rect 148594 144304 148600 144316
rect 148652 144304 148658 144356
rect 156414 144304 156420 144356
rect 156472 144344 156478 144356
rect 191006 144344 191012 144356
rect 156472 144316 191012 144344
rect 156472 144304 156478 144316
rect 191006 144304 191012 144316
rect 191064 144304 191070 144356
rect 115290 144236 115296 144288
rect 115348 144276 115354 144288
rect 131390 144276 131396 144288
rect 115348 144248 131396 144276
rect 115348 144236 115354 144248
rect 131390 144236 131396 144248
rect 131448 144276 131454 144288
rect 188614 144276 188620 144288
rect 131448 144248 188620 144276
rect 131448 144236 131454 144248
rect 188614 144236 188620 144248
rect 188672 144236 188678 144288
rect 116670 144168 116676 144220
rect 116728 144208 116734 144220
rect 129366 144208 129372 144220
rect 116728 144180 129372 144208
rect 116728 144168 116734 144180
rect 129366 144168 129372 144180
rect 129424 144168 129430 144220
rect 130010 144168 130016 144220
rect 130068 144208 130074 144220
rect 189810 144208 189816 144220
rect 130068 144180 189816 144208
rect 130068 144168 130074 144180
rect 189810 144168 189816 144180
rect 189868 144168 189874 144220
rect 188154 143896 188160 143948
rect 188212 143896 188218 143948
rect 188172 143676 188200 143896
rect 188154 143624 188160 143676
rect 188212 143624 188218 143676
rect 119982 143556 119988 143608
rect 120040 143596 120046 143608
rect 145282 143596 145288 143608
rect 120040 143568 145288 143596
rect 120040 143556 120046 143568
rect 145282 143556 145288 143568
rect 145340 143556 145346 143608
rect 187878 143556 187884 143608
rect 187936 143596 187942 143608
rect 188062 143596 188068 143608
rect 187936 143568 188068 143596
rect 187936 143556 187942 143568
rect 188062 143556 188068 143568
rect 188120 143556 188126 143608
rect 113726 143488 113732 143540
rect 113784 143528 113790 143540
rect 123846 143528 123852 143540
rect 113784 143500 123852 143528
rect 113784 143488 113790 143500
rect 123846 143488 123852 143500
rect 123904 143488 123910 143540
rect 124030 143488 124036 143540
rect 124088 143528 124094 143540
rect 124582 143528 124588 143540
rect 124088 143500 124588 143528
rect 124088 143488 124094 143500
rect 124582 143488 124588 143500
rect 124640 143488 124646 143540
rect 131482 143528 131488 143540
rect 125888 143500 131488 143528
rect 119798 143420 119804 143472
rect 119856 143460 119862 143472
rect 125888 143460 125916 143500
rect 131482 143488 131488 143500
rect 131540 143488 131546 143540
rect 131574 143488 131580 143540
rect 131632 143528 131638 143540
rect 580350 143528 580356 143540
rect 131632 143500 580356 143528
rect 131632 143488 131638 143500
rect 580350 143488 580356 143500
rect 580408 143488 580414 143540
rect 119856 143432 125916 143460
rect 119856 143420 119862 143432
rect 131114 143420 131120 143472
rect 131172 143460 131178 143472
rect 137554 143460 137560 143472
rect 131172 143432 137560 143460
rect 131172 143420 131178 143432
rect 137554 143420 137560 143432
rect 137612 143420 137618 143472
rect 146294 143420 146300 143472
rect 146352 143460 146358 143472
rect 149146 143460 149152 143472
rect 146352 143432 149152 143460
rect 146352 143420 146358 143432
rect 149146 143420 149152 143432
rect 149204 143420 149210 143472
rect 175458 143420 175464 143472
rect 175516 143460 175522 143472
rect 179506 143460 179512 143472
rect 175516 143432 179512 143460
rect 175516 143420 175522 143432
rect 179506 143420 179512 143432
rect 179564 143420 179570 143472
rect 181530 143420 181536 143472
rect 181588 143460 181594 143472
rect 187050 143460 187056 143472
rect 181588 143432 187056 143460
rect 181588 143420 181594 143432
rect 187050 143420 187056 143432
rect 187108 143420 187114 143472
rect 187418 143420 187424 143472
rect 187476 143460 187482 143472
rect 187878 143460 187884 143472
rect 187476 143432 187884 143460
rect 187476 143420 187482 143432
rect 187878 143420 187884 143432
rect 187936 143420 187942 143472
rect 193674 143460 193680 143472
rect 187988 143432 193680 143460
rect 120810 143352 120816 143404
rect 120868 143392 120874 143404
rect 133138 143392 133144 143404
rect 120868 143364 133144 143392
rect 120868 143352 120874 143364
rect 133138 143352 133144 143364
rect 133196 143352 133202 143404
rect 174630 143352 174636 143404
rect 174688 143392 174694 143404
rect 179690 143392 179696 143404
rect 174688 143364 179696 143392
rect 174688 143352 174694 143364
rect 179690 143352 179696 143364
rect 179748 143352 179754 143404
rect 185670 143352 185676 143404
rect 185728 143392 185734 143404
rect 187988 143392 188016 143432
rect 193674 143420 193680 143432
rect 193732 143420 193738 143472
rect 195054 143392 195060 143404
rect 185728 143364 188016 143392
rect 188080 143364 195060 143392
rect 185728 143352 185734 143364
rect 115106 143284 115112 143336
rect 115164 143324 115170 143336
rect 123754 143324 123760 143336
rect 115164 143296 123760 143324
rect 115164 143284 115170 143296
rect 123754 143284 123760 143296
rect 123812 143284 123818 143336
rect 123846 143284 123852 143336
rect 123904 143324 123910 143336
rect 124858 143324 124864 143336
rect 123904 143296 124864 143324
rect 123904 143284 123910 143296
rect 124858 143284 124864 143296
rect 124916 143284 124922 143336
rect 131206 143284 131212 143336
rect 131264 143324 131270 143336
rect 135438 143324 135444 143336
rect 131264 143296 135444 143324
rect 131264 143284 131270 143296
rect 135438 143284 135444 143296
rect 135496 143284 135502 143336
rect 172974 143284 172980 143336
rect 173032 143324 173038 143336
rect 178402 143324 178408 143336
rect 173032 143296 178408 143324
rect 173032 143284 173038 143296
rect 178402 143284 178408 143296
rect 178460 143284 178466 143336
rect 180766 143296 182496 143324
rect 122190 143216 122196 143268
rect 122248 143256 122254 143268
rect 136634 143256 136640 143268
rect 122248 143228 136640 143256
rect 122248 143216 122254 143228
rect 136634 143216 136640 143228
rect 136692 143216 136698 143268
rect 176562 143216 176568 143268
rect 176620 143256 176626 143268
rect 180766 143256 180794 143296
rect 182468 143256 182496 143296
rect 185946 143284 185952 143336
rect 186004 143324 186010 143336
rect 188080 143324 188108 143364
rect 195054 143352 195060 143364
rect 195112 143352 195118 143404
rect 189534 143324 189540 143336
rect 186004 143296 188108 143324
rect 188264 143296 189540 143324
rect 186004 143284 186010 143296
rect 188264 143256 188292 143296
rect 189534 143284 189540 143296
rect 189592 143284 189598 143336
rect 195238 143324 195244 143336
rect 190426 143296 195244 143324
rect 176620 143228 180794 143256
rect 182100 143228 182404 143256
rect 182468 143228 188292 143256
rect 176620 143216 176626 143228
rect 114002 143148 114008 143200
rect 114060 143188 114066 143200
rect 129550 143188 129556 143200
rect 114060 143160 129556 143188
rect 114060 143148 114066 143160
rect 129550 143148 129556 143160
rect 129608 143148 129614 143200
rect 129826 143148 129832 143200
rect 129884 143188 129890 143200
rect 135898 143188 135904 143200
rect 129884 143160 135904 143188
rect 129884 143148 129890 143160
rect 135898 143148 135904 143160
rect 135956 143148 135962 143200
rect 169662 143148 169668 143200
rect 169720 143188 169726 143200
rect 179598 143188 179604 143200
rect 169720 143160 179604 143188
rect 169720 143148 169726 143160
rect 179598 143148 179604 143160
rect 179656 143148 179662 143200
rect 118326 143080 118332 143132
rect 118384 143120 118390 143132
rect 134794 143120 134800 143132
rect 118384 143092 134800 143120
rect 118384 143080 118390 143092
rect 134794 143080 134800 143092
rect 134852 143080 134858 143132
rect 177390 143080 177396 143132
rect 177448 143120 177454 143132
rect 179414 143120 179420 143132
rect 177448 143092 179420 143120
rect 177448 143080 177454 143092
rect 179414 143080 179420 143092
rect 179472 143080 179478 143132
rect 115566 143012 115572 143064
rect 115624 143052 115630 143064
rect 132586 143052 132592 143064
rect 115624 143024 132592 143052
rect 115624 143012 115630 143024
rect 132586 143012 132592 143024
rect 132644 143012 132650 143064
rect 170214 143012 170220 143064
rect 170272 143052 170278 143064
rect 182100 143052 182128 143228
rect 170272 143024 182128 143052
rect 182376 143052 182404 143228
rect 188430 143216 188436 143268
rect 188488 143256 188494 143268
rect 190426 143256 190454 143296
rect 195238 143284 195244 143296
rect 195296 143284 195302 143336
rect 188488 143228 190454 143256
rect 188488 143216 188494 143228
rect 182450 143148 182456 143200
rect 182508 143188 182514 143200
rect 196434 143188 196440 143200
rect 182508 143160 196440 143188
rect 182508 143148 182514 143160
rect 196434 143148 196440 143160
rect 196492 143148 196498 143200
rect 184474 143080 184480 143132
rect 184532 143120 184538 143132
rect 197998 143120 198004 143132
rect 184532 143092 198004 143120
rect 184532 143080 184538 143092
rect 197998 143080 198004 143092
rect 198056 143080 198062 143132
rect 191098 143052 191104 143064
rect 182376 143024 191104 143052
rect 170272 143012 170278 143024
rect 191098 143012 191104 143024
rect 191156 143012 191162 143064
rect 120902 142944 120908 142996
rect 120960 142984 120966 142996
rect 139762 142984 139768 142996
rect 120960 142956 139768 142984
rect 120960 142944 120966 142956
rect 139762 142944 139768 142956
rect 139820 142944 139826 142996
rect 168282 142944 168288 142996
rect 168340 142984 168346 142996
rect 182082 142984 182088 142996
rect 168340 142956 182088 142984
rect 168340 142944 168346 142956
rect 182082 142944 182088 142956
rect 182140 142944 182146 142996
rect 120994 142876 121000 142928
rect 121052 142916 121058 142928
rect 141510 142916 141516 142928
rect 121052 142888 141516 142916
rect 121052 142876 121058 142888
rect 141510 142876 141516 142888
rect 141568 142876 141574 142928
rect 166902 142876 166908 142928
rect 166960 142916 166966 142928
rect 191190 142916 191196 142928
rect 166960 142888 191196 142916
rect 166960 142876 166966 142888
rect 191190 142876 191196 142888
rect 191248 142876 191254 142928
rect 121086 142808 121092 142860
rect 121144 142848 121150 142860
rect 151354 142848 151360 142860
rect 121144 142820 151360 142848
rect 121144 142808 121150 142820
rect 151354 142808 151360 142820
rect 151412 142808 151418 142860
rect 158622 142808 158628 142860
rect 158680 142848 158686 142860
rect 188246 142848 188252 142860
rect 158680 142820 188252 142848
rect 158680 142808 158686 142820
rect 188246 142808 188252 142820
rect 188304 142808 188310 142860
rect 119614 142740 119620 142792
rect 119672 142780 119678 142792
rect 128446 142780 128452 142792
rect 119672 142752 128452 142780
rect 119672 142740 119678 142752
rect 128446 142740 128452 142752
rect 128504 142740 128510 142792
rect 129366 142740 129372 142792
rect 129424 142780 129430 142792
rect 131574 142780 131580 142792
rect 129424 142752 131580 142780
rect 129424 142740 129430 142752
rect 131574 142740 131580 142752
rect 131632 142740 131638 142792
rect 183094 142740 183100 142792
rect 183152 142780 183158 142792
rect 190914 142780 190920 142792
rect 183152 142752 190920 142780
rect 183152 142740 183158 142752
rect 190914 142740 190920 142752
rect 190972 142740 190978 142792
rect 123754 142672 123760 142724
rect 123812 142712 123818 142724
rect 129090 142712 129096 142724
rect 123812 142684 129096 142712
rect 123812 142672 123818 142684
rect 129090 142672 129096 142684
rect 129148 142672 129154 142724
rect 131206 142672 131212 142724
rect 131264 142712 131270 142724
rect 131390 142712 131396 142724
rect 131264 142684 131396 142712
rect 131264 142672 131270 142684
rect 131390 142672 131396 142684
rect 131448 142672 131454 142724
rect 177942 142672 177948 142724
rect 178000 142712 178006 142724
rect 178218 142712 178224 142724
rect 178000 142684 178224 142712
rect 178000 142672 178006 142684
rect 178218 142672 178224 142684
rect 178276 142672 178282 142724
rect 182082 142672 182088 142724
rect 182140 142712 182146 142724
rect 189442 142712 189448 142724
rect 182140 142684 189448 142712
rect 182140 142672 182146 142684
rect 189442 142672 189448 142684
rect 189500 142672 189506 142724
rect 183738 142604 183744 142656
rect 183796 142644 183802 142656
rect 188430 142644 188436 142656
rect 183796 142616 188436 142644
rect 183796 142604 183802 142616
rect 188430 142604 188436 142616
rect 188488 142604 188494 142656
rect 129918 142264 129924 142316
rect 129976 142304 129982 142316
rect 134242 142304 134248 142316
rect 129976 142276 134248 142304
rect 129976 142264 129982 142276
rect 134242 142264 134248 142276
rect 134300 142264 134306 142316
rect 129734 142196 129740 142248
rect 129792 142236 129798 142248
rect 133874 142236 133880 142248
rect 129792 142208 133880 142236
rect 129792 142196 129798 142208
rect 133874 142196 133880 142208
rect 133932 142196 133938 142248
rect 155678 142196 155684 142248
rect 155736 142236 155742 142248
rect 157334 142236 157340 142248
rect 155736 142208 157340 142236
rect 155736 142196 155742 142208
rect 157334 142196 157340 142208
rect 157392 142196 157398 142248
rect 159174 142196 159180 142248
rect 159232 142236 159238 142248
rect 161474 142236 161480 142248
rect 159232 142208 161480 142236
rect 159232 142196 159238 142208
rect 161474 142196 161480 142208
rect 161532 142196 161538 142248
rect 3418 142128 3424 142180
rect 3476 142168 3482 142180
rect 183738 142168 183744 142180
rect 3476 142140 183744 142168
rect 3476 142128 3482 142140
rect 183738 142128 183744 142140
rect 183796 142128 183802 142180
rect 185946 142128 185952 142180
rect 186004 142168 186010 142180
rect 187878 142168 187884 142180
rect 186004 142140 187884 142168
rect 186004 142128 186010 142140
rect 187878 142128 187884 142140
rect 187936 142128 187942 142180
rect 161474 142060 161480 142112
rect 161532 142100 161538 142112
rect 192294 142100 192300 142112
rect 161532 142072 192300 142100
rect 161532 142060 161538 142072
rect 192294 142060 192300 142072
rect 192352 142060 192358 142112
rect 118418 141992 118424 142044
rect 118476 142032 118482 142044
rect 126882 142032 126888 142044
rect 118476 142004 126888 142032
rect 118476 141992 118482 142004
rect 126882 141992 126888 142004
rect 126940 141992 126946 142044
rect 115474 141924 115480 141976
rect 115532 141964 115538 141976
rect 127342 141964 127348 141976
rect 115532 141936 127348 141964
rect 115532 141924 115538 141936
rect 127342 141924 127348 141936
rect 127400 141924 127406 141976
rect 180334 141924 180340 141976
rect 180392 141964 180398 141976
rect 187234 141964 187240 141976
rect 180392 141936 187240 141964
rect 180392 141924 180398 141936
rect 187234 141924 187240 141936
rect 187292 141924 187298 141976
rect 115290 141856 115296 141908
rect 115348 141896 115354 141908
rect 130378 141896 130384 141908
rect 115348 141868 130384 141896
rect 115348 141856 115354 141868
rect 130378 141856 130384 141868
rect 130436 141856 130442 141908
rect 182082 141856 182088 141908
rect 182140 141896 182146 141908
rect 192110 141896 192116 141908
rect 182140 141868 192116 141896
rect 182140 141856 182146 141868
rect 192110 141856 192116 141868
rect 192168 141856 192174 141908
rect 116578 141788 116584 141840
rect 116636 141828 116642 141840
rect 131758 141828 131764 141840
rect 116636 141800 131764 141828
rect 116636 141788 116642 141800
rect 131758 141788 131764 141800
rect 131816 141788 131822 141840
rect 183186 141788 183192 141840
rect 183244 141828 183250 141840
rect 196434 141828 196440 141840
rect 183244 141800 196440 141828
rect 183244 141788 183250 141800
rect 196434 141788 196440 141800
rect 196492 141788 196498 141840
rect 113634 141720 113640 141772
rect 113692 141760 113698 141772
rect 132862 141760 132868 141772
rect 113692 141732 132868 141760
rect 113692 141720 113698 141732
rect 132862 141720 132868 141732
rect 132920 141720 132926 141772
rect 175182 141720 175188 141772
rect 175240 141760 175246 141772
rect 187326 141760 187332 141772
rect 175240 141732 187332 141760
rect 175240 141720 175246 141732
rect 187326 141720 187332 141732
rect 187384 141720 187390 141772
rect 118142 141652 118148 141704
rect 118200 141692 118206 141704
rect 140314 141692 140320 141704
rect 118200 141664 140320 141692
rect 118200 141652 118206 141664
rect 140314 141652 140320 141664
rect 140372 141652 140378 141704
rect 173526 141652 173532 141704
rect 173584 141692 173590 141704
rect 190822 141692 190828 141704
rect 173584 141664 190828 141692
rect 173584 141652 173590 141664
rect 190822 141652 190828 141664
rect 190880 141652 190886 141704
rect 114186 141584 114192 141636
rect 114244 141624 114250 141636
rect 137002 141624 137008 141636
rect 114244 141596 137008 141624
rect 114244 141584 114250 141596
rect 137002 141584 137008 141596
rect 137060 141584 137066 141636
rect 171870 141584 171876 141636
rect 171928 141624 171934 141636
rect 189350 141624 189356 141636
rect 171928 141596 189356 141624
rect 171928 141584 171934 141596
rect 189350 141584 189356 141596
rect 189408 141584 189414 141636
rect 119982 141516 119988 141568
rect 120040 141556 120046 141568
rect 151906 141556 151912 141568
rect 120040 141528 151912 141556
rect 120040 141516 120046 141528
rect 151906 141516 151912 141528
rect 151964 141516 151970 141568
rect 167454 141516 167460 141568
rect 167512 141556 167518 141568
rect 192202 141556 192208 141568
rect 167512 141528 192208 141556
rect 167512 141516 167518 141528
rect 192202 141516 192208 141528
rect 192260 141516 192266 141568
rect 119522 141448 119528 141500
rect 119580 141488 119586 141500
rect 142246 141488 142252 141500
rect 119580 141460 142252 141488
rect 119580 141448 119586 141460
rect 142246 141448 142252 141460
rect 142304 141448 142310 141500
rect 164326 141448 164332 141500
rect 164384 141488 164390 141500
rect 189534 141488 189540 141500
rect 164384 141460 189540 141488
rect 164384 141448 164390 141460
rect 189534 141448 189540 141460
rect 189592 141448 189598 141500
rect 119430 141380 119436 141432
rect 119488 141420 119494 141432
rect 153562 141420 153568 141432
rect 119488 141392 153568 141420
rect 119488 141380 119494 141392
rect 153562 141380 153568 141392
rect 153620 141380 153626 141432
rect 162854 141380 162860 141432
rect 162912 141420 162918 141432
rect 197998 141420 198004 141432
rect 162912 141392 198004 141420
rect 162912 141380 162918 141392
rect 197998 141380 198004 141392
rect 198056 141380 198062 141432
rect 120994 141312 121000 141364
rect 121052 141352 121058 141364
rect 126514 141352 126520 141364
rect 121052 141324 126520 141352
rect 121052 141312 121058 141324
rect 126514 141312 126520 141324
rect 126572 141312 126578 141364
rect 118234 141244 118240 141296
rect 118292 141284 118298 141296
rect 125410 141284 125416 141296
rect 118292 141256 125416 141284
rect 118292 141244 118298 141256
rect 125410 141244 125416 141256
rect 125468 141244 125474 141296
rect 129550 141040 129556 141092
rect 129608 141080 129614 141092
rect 187970 141080 187976 141092
rect 129608 141052 187976 141080
rect 129608 141040 129614 141052
rect 187970 141040 187976 141052
rect 188028 141040 188034 141092
rect 117774 140972 117780 141024
rect 117832 141012 117838 141024
rect 182082 141012 182088 141024
rect 117832 140984 182088 141012
rect 117832 140972 117838 140984
rect 182082 140972 182088 140984
rect 182140 140972 182146 141024
rect 8938 140904 8944 140956
rect 8996 140944 9002 140956
rect 182818 140944 182824 140956
rect 8996 140916 182824 140944
rect 8996 140904 9002 140916
rect 182818 140904 182824 140916
rect 182876 140904 182882 140956
rect 184566 140904 184572 140956
rect 184624 140944 184630 140956
rect 188430 140944 188436 140956
rect 184624 140916 188436 140944
rect 184624 140904 184630 140916
rect 188430 140904 188436 140916
rect 188488 140904 188494 140956
rect 126882 140836 126888 140888
rect 126940 140876 126946 140888
rect 464338 140876 464344 140888
rect 126940 140848 464344 140876
rect 126940 140836 126946 140848
rect 464338 140836 464344 140848
rect 464396 140836 464402 140888
rect 124582 140768 124588 140820
rect 124640 140808 124646 140820
rect 124950 140808 124956 140820
rect 124640 140780 124956 140808
rect 124640 140768 124646 140780
rect 124950 140768 124956 140780
rect 125008 140808 125014 140820
rect 485038 140808 485044 140820
rect 125008 140780 485044 140808
rect 125008 140768 125014 140780
rect 485038 140768 485044 140780
rect 485096 140768 485102 140820
rect 125962 140700 125968 140752
rect 126020 140740 126026 140752
rect 126606 140740 126612 140752
rect 126020 140712 126612 140740
rect 126020 140700 126026 140712
rect 126606 140700 126612 140712
rect 126664 140700 126670 140752
rect 126974 140700 126980 140752
rect 127032 140740 127038 140752
rect 127710 140740 127716 140752
rect 127032 140712 127716 140740
rect 127032 140700 127038 140712
rect 127710 140700 127716 140712
rect 127768 140700 127774 140752
rect 131298 140700 131304 140752
rect 131356 140740 131362 140752
rect 132310 140740 132316 140752
rect 131356 140712 132316 140740
rect 131356 140700 131362 140712
rect 132310 140700 132316 140712
rect 132368 140700 132374 140752
rect 178034 140700 178040 140752
rect 178092 140740 178098 140752
rect 178954 140740 178960 140752
rect 178092 140712 178960 140740
rect 178092 140700 178098 140712
rect 178954 140700 178960 140712
rect 179012 140700 179018 140752
rect 184750 140700 184756 140752
rect 184808 140740 184814 140752
rect 192018 140740 192024 140752
rect 184808 140712 192024 140740
rect 184808 140700 184814 140712
rect 192018 140700 192024 140712
rect 192076 140700 192082 140752
rect 120626 140632 120632 140684
rect 120684 140672 120690 140684
rect 126330 140672 126336 140684
rect 120684 140644 126336 140672
rect 120684 140632 120690 140644
rect 126330 140632 126336 140644
rect 126388 140632 126394 140684
rect 172514 140632 172520 140684
rect 172572 140672 172578 140684
rect 180150 140672 180156 140684
rect 172572 140644 180156 140672
rect 172572 140632 172578 140644
rect 180150 140632 180156 140644
rect 180208 140632 180214 140684
rect 118142 140564 118148 140616
rect 118200 140604 118206 140616
rect 126238 140604 126244 140616
rect 118200 140576 126244 140604
rect 118200 140564 118206 140576
rect 126238 140564 126244 140576
rect 126296 140564 126302 140616
rect 171686 140564 171692 140616
rect 171744 140604 171750 140616
rect 179046 140604 179052 140616
rect 171744 140576 179052 140604
rect 171744 140564 171750 140576
rect 179046 140564 179052 140576
rect 179104 140564 179110 140616
rect 180242 140564 180248 140616
rect 180300 140604 180306 140616
rect 188246 140604 188252 140616
rect 180300 140576 188252 140604
rect 180300 140564 180306 140576
rect 188246 140564 188252 140576
rect 188304 140564 188310 140616
rect 117866 140496 117872 140548
rect 117924 140536 117930 140548
rect 126422 140536 126428 140548
rect 117924 140508 126428 140536
rect 117924 140496 117930 140508
rect 126422 140496 126428 140508
rect 126480 140496 126486 140548
rect 184106 140496 184112 140548
rect 184164 140536 184170 140548
rect 188614 140536 188620 140548
rect 184164 140508 188620 140536
rect 184164 140496 184170 140508
rect 188614 140496 188620 140508
rect 188672 140496 188678 140548
rect 120718 140428 120724 140480
rect 120776 140468 120782 140480
rect 147030 140468 147036 140480
rect 120776 140440 147036 140468
rect 120776 140428 120782 140440
rect 147030 140428 147036 140440
rect 147088 140428 147094 140480
rect 182910 140428 182916 140480
rect 182968 140468 182974 140480
rect 190822 140468 190828 140480
rect 182968 140440 190828 140468
rect 182968 140428 182974 140440
rect 190822 140428 190828 140440
rect 190880 140428 190886 140480
rect 119246 140360 119252 140412
rect 119304 140400 119310 140412
rect 146938 140400 146944 140412
rect 119304 140372 146944 140400
rect 119304 140360 119310 140372
rect 146938 140360 146944 140372
rect 146996 140360 147002 140412
rect 185762 140360 185768 140412
rect 185820 140400 185826 140412
rect 193858 140400 193864 140412
rect 185820 140372 193864 140400
rect 185820 140360 185826 140372
rect 193858 140360 193864 140372
rect 193916 140360 193922 140412
rect 120534 140292 120540 140344
rect 120592 140332 120598 140344
rect 148226 140332 148232 140344
rect 120592 140304 148232 140332
rect 120592 140292 120598 140304
rect 148226 140292 148232 140304
rect 148284 140292 148290 140344
rect 181438 140292 181444 140344
rect 181496 140332 181502 140344
rect 189902 140332 189908 140344
rect 181496 140304 189908 140332
rect 181496 140292 181502 140304
rect 189902 140292 189908 140304
rect 189960 140292 189966 140344
rect 117958 140224 117964 140276
rect 118016 140264 118022 140276
rect 145558 140264 145564 140276
rect 118016 140236 145564 140264
rect 118016 140224 118022 140236
rect 145558 140224 145564 140236
rect 145616 140224 145622 140276
rect 180058 140224 180064 140276
rect 180116 140264 180122 140276
rect 189350 140264 189356 140276
rect 180116 140236 189356 140264
rect 180116 140224 180122 140236
rect 189350 140224 189356 140236
rect 189408 140224 189414 140276
rect 118050 140156 118056 140208
rect 118108 140196 118114 140208
rect 147950 140196 147956 140208
rect 118108 140168 147956 140196
rect 118108 140156 118114 140168
rect 147950 140156 147956 140168
rect 148008 140156 148014 140208
rect 184290 140156 184296 140208
rect 184348 140196 184354 140208
rect 189810 140196 189816 140208
rect 184348 140168 189816 140196
rect 184348 140156 184354 140168
rect 189810 140156 189816 140168
rect 189868 140156 189874 140208
rect 121914 140088 121920 140140
rect 121972 140128 121978 140140
rect 152458 140128 152464 140140
rect 121972 140100 152464 140128
rect 121972 140088 121978 140100
rect 152458 140088 152464 140100
rect 152516 140088 152522 140140
rect 169846 140088 169852 140140
rect 169904 140128 169910 140140
rect 169904 140100 184060 140128
rect 169904 140088 169910 140100
rect 119338 140020 119344 140072
rect 119396 140060 119402 140072
rect 129274 140060 129280 140072
rect 119396 140032 129280 140060
rect 119396 140020 119402 140032
rect 129274 140020 129280 140032
rect 129332 140020 129338 140072
rect 129734 140020 129740 140072
rect 129792 140060 129798 140072
rect 184032 140060 184060 140100
rect 184658 140088 184664 140140
rect 184716 140128 184722 140140
rect 187234 140128 187240 140140
rect 184716 140100 187240 140128
rect 184716 140088 184722 140100
rect 187234 140088 187240 140100
rect 187292 140088 187298 140140
rect 187326 140060 187332 140072
rect 129792 140032 180794 140060
rect 184032 140032 187332 140060
rect 129792 140020 129798 140032
rect 130010 139952 130016 140004
rect 130068 139992 130074 140004
rect 130470 139992 130476 140004
rect 130068 139964 130476 139992
rect 130068 139952 130074 139964
rect 130470 139952 130476 139964
rect 130528 139952 130534 140004
rect 180766 139992 180794 140032
rect 187326 140020 187332 140032
rect 187384 140020 187390 140072
rect 188062 139992 188068 140004
rect 180766 139964 188068 139992
rect 188062 139952 188068 139964
rect 188120 139952 188126 140004
rect 194042 139992 194048 140004
rect 188172 139964 194048 139992
rect 184382 139884 184388 139936
rect 184440 139924 184446 139936
rect 188172 139924 188200 139964
rect 194042 139952 194048 139964
rect 194100 139952 194106 140004
rect 184440 139896 188200 139924
rect 184440 139884 184446 139896
rect 188614 139884 188620 139936
rect 188672 139924 188678 139936
rect 192294 139924 192300 139936
rect 188672 139896 192300 139924
rect 188672 139884 188678 139896
rect 192294 139884 192300 139896
rect 192352 139884 192358 139936
rect 171134 139816 171140 139868
rect 171192 139856 171198 139868
rect 196250 139856 196256 139868
rect 171192 139828 185624 139856
rect 171192 139816 171198 139828
rect 128814 139748 128820 139800
rect 128872 139788 128878 139800
rect 183462 139788 183468 139800
rect 128872 139760 183468 139788
rect 128872 139748 128878 139760
rect 183462 139748 183468 139760
rect 183520 139748 183526 139800
rect 125870 139680 125876 139732
rect 125928 139720 125934 139732
rect 184658 139720 184664 139732
rect 125928 139692 184664 139720
rect 125928 139680 125934 139692
rect 184658 139680 184664 139692
rect 184716 139680 184722 139732
rect 185596 139720 185624 139828
rect 190426 139828 196256 139856
rect 190426 139720 190454 139828
rect 196250 139816 196256 139828
rect 196308 139816 196314 139868
rect 185596 139692 190454 139720
rect 118694 139612 118700 139664
rect 118752 139652 118758 139664
rect 180058 139652 180064 139664
rect 118752 139624 180064 139652
rect 118752 139612 118758 139624
rect 180058 139612 180064 139624
rect 180116 139612 180122 139664
rect 122834 139544 122840 139596
rect 122892 139584 122898 139596
rect 123846 139584 123852 139596
rect 122892 139556 123852 139584
rect 122892 139544 122898 139556
rect 123846 139544 123852 139556
rect 123904 139584 123910 139596
rect 184566 139584 184572 139596
rect 123904 139556 184572 139584
rect 123904 139544 123910 139556
rect 184566 139544 184572 139556
rect 184624 139544 184630 139596
rect 31018 139476 31024 139528
rect 31076 139516 31082 139528
rect 181162 139516 181168 139528
rect 31076 139488 181168 139516
rect 31076 139476 31082 139488
rect 181162 139476 181168 139488
rect 181220 139476 181226 139528
rect 185578 139476 185584 139528
rect 185636 139516 185642 139528
rect 187418 139516 187424 139528
rect 185636 139488 187424 139516
rect 185636 139476 185642 139488
rect 187418 139476 187424 139488
rect 187476 139476 187482 139528
rect 13078 139408 13084 139460
rect 13136 139448 13142 139460
rect 185026 139448 185032 139460
rect 13136 139420 185032 139448
rect 13136 139408 13142 139420
rect 185026 139408 185032 139420
rect 185084 139408 185090 139460
rect 186130 139408 186136 139460
rect 186188 139448 186194 139460
rect 187142 139448 187148 139460
rect 186188 139420 187148 139448
rect 186188 139408 186194 139420
rect 187142 139408 187148 139420
rect 187200 139408 187206 139460
rect 188246 139448 188252 139460
rect 187896 139420 188252 139448
rect 186038 139340 186044 139392
rect 186096 139380 186102 139392
rect 186866 139380 186872 139392
rect 186096 139352 186872 139380
rect 186096 139340 186102 139352
rect 186866 139340 186872 139352
rect 186924 139340 186930 139392
rect 187896 139312 187924 139420
rect 188246 139408 188252 139420
rect 188304 139408 188310 139460
rect 187970 139340 187976 139392
rect 188028 139380 188034 139392
rect 580166 139380 580172 139392
rect 188028 139352 580172 139380
rect 188028 139340 188034 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 187896 139284 188016 139312
rect 187988 139256 188016 139284
rect 187970 139204 187976 139256
rect 188028 139204 188034 139256
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 118694 137952 118700 137964
rect 3568 137924 118700 137952
rect 3568 137912 3574 137924
rect 118694 137912 118700 137924
rect 118752 137912 118758 137964
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 31018 111772 31024 111784
rect 3200 111744 31024 111772
rect 3200 111732 3206 111744
rect 31018 111732 31024 111744
rect 31076 111732 31082 111784
rect 464338 86912 464344 86964
rect 464396 86952 464402 86964
rect 580166 86952 580172 86964
rect 464396 86924 580172 86952
rect 464396 86912 464402 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 117774 85524 117780 85536
rect 3568 85496 117780 85524
rect 3568 85484 3574 85496
rect 117774 85484 117780 85496
rect 117832 85484 117838 85536
rect 150682 81212 177988 81240
rect 123018 81064 123024 81116
rect 123076 81104 123082 81116
rect 123076 81076 132494 81104
rect 123076 81064 123082 81076
rect 132466 81036 132494 81076
rect 122806 81008 124720 81036
rect 132466 81008 140774 81036
rect 119062 80928 119068 80980
rect 119120 80968 119126 80980
rect 122806 80968 122834 81008
rect 119120 80940 122834 80968
rect 119120 80928 119126 80940
rect 122282 80860 122288 80912
rect 122340 80900 122346 80912
rect 123018 80900 123024 80912
rect 122340 80872 123024 80900
rect 122340 80860 122346 80872
rect 123018 80860 123024 80872
rect 123076 80860 123082 80912
rect 124692 80900 124720 81008
rect 133846 80940 138704 80968
rect 133846 80900 133874 80940
rect 124692 80872 133874 80900
rect 108206 80792 108212 80844
rect 108264 80832 108270 80844
rect 108264 80804 132172 80832
rect 108264 80792 108270 80804
rect 85574 80724 85580 80776
rect 85632 80764 85638 80776
rect 105630 80764 105636 80776
rect 85632 80736 105636 80764
rect 85632 80724 85638 80736
rect 105630 80724 105636 80736
rect 105688 80764 105694 80776
rect 105688 80736 125594 80764
rect 105688 80724 105694 80736
rect 71774 80656 71780 80708
rect 71832 80696 71838 80708
rect 108206 80696 108212 80708
rect 71832 80668 108212 80696
rect 71832 80656 71838 80668
rect 108206 80656 108212 80668
rect 108264 80656 108270 80708
rect 119982 80656 119988 80708
rect 120040 80696 120046 80708
rect 125566 80696 125594 80736
rect 132144 80708 132172 80804
rect 131942 80696 131948 80708
rect 120040 80668 122834 80696
rect 125566 80668 131948 80696
rect 120040 80656 120046 80668
rect 104250 80424 104256 80436
rect 104176 80396 104256 80424
rect 104176 80232 104204 80396
rect 104250 80384 104256 80396
rect 104308 80384 104314 80436
rect 122806 80424 122834 80668
rect 131942 80656 131948 80668
rect 132000 80656 132006 80708
rect 132126 80656 132132 80708
rect 132184 80656 132190 80708
rect 138676 80696 138704 80940
rect 140746 80764 140774 81008
rect 140746 80736 146754 80764
rect 138676 80668 144822 80696
rect 132218 80588 132224 80640
rect 132276 80628 132282 80640
rect 132276 80600 142154 80628
rect 132276 80588 132282 80600
rect 142126 80492 142154 80600
rect 142126 80464 144500 80492
rect 132218 80424 132224 80436
rect 122806 80396 132224 80424
rect 132218 80384 132224 80396
rect 132276 80384 132282 80436
rect 131850 80316 131856 80368
rect 131908 80356 131914 80368
rect 131908 80328 142154 80356
rect 131908 80316 131914 80328
rect 122806 80260 125594 80288
rect 104158 80180 104164 80232
rect 104216 80180 104222 80232
rect 110966 80044 110972 80096
rect 111024 80084 111030 80096
rect 122806 80084 122834 80260
rect 125566 80152 125594 80260
rect 131022 80248 131028 80300
rect 131080 80288 131086 80300
rect 131080 80260 141970 80288
rect 131080 80248 131086 80260
rect 127526 80180 127532 80232
rect 127584 80220 127590 80232
rect 127584 80192 141878 80220
rect 127584 80180 127590 80192
rect 125566 80124 140866 80152
rect 111024 80056 122834 80084
rect 111024 80044 111030 80056
rect 131942 80044 131948 80096
rect 132000 80084 132006 80096
rect 132000 80056 139118 80084
rect 132000 80044 132006 80056
rect 132742 79988 133230 80016
rect 132742 79960 132770 79988
rect 132724 79908 132730 79960
rect 132782 79908 132788 79960
rect 133092 79908 133098 79960
rect 133150 79908 133156 79960
rect 126974 79840 126980 79892
rect 127032 79880 127038 79892
rect 132908 79880 132914 79892
rect 127032 79852 132914 79880
rect 127032 79840 127038 79852
rect 132908 79840 132914 79852
rect 132966 79840 132972 79892
rect 119246 79636 119252 79688
rect 119304 79676 119310 79688
rect 132402 79676 132408 79688
rect 119304 79648 132408 79676
rect 119304 79636 119310 79648
rect 132402 79636 132408 79648
rect 132460 79636 132466 79688
rect 133110 79620 133138 79908
rect 106826 79568 106832 79620
rect 106884 79608 106890 79620
rect 106884 79580 127664 79608
rect 106884 79568 106890 79580
rect 113818 79500 113824 79552
rect 113876 79540 113882 79552
rect 125686 79540 125692 79552
rect 113876 79512 125692 79540
rect 113876 79500 113882 79512
rect 125686 79500 125692 79512
rect 125744 79540 125750 79552
rect 127434 79540 127440 79552
rect 125744 79512 127440 79540
rect 125744 79500 125750 79512
rect 127434 79500 127440 79512
rect 127492 79500 127498 79552
rect 111058 79432 111064 79484
rect 111116 79472 111122 79484
rect 125594 79472 125600 79484
rect 111116 79444 125600 79472
rect 111116 79432 111122 79444
rect 125594 79432 125600 79444
rect 125652 79472 125658 79484
rect 127526 79472 127532 79484
rect 125652 79444 127532 79472
rect 125652 79432 125658 79444
rect 127526 79432 127532 79444
rect 127584 79432 127590 79484
rect 127636 79472 127664 79580
rect 133046 79568 133052 79620
rect 133104 79580 133138 79620
rect 133202 79608 133230 79988
rect 133754 79988 134886 80016
rect 133368 79908 133374 79960
rect 133426 79908 133432 79960
rect 133644 79908 133650 79960
rect 133702 79908 133708 79960
rect 133386 79756 133414 79908
rect 133460 79840 133466 79892
rect 133518 79880 133524 79892
rect 133518 79840 133552 79880
rect 133386 79716 133420 79756
rect 133414 79704 133420 79716
rect 133472 79704 133478 79756
rect 133322 79608 133328 79620
rect 133202 79580 133328 79608
rect 133104 79568 133110 79580
rect 133322 79568 133328 79580
rect 133380 79568 133386 79620
rect 132862 79500 132868 79552
rect 132920 79540 132926 79552
rect 133524 79540 133552 79840
rect 133662 79688 133690 79908
rect 133754 79812 133782 79988
rect 134858 79960 134886 79988
rect 139090 79960 139118 80056
rect 140838 79960 140866 80124
rect 141850 79960 141878 80192
rect 133828 79908 133834 79960
rect 133886 79908 133892 79960
rect 134012 79948 134018 79960
rect 133984 79908 134018 79948
rect 134070 79908 134076 79960
rect 134104 79908 134110 79960
rect 134162 79908 134168 79960
rect 134656 79908 134662 79960
rect 134714 79908 134720 79960
rect 134840 79908 134846 79960
rect 134898 79908 134904 79960
rect 135300 79948 135306 79960
rect 135226 79920 135306 79948
rect 133846 79880 133874 79908
rect 133846 79852 133920 79880
rect 133892 79824 133920 79852
rect 133984 79824 134012 79908
rect 133754 79784 133828 79812
rect 133662 79648 133696 79688
rect 133690 79636 133696 79648
rect 133748 79636 133754 79688
rect 133598 79568 133604 79620
rect 133656 79608 133662 79620
rect 133800 79608 133828 79784
rect 133874 79772 133880 79824
rect 133932 79772 133938 79824
rect 133966 79772 133972 79824
rect 134024 79772 134030 79824
rect 134122 79756 134150 79908
rect 134472 79840 134478 79892
rect 134530 79840 134536 79892
rect 134196 79772 134202 79824
rect 134254 79772 134260 79824
rect 134058 79704 134064 79756
rect 134116 79716 134150 79756
rect 134116 79704 134122 79716
rect 134214 79620 134242 79772
rect 133656 79580 133828 79608
rect 133656 79568 133662 79580
rect 134150 79568 134156 79620
rect 134208 79580 134242 79620
rect 134208 79568 134214 79580
rect 134334 79568 134340 79620
rect 134392 79568 134398 79620
rect 134490 79608 134518 79840
rect 134674 79824 134702 79908
rect 134932 79880 134938 79892
rect 134904 79840 134938 79880
rect 134990 79840 134996 79892
rect 134656 79772 134662 79824
rect 134714 79772 134720 79824
rect 134748 79704 134754 79756
rect 134806 79704 134812 79756
rect 134444 79580 134518 79608
rect 132920 79512 133552 79540
rect 132920 79500 132926 79512
rect 134352 79484 134380 79568
rect 127636 79444 133046 79472
rect 111242 79364 111248 79416
rect 111300 79404 111306 79416
rect 128354 79404 128360 79416
rect 111300 79376 128360 79404
rect 111300 79364 111306 79376
rect 128354 79364 128360 79376
rect 128412 79404 128418 79416
rect 131022 79404 131028 79416
rect 128412 79376 131028 79404
rect 128412 79364 128418 79376
rect 131022 79364 131028 79376
rect 131080 79364 131086 79416
rect 132678 79404 132684 79416
rect 131132 79376 132684 79404
rect 100110 79296 100116 79348
rect 100168 79336 100174 79348
rect 100294 79336 100300 79348
rect 100168 79308 100300 79336
rect 100168 79296 100174 79308
rect 100294 79296 100300 79308
rect 100352 79296 100358 79348
rect 112438 79296 112444 79348
rect 112496 79336 112502 79348
rect 130378 79336 130384 79348
rect 112496 79308 130384 79336
rect 112496 79296 112502 79308
rect 130378 79296 130384 79308
rect 130436 79336 130442 79348
rect 131132 79336 131160 79376
rect 132678 79364 132684 79376
rect 132736 79364 132742 79416
rect 133018 79404 133046 79444
rect 134334 79432 134340 79484
rect 134392 79432 134398 79484
rect 134444 79472 134472 79580
rect 134610 79500 134616 79552
rect 134668 79540 134674 79552
rect 134766 79540 134794 79704
rect 134904 79688 134932 79840
rect 134886 79636 134892 79688
rect 134944 79636 134950 79688
rect 135226 79676 135254 79920
rect 135300 79908 135306 79920
rect 135358 79908 135364 79960
rect 136220 79908 136226 79960
rect 136278 79908 136284 79960
rect 136312 79908 136318 79960
rect 136370 79908 136376 79960
rect 136588 79908 136594 79960
rect 136646 79908 136652 79960
rect 136956 79908 136962 79960
rect 137014 79908 137020 79960
rect 137048 79908 137054 79960
rect 137106 79908 137112 79960
rect 137232 79908 137238 79960
rect 137290 79908 137296 79960
rect 137508 79908 137514 79960
rect 137566 79908 137572 79960
rect 138244 79908 138250 79960
rect 138302 79908 138308 79960
rect 138888 79908 138894 79960
rect 138946 79908 138952 79960
rect 139072 79908 139078 79960
rect 139130 79908 139136 79960
rect 139440 79908 139446 79960
rect 139498 79908 139504 79960
rect 139624 79908 139630 79960
rect 139682 79908 139688 79960
rect 139716 79908 139722 79960
rect 139774 79908 139780 79960
rect 140636 79948 140642 79960
rect 140608 79908 140642 79948
rect 140694 79908 140700 79960
rect 140820 79908 140826 79960
rect 140878 79908 140884 79960
rect 141004 79908 141010 79960
rect 141062 79908 141068 79960
rect 141188 79948 141194 79960
rect 141160 79908 141194 79948
rect 141246 79908 141252 79960
rect 141556 79908 141562 79960
rect 141614 79948 141620 79960
rect 141614 79920 141786 79948
rect 141614 79908 141620 79920
rect 135760 79880 135766 79892
rect 135180 79648 135254 79676
rect 135318 79852 135766 79880
rect 134668 79512 134794 79540
rect 134668 79500 134674 79512
rect 135070 79472 135076 79484
rect 134444 79444 135076 79472
rect 135070 79432 135076 79444
rect 135128 79432 135134 79484
rect 135180 79472 135208 79648
rect 135318 79620 135346 79852
rect 135760 79840 135766 79852
rect 135818 79840 135824 79892
rect 135944 79840 135950 79892
rect 136002 79840 136008 79892
rect 136036 79840 136042 79892
rect 136094 79840 136100 79892
rect 135576 79772 135582 79824
rect 135634 79772 135640 79824
rect 135962 79812 135990 79840
rect 135824 79784 135990 79812
rect 135254 79568 135260 79620
rect 135312 79580 135346 79620
rect 135594 79620 135622 79772
rect 135594 79580 135628 79620
rect 135312 79568 135318 79580
rect 135622 79568 135628 79580
rect 135680 79568 135686 79620
rect 135824 79540 135852 79784
rect 136054 79744 136082 79840
rect 135916 79716 136082 79744
rect 135916 79608 135944 79716
rect 135990 79636 135996 79688
rect 136048 79676 136054 79688
rect 136238 79676 136266 79908
rect 136048 79648 136266 79676
rect 136048 79636 136054 79648
rect 136330 79620 136358 79908
rect 136404 79772 136410 79824
rect 136462 79772 136468 79824
rect 136422 79688 136450 79772
rect 136422 79648 136456 79688
rect 136450 79636 136456 79648
rect 136508 79636 136514 79688
rect 136606 79620 136634 79908
rect 136974 79812 137002 79908
rect 136928 79784 137002 79812
rect 136818 79704 136824 79756
rect 136876 79704 136882 79756
rect 136174 79608 136180 79620
rect 135916 79580 136180 79608
rect 136174 79568 136180 79580
rect 136232 79568 136238 79620
rect 136330 79580 136364 79620
rect 136358 79568 136364 79580
rect 136416 79568 136422 79620
rect 136542 79568 136548 79620
rect 136600 79580 136634 79620
rect 136600 79568 136606 79580
rect 135732 79512 135852 79540
rect 135732 79484 135760 79512
rect 136082 79500 136088 79552
rect 136140 79540 136146 79552
rect 136836 79540 136864 79704
rect 136928 79688 136956 79784
rect 137066 79744 137094 79908
rect 137020 79716 137094 79744
rect 136910 79636 136916 79688
rect 136968 79636 136974 79688
rect 137020 79620 137048 79716
rect 137094 79636 137100 79688
rect 137152 79676 137158 79688
rect 137250 79676 137278 79908
rect 137416 79880 137422 79892
rect 137152 79648 137278 79676
rect 137342 79852 137422 79880
rect 137152 79636 137158 79648
rect 137342 79620 137370 79852
rect 137416 79840 137422 79852
rect 137474 79840 137480 79892
rect 137526 79756 137554 79908
rect 137784 79840 137790 79892
rect 137842 79840 137848 79892
rect 137462 79704 137468 79756
rect 137520 79716 137554 79756
rect 137520 79704 137526 79716
rect 137802 79688 137830 79840
rect 137802 79648 137836 79688
rect 137830 79636 137836 79648
rect 137888 79636 137894 79688
rect 138106 79636 138112 79688
rect 138164 79676 138170 79688
rect 138262 79676 138290 79908
rect 138906 79744 138934 79908
rect 138980 79840 138986 79892
rect 139038 79840 139044 79892
rect 139458 79880 139486 79908
rect 139320 79852 139486 79880
rect 138400 79716 138934 79744
rect 138400 79688 138428 79716
rect 138164 79648 138290 79676
rect 138164 79636 138170 79648
rect 138382 79636 138388 79688
rect 138440 79636 138446 79688
rect 138474 79636 138480 79688
rect 138532 79676 138538 79688
rect 138998 79676 139026 79840
rect 138532 79648 139026 79676
rect 138532 79636 138538 79648
rect 137002 79568 137008 79620
rect 137060 79568 137066 79620
rect 137278 79568 137284 79620
rect 137336 79580 137370 79620
rect 137336 79568 137342 79580
rect 136140 79512 136864 79540
rect 139320 79540 139348 79852
rect 139642 79812 139670 79908
rect 139412 79784 139670 79812
rect 139412 79608 139440 79784
rect 139734 79744 139762 79908
rect 139808 79840 139814 79892
rect 139866 79880 139872 79892
rect 139866 79852 140084 79880
rect 139866 79840 139872 79852
rect 139504 79716 139762 79744
rect 139504 79688 139532 79716
rect 139486 79636 139492 79688
rect 139544 79636 139550 79688
rect 139578 79608 139584 79620
rect 139412 79580 139584 79608
rect 139578 79568 139584 79580
rect 139636 79568 139642 79620
rect 140056 79552 140084 79852
rect 140176 79840 140182 79892
rect 140234 79840 140240 79892
rect 140452 79840 140458 79892
rect 140510 79840 140516 79892
rect 139762 79540 139768 79552
rect 139320 79512 139768 79540
rect 136140 79500 136146 79512
rect 139762 79500 139768 79512
rect 139820 79500 139826 79552
rect 140038 79500 140044 79552
rect 140096 79500 140102 79552
rect 135530 79472 135536 79484
rect 135180 79444 135536 79472
rect 135530 79432 135536 79444
rect 135588 79432 135594 79484
rect 135714 79432 135720 79484
rect 135772 79432 135778 79484
rect 137002 79432 137008 79484
rect 137060 79472 137066 79484
rect 137922 79472 137928 79484
rect 137060 79444 137928 79472
rect 137060 79432 137066 79444
rect 137922 79432 137928 79444
rect 137980 79432 137986 79484
rect 140194 79404 140222 79840
rect 140314 79636 140320 79688
rect 140372 79676 140378 79688
rect 140470 79676 140498 79840
rect 140608 79824 140636 79908
rect 141022 79880 141050 79908
rect 140792 79852 141050 79880
rect 140590 79772 140596 79824
rect 140648 79772 140654 79824
rect 140372 79648 140498 79676
rect 140372 79636 140378 79648
rect 140792 79620 140820 79852
rect 141050 79704 141056 79756
rect 141108 79704 141114 79756
rect 141068 79676 141096 79704
rect 141160 79688 141188 79908
rect 141280 79840 141286 79892
rect 141338 79880 141344 79892
rect 141338 79840 141372 79880
rect 141464 79840 141470 79892
rect 141522 79840 141528 79892
rect 141648 79840 141654 79892
rect 141706 79840 141712 79892
rect 140976 79648 141096 79676
rect 140774 79568 140780 79620
rect 140832 79568 140838 79620
rect 140976 79540 141004 79648
rect 141142 79636 141148 79688
rect 141200 79636 141206 79688
rect 141050 79568 141056 79620
rect 141108 79608 141114 79620
rect 141344 79608 141372 79840
rect 141108 79580 141372 79608
rect 141108 79568 141114 79580
rect 141234 79540 141240 79552
rect 140976 79512 141240 79540
rect 141234 79500 141240 79512
rect 141292 79500 141298 79552
rect 141326 79500 141332 79552
rect 141384 79540 141390 79552
rect 141482 79540 141510 79840
rect 141384 79512 141510 79540
rect 141384 79500 141390 79512
rect 141510 79432 141516 79484
rect 141568 79472 141574 79484
rect 141666 79472 141694 79840
rect 141758 79540 141786 79920
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 141942 79948 141970 80260
rect 142126 80152 142154 80328
rect 142126 80124 143534 80152
rect 143506 80016 143534 80124
rect 143506 79988 144362 80016
rect 142384 79948 142390 79960
rect 141942 79920 142390 79948
rect 142384 79908 142390 79920
rect 142442 79908 142448 79960
rect 143396 79948 143402 79960
rect 142770 79920 143402 79948
rect 142476 79840 142482 79892
rect 142534 79840 142540 79892
rect 142770 79880 142798 79920
rect 143396 79908 143402 79920
rect 143454 79908 143460 79960
rect 143580 79908 143586 79960
rect 143638 79908 143644 79960
rect 142632 79852 142798 79880
rect 142200 79772 142206 79824
rect 142258 79772 142264 79824
rect 141970 79636 141976 79688
rect 142028 79676 142034 79688
rect 142218 79676 142246 79772
rect 142028 79648 142246 79676
rect 142028 79636 142034 79648
rect 142062 79540 142068 79552
rect 141758 79512 142068 79540
rect 142062 79500 142068 79512
rect 142120 79500 142126 79552
rect 142494 79540 142522 79840
rect 142632 79620 142660 79852
rect 142936 79840 142942 79892
rect 142994 79880 143000 79892
rect 142994 79840 143028 79880
rect 143212 79840 143218 79892
rect 143270 79840 143276 79892
rect 143488 79840 143494 79892
rect 143546 79840 143552 79892
rect 142752 79772 142758 79824
rect 142810 79772 142816 79824
rect 142770 79620 142798 79772
rect 142614 79568 142620 79620
rect 142672 79568 142678 79620
rect 142770 79580 142804 79620
rect 142798 79568 142804 79580
rect 142856 79568 142862 79620
rect 142890 79540 142896 79552
rect 142494 79512 142896 79540
rect 142890 79500 142896 79512
rect 142948 79500 142954 79552
rect 141568 79444 141694 79472
rect 141568 79432 141574 79444
rect 142522 79432 142528 79484
rect 142580 79472 142586 79484
rect 143000 79472 143028 79840
rect 143230 79484 143258 79840
rect 143506 79812 143534 79840
rect 143460 79784 143534 79812
rect 143460 79484 143488 79784
rect 143598 79756 143626 79908
rect 143672 79840 143678 79892
rect 143730 79840 143736 79892
rect 144132 79880 144138 79892
rect 143828 79852 144138 79880
rect 143534 79704 143540 79756
rect 143592 79716 143626 79756
rect 143592 79704 143598 79716
rect 142580 79444 143028 79472
rect 142580 79432 142586 79444
rect 143166 79432 143172 79484
rect 143224 79444 143258 79484
rect 143224 79432 143230 79444
rect 143442 79432 143448 79484
rect 143500 79432 143506 79484
rect 133018 79376 140222 79404
rect 141142 79364 141148 79416
rect 141200 79404 141206 79416
rect 141602 79404 141608 79416
rect 141200 79376 141608 79404
rect 141200 79364 141206 79376
rect 141602 79364 141608 79376
rect 141660 79364 141666 79416
rect 143690 79336 143718 79840
rect 143828 79688 143856 79852
rect 144132 79840 144138 79852
rect 144190 79840 144196 79892
rect 143948 79772 143954 79824
rect 144006 79772 144012 79824
rect 143966 79688 143994 79772
rect 143810 79636 143816 79688
rect 143868 79636 143874 79688
rect 143966 79648 144000 79688
rect 143994 79636 144000 79648
rect 144052 79636 144058 79688
rect 144334 79552 144362 79988
rect 144334 79512 144368 79552
rect 144362 79500 144368 79512
rect 144420 79500 144426 79552
rect 144472 79472 144500 80464
rect 144794 80016 144822 80668
rect 146726 80016 146754 80736
rect 150682 80152 150710 81212
rect 177960 81036 177988 81212
rect 177960 81008 178034 81036
rect 178006 80968 178034 81008
rect 187666 81008 193214 81036
rect 187666 80968 187694 81008
rect 150498 80124 150710 80152
rect 151878 80940 155954 80968
rect 178006 80940 187694 80968
rect 144794 79988 145236 80016
rect 146726 79988 149238 80016
rect 144776 79908 144782 79960
rect 144834 79908 144840 79960
rect 144868 79908 144874 79960
rect 144926 79908 144932 79960
rect 144592 79840 144598 79892
rect 144650 79840 144656 79892
rect 144610 79688 144638 79840
rect 144794 79824 144822 79908
rect 144886 79880 144914 79908
rect 145208 79880 145236 79988
rect 149210 79960 149238 79988
rect 145696 79908 145702 79960
rect 145754 79908 145760 79960
rect 145788 79908 145794 79960
rect 145846 79908 145852 79960
rect 145972 79908 145978 79960
rect 146030 79908 146036 79960
rect 146064 79908 146070 79960
rect 146122 79948 146128 79960
rect 146122 79908 146156 79948
rect 146248 79908 146254 79960
rect 146306 79948 146312 79960
rect 146306 79920 146662 79948
rect 146306 79908 146312 79920
rect 145512 79880 145518 79892
rect 144886 79852 144960 79880
rect 144794 79784 144828 79824
rect 144822 79772 144828 79784
rect 144880 79772 144886 79824
rect 144610 79648 144644 79688
rect 144638 79636 144644 79648
rect 144696 79636 144702 79688
rect 144546 79500 144552 79552
rect 144604 79540 144610 79552
rect 144932 79540 144960 79852
rect 145208 79852 145518 79880
rect 145208 79552 145236 79852
rect 145512 79840 145518 79852
rect 145570 79840 145576 79892
rect 145558 79704 145564 79756
rect 145616 79704 145622 79756
rect 144604 79512 144960 79540
rect 144604 79500 144610 79512
rect 145190 79500 145196 79552
rect 145248 79500 145254 79552
rect 145576 79540 145604 79704
rect 145714 79688 145742 79908
rect 145650 79636 145656 79688
rect 145708 79648 145742 79688
rect 145708 79636 145714 79648
rect 145650 79540 145656 79552
rect 145576 79512 145656 79540
rect 145650 79500 145656 79512
rect 145708 79500 145714 79552
rect 144472 79444 144592 79472
rect 144454 79336 144460 79348
rect 130436 79308 131160 79336
rect 131224 79308 144460 79336
rect 130436 79296 130442 79308
rect 123294 79228 123300 79280
rect 123352 79268 123358 79280
rect 131224 79268 131252 79308
rect 144454 79296 144460 79308
rect 144512 79296 144518 79348
rect 144564 79336 144592 79444
rect 145006 79432 145012 79484
rect 145064 79472 145070 79484
rect 145806 79472 145834 79908
rect 145990 79824 146018 79908
rect 146128 79824 146156 79908
rect 146340 79880 146346 79892
rect 146312 79840 146346 79880
rect 146398 79840 146404 79892
rect 146524 79840 146530 79892
rect 146582 79840 146588 79892
rect 145990 79784 146024 79824
rect 146018 79772 146024 79784
rect 146076 79772 146082 79824
rect 146110 79772 146116 79824
rect 146168 79772 146174 79824
rect 146312 79756 146340 79840
rect 146294 79704 146300 79756
rect 146352 79704 146358 79756
rect 146542 79620 146570 79840
rect 146634 79812 146662 79920
rect 146708 79908 146714 79960
rect 146766 79948 146772 79960
rect 146984 79948 146990 79960
rect 146766 79908 146800 79948
rect 146634 79784 146708 79812
rect 146680 79756 146708 79784
rect 146662 79704 146668 79756
rect 146720 79704 146726 79756
rect 146542 79580 146576 79620
rect 146570 79568 146576 79580
rect 146628 79568 146634 79620
rect 146772 79484 146800 79908
rect 146956 79908 146990 79948
rect 147042 79908 147048 79960
rect 147076 79908 147082 79960
rect 147134 79908 147140 79960
rect 147168 79908 147174 79960
rect 147226 79908 147232 79960
rect 147444 79908 147450 79960
rect 147502 79908 147508 79960
rect 147536 79908 147542 79960
rect 147594 79908 147600 79960
rect 147904 79908 147910 79960
rect 147962 79948 147968 79960
rect 147962 79908 147996 79948
rect 148088 79908 148094 79960
rect 148146 79948 148152 79960
rect 148824 79948 148830 79960
rect 148146 79920 148594 79948
rect 148146 79908 148152 79920
rect 146956 79756 146984 79908
rect 147094 79880 147122 79908
rect 147048 79852 147122 79880
rect 146938 79704 146944 79756
rect 146996 79704 147002 79756
rect 147048 79688 147076 79852
rect 147186 79812 147214 79908
rect 147140 79784 147214 79812
rect 147462 79812 147490 79908
rect 147554 79880 147582 79908
rect 147554 79852 147720 79880
rect 147462 79784 147628 79812
rect 147140 79688 147168 79784
rect 147214 79704 147220 79756
rect 147272 79744 147278 79756
rect 147490 79744 147496 79756
rect 147272 79716 147496 79744
rect 147272 79704 147278 79716
rect 147490 79704 147496 79716
rect 147548 79704 147554 79756
rect 147030 79636 147036 79688
rect 147088 79636 147094 79688
rect 147122 79636 147128 79688
rect 147180 79636 147186 79688
rect 147214 79568 147220 79620
rect 147272 79608 147278 79620
rect 147600 79608 147628 79784
rect 147272 79580 147628 79608
rect 147272 79568 147278 79580
rect 147398 79500 147404 79552
rect 147456 79540 147462 79552
rect 147582 79540 147588 79552
rect 147456 79512 147588 79540
rect 147456 79500 147462 79512
rect 147582 79500 147588 79512
rect 147640 79540 147646 79552
rect 147692 79540 147720 79852
rect 147812 79840 147818 79892
rect 147870 79880 147876 79892
rect 147870 79840 147904 79880
rect 147766 79704 147772 79756
rect 147824 79704 147830 79756
rect 147784 79620 147812 79704
rect 147876 79688 147904 79840
rect 147858 79636 147864 79688
rect 147916 79636 147922 79688
rect 147968 79620 147996 79908
rect 148272 79840 148278 79892
rect 148330 79840 148336 79892
rect 148364 79840 148370 79892
rect 148422 79840 148428 79892
rect 148290 79756 148318 79840
rect 148226 79704 148232 79756
rect 148284 79716 148318 79756
rect 148284 79704 148290 79716
rect 148382 79688 148410 79840
rect 148318 79636 148324 79688
rect 148376 79648 148410 79688
rect 148376 79636 148382 79648
rect 147766 79568 147772 79620
rect 147824 79568 147830 79620
rect 147950 79568 147956 79620
rect 148008 79568 148014 79620
rect 147640 79512 147720 79540
rect 147640 79500 147646 79512
rect 148566 79484 148594 79920
rect 148704 79920 148830 79948
rect 148704 79688 148732 79920
rect 148824 79908 148830 79920
rect 148882 79908 148888 79960
rect 148916 79908 148922 79960
rect 148974 79908 148980 79960
rect 149100 79908 149106 79960
rect 149158 79908 149164 79960
rect 149192 79908 149198 79960
rect 149250 79908 149256 79960
rect 149652 79948 149658 79960
rect 149394 79920 149658 79948
rect 148934 79880 148962 79908
rect 148796 79852 148962 79880
rect 148686 79636 148692 79688
rect 148744 79636 148750 79688
rect 145064 79444 145834 79472
rect 145064 79432 145070 79444
rect 146754 79432 146760 79484
rect 146812 79432 146818 79484
rect 148566 79444 148600 79484
rect 148594 79432 148600 79444
rect 148652 79432 148658 79484
rect 147398 79364 147404 79416
rect 147456 79404 147462 79416
rect 148796 79404 148824 79852
rect 149118 79824 149146 79908
rect 149210 79880 149238 79908
rect 149210 79852 149284 79880
rect 148870 79772 148876 79824
rect 148928 79772 148934 79824
rect 149118 79784 149152 79824
rect 149146 79772 149152 79784
rect 149204 79772 149210 79824
rect 148888 79676 148916 79772
rect 149054 79676 149060 79688
rect 148888 79648 149060 79676
rect 149054 79636 149060 79648
rect 149112 79636 149118 79688
rect 149256 79676 149284 79852
rect 149164 79648 149284 79676
rect 149164 79540 149192 79648
rect 149238 79568 149244 79620
rect 149296 79608 149302 79620
rect 149394 79608 149422 79920
rect 149652 79908 149658 79920
rect 149710 79908 149716 79960
rect 149744 79908 149750 79960
rect 149802 79908 149808 79960
rect 149836 79908 149842 79960
rect 149894 79908 149900 79960
rect 149468 79840 149474 79892
rect 149526 79840 149532 79892
rect 149486 79744 149514 79840
rect 149762 79824 149790 79908
rect 149854 79880 149882 79908
rect 149854 79852 149928 79880
rect 149698 79772 149704 79824
rect 149756 79784 149790 79824
rect 149756 79772 149762 79784
rect 149790 79744 149796 79756
rect 149486 79716 149796 79744
rect 149790 79704 149796 79716
rect 149848 79704 149854 79756
rect 149900 79688 149928 79852
rect 150112 79840 150118 79892
rect 150170 79840 150176 79892
rect 149882 79636 149888 79688
rect 149940 79636 149946 79688
rect 149296 79580 149422 79608
rect 150130 79608 150158 79840
rect 150498 79812 150526 80124
rect 151878 80084 151906 80940
rect 155926 80764 155954 80940
rect 187418 80860 187424 80912
rect 187476 80900 187482 80912
rect 188614 80900 188620 80912
rect 187476 80872 188620 80900
rect 187476 80860 187482 80872
rect 188614 80860 188620 80872
rect 188672 80860 188678 80912
rect 193186 80900 193214 81008
rect 206094 80900 206100 80912
rect 193186 80872 206100 80900
rect 206094 80860 206100 80872
rect 206152 80900 206158 80912
rect 234614 80900 234620 80912
rect 206152 80872 234620 80900
rect 206152 80860 206158 80872
rect 234614 80860 234620 80872
rect 234672 80860 234678 80912
rect 186774 80832 186780 80844
rect 158686 80804 178172 80832
rect 158686 80764 158714 80804
rect 155926 80736 158714 80764
rect 162734 80736 175090 80764
rect 162734 80492 162762 80736
rect 153350 80464 162762 80492
rect 162826 80668 174630 80696
rect 153350 80084 153378 80464
rect 162826 80424 162854 80668
rect 150590 80056 151906 80084
rect 152062 80056 153378 80084
rect 153442 80396 162854 80424
rect 167656 80600 172790 80628
rect 150590 79880 150618 80056
rect 152062 79960 152090 80056
rect 153442 79960 153470 80396
rect 154822 80328 155954 80356
rect 154822 79960 154850 80328
rect 155926 80288 155954 80328
rect 167656 80288 167684 80600
rect 155926 80260 167684 80288
rect 168852 80532 172698 80560
rect 168852 80220 168880 80532
rect 172670 80424 172698 80532
rect 172762 80492 172790 80600
rect 174602 80560 174630 80668
rect 175062 80628 175090 80736
rect 177960 80736 178080 80764
rect 177960 80708 177988 80736
rect 178052 80708 178080 80736
rect 177942 80656 177948 80708
rect 178000 80656 178006 80708
rect 178034 80656 178040 80708
rect 178092 80656 178098 80708
rect 178144 80696 178172 80804
rect 178696 80804 186780 80832
rect 178586 80696 178592 80708
rect 178144 80668 178592 80696
rect 178586 80656 178592 80668
rect 178644 80656 178650 80708
rect 178696 80628 178724 80804
rect 186774 80792 186780 80804
rect 186832 80832 186838 80844
rect 252554 80832 252560 80844
rect 186832 80804 252560 80832
rect 186832 80792 186838 80804
rect 252554 80792 252560 80804
rect 252612 80792 252618 80844
rect 188154 80764 188160 80776
rect 175062 80600 178724 80628
rect 180444 80736 188160 80764
rect 180444 80560 180472 80736
rect 188154 80724 188160 80736
rect 188212 80764 188218 80776
rect 270494 80764 270500 80776
rect 188212 80736 270500 80764
rect 188212 80724 188218 80736
rect 270494 80724 270500 80736
rect 270552 80724 270558 80776
rect 188614 80656 188620 80708
rect 188672 80696 188678 80708
rect 189258 80696 189264 80708
rect 188672 80668 189264 80696
rect 188672 80656 188678 80668
rect 189258 80656 189264 80668
rect 189316 80696 189322 80708
rect 288434 80696 288440 80708
rect 189316 80668 288440 80696
rect 189316 80656 189322 80668
rect 288434 80656 288440 80668
rect 288492 80656 288498 80708
rect 174602 80532 180472 80560
rect 187418 80492 187424 80504
rect 172762 80464 187424 80492
rect 187418 80452 187424 80464
rect 187476 80452 187482 80504
rect 172670 80396 179414 80424
rect 178770 80356 178776 80368
rect 155926 80192 168880 80220
rect 172762 80328 178776 80356
rect 150664 79908 150670 79960
rect 150722 79948 150728 79960
rect 150722 79920 151078 79948
rect 150722 79908 150728 79920
rect 150940 79880 150946 79892
rect 150590 79852 150946 79880
rect 150940 79840 150946 79852
rect 150998 79840 151004 79892
rect 151050 79812 151078 79920
rect 151216 79908 151222 79960
rect 151274 79908 151280 79960
rect 151400 79948 151406 79960
rect 151372 79908 151406 79948
rect 151458 79908 151464 79960
rect 152044 79908 152050 79960
rect 152102 79908 152108 79960
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 152872 79908 152878 79960
rect 152930 79908 152936 79960
rect 152964 79908 152970 79960
rect 153022 79908 153028 79960
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 154160 79948 154166 79960
rect 154132 79908 154166 79948
rect 154218 79908 154224 79960
rect 154252 79908 154258 79960
rect 154310 79908 154316 79960
rect 154344 79908 154350 79960
rect 154402 79908 154408 79960
rect 154436 79908 154442 79960
rect 154494 79948 154500 79960
rect 154494 79908 154528 79948
rect 154804 79908 154810 79960
rect 154862 79908 154868 79960
rect 154988 79908 154994 79960
rect 155046 79908 155052 79960
rect 155172 79908 155178 79960
rect 155230 79908 155236 79960
rect 151234 79824 151262 79908
rect 150498 79784 151078 79812
rect 151170 79772 151176 79824
rect 151228 79784 151262 79824
rect 151228 79772 151234 79784
rect 150342 79704 150348 79756
rect 150400 79704 150406 79756
rect 150360 79676 150388 79704
rect 151372 79688 151400 79908
rect 151860 79840 151866 79892
rect 151918 79840 151924 79892
rect 150434 79676 150440 79688
rect 150360 79648 150440 79676
rect 150434 79636 150440 79648
rect 150492 79636 150498 79688
rect 151354 79636 151360 79688
rect 151412 79636 151418 79688
rect 151878 79620 151906 79840
rect 152228 79772 152234 79824
rect 152286 79772 152292 79824
rect 152246 79688 152274 79772
rect 152182 79636 152188 79688
rect 152240 79648 152274 79688
rect 152240 79636 152246 79648
rect 150986 79608 150992 79620
rect 150130 79580 150992 79608
rect 149296 79568 149302 79580
rect 150986 79568 150992 79580
rect 151044 79568 151050 79620
rect 151814 79568 151820 79620
rect 151872 79580 151906 79620
rect 152430 79608 152458 79908
rect 152688 79880 152694 79892
rect 152660 79840 152694 79880
rect 152746 79840 152752 79892
rect 152660 79688 152688 79840
rect 152642 79636 152648 79688
rect 152700 79636 152706 79688
rect 152550 79608 152556 79620
rect 152430 79580 152556 79608
rect 151872 79568 151878 79580
rect 152550 79568 152556 79580
rect 152608 79568 152614 79620
rect 152890 79608 152918 79908
rect 152982 79824 153010 79908
rect 153148 79840 153154 79892
rect 153206 79840 153212 79892
rect 153700 79840 153706 79892
rect 153758 79880 153764 79892
rect 153758 79840 153792 79880
rect 152964 79772 152970 79824
rect 153022 79772 153028 79824
rect 153010 79636 153016 79688
rect 153068 79676 153074 79688
rect 153166 79676 153194 79840
rect 153068 79648 153194 79676
rect 153068 79636 153074 79648
rect 153764 79620 153792 79840
rect 153884 79812 153890 79824
rect 153856 79772 153890 79812
rect 153942 79772 153948 79824
rect 153286 79608 153292 79620
rect 152890 79580 153292 79608
rect 153286 79568 153292 79580
rect 153344 79568 153350 79620
rect 153746 79568 153752 79620
rect 153804 79568 153810 79620
rect 150158 79540 150164 79552
rect 149164 79512 150164 79540
rect 150158 79500 150164 79512
rect 150216 79500 150222 79552
rect 153470 79500 153476 79552
rect 153528 79540 153534 79552
rect 153856 79540 153884 79772
rect 154132 79744 154160 79908
rect 154270 79824 154298 79908
rect 154206 79772 154212 79824
rect 154264 79784 154298 79824
rect 154362 79824 154390 79908
rect 154362 79784 154396 79824
rect 154264 79772 154270 79784
rect 154390 79772 154396 79784
rect 154448 79772 154454 79824
rect 153948 79716 154160 79744
rect 153948 79620 153976 79716
rect 154298 79636 154304 79688
rect 154356 79676 154362 79688
rect 154500 79676 154528 79908
rect 154620 79840 154626 79892
rect 154678 79880 154684 79892
rect 154678 79840 154712 79880
rect 154684 79688 154712 79840
rect 154758 79704 154764 79756
rect 154816 79744 154822 79756
rect 155006 79744 155034 79908
rect 154816 79716 155034 79744
rect 154816 79704 154822 79716
rect 154356 79648 154528 79676
rect 154356 79636 154362 79648
rect 154666 79636 154672 79688
rect 154724 79636 154730 79688
rect 153930 79568 153936 79620
rect 153988 79568 153994 79620
rect 154942 79568 154948 79620
rect 155000 79608 155006 79620
rect 155190 79608 155218 79908
rect 155926 79892 155954 80192
rect 172762 80084 172790 80328
rect 178770 80316 178776 80328
rect 178828 80316 178834 80368
rect 179386 80288 179414 80396
rect 185210 80288 185216 80300
rect 179386 80260 185216 80288
rect 185210 80248 185216 80260
rect 185268 80248 185274 80300
rect 177758 80220 177764 80232
rect 168530 80056 172790 80084
rect 173038 80192 177764 80220
rect 156662 79988 156920 80016
rect 156276 79908 156282 79960
rect 156334 79908 156340 79960
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 156552 79908 156558 79960
rect 156610 79908 156616 79960
rect 155356 79880 155362 79892
rect 155000 79580 155218 79608
rect 155328 79840 155362 79880
rect 155414 79840 155420 79892
rect 155908 79840 155914 79892
rect 155966 79840 155972 79892
rect 156184 79840 156190 79892
rect 156242 79840 156248 79892
rect 155000 79568 155006 79580
rect 153528 79512 153884 79540
rect 153528 79500 153534 79512
rect 155126 79500 155132 79552
rect 155184 79540 155190 79552
rect 155328 79540 155356 79840
rect 155448 79772 155454 79824
rect 155506 79812 155512 79824
rect 155506 79772 155540 79812
rect 155512 79688 155540 79772
rect 155494 79636 155500 79688
rect 155552 79636 155558 79688
rect 156202 79552 156230 79840
rect 155184 79512 155356 79540
rect 155184 79500 155190 79512
rect 156138 79500 156144 79552
rect 156196 79512 156230 79552
rect 156196 79500 156202 79512
rect 156294 79484 156322 79908
rect 156230 79432 156236 79484
rect 156288 79444 156322 79484
rect 156386 79472 156414 79908
rect 156570 79744 156598 79908
rect 156524 79716 156598 79744
rect 156524 79608 156552 79716
rect 156662 79688 156690 79988
rect 156892 79960 156920 79988
rect 157674 79988 157886 80016
rect 157674 79960 157702 79988
rect 156736 79908 156742 79960
rect 156794 79908 156800 79960
rect 156892 79920 156926 79960
rect 156920 79908 156926 79920
rect 156978 79908 156984 79960
rect 157288 79908 157294 79960
rect 157346 79948 157352 79960
rect 157472 79948 157478 79960
rect 157346 79908 157380 79948
rect 156754 79756 156782 79908
rect 156828 79840 156834 79892
rect 156886 79880 156892 79892
rect 156886 79840 156920 79880
rect 156754 79716 156788 79756
rect 156782 79704 156788 79716
rect 156840 79704 156846 79756
rect 156892 79688 156920 79840
rect 156598 79636 156604 79688
rect 156656 79676 156690 79688
rect 156656 79648 156828 79676
rect 156656 79636 156662 79648
rect 156690 79608 156696 79620
rect 156524 79580 156696 79608
rect 156690 79568 156696 79580
rect 156748 79568 156754 79620
rect 156800 79608 156828 79648
rect 156874 79636 156880 79688
rect 156932 79636 156938 79688
rect 157242 79608 157248 79620
rect 156800 79580 157248 79608
rect 157242 79568 157248 79580
rect 157300 79568 157306 79620
rect 157058 79472 157064 79484
rect 156386 79444 157064 79472
rect 156288 79432 156294 79444
rect 157058 79432 157064 79444
rect 157116 79432 157122 79484
rect 147456 79376 148824 79404
rect 147456 79364 147462 79376
rect 152642 79336 152648 79348
rect 144564 79308 152648 79336
rect 152642 79296 152648 79308
rect 152700 79296 152706 79348
rect 156966 79296 156972 79348
rect 157024 79336 157030 79348
rect 157352 79336 157380 79908
rect 157444 79908 157478 79948
rect 157530 79908 157536 79960
rect 157564 79908 157570 79960
rect 157622 79908 157628 79960
rect 157656 79908 157662 79960
rect 157714 79908 157720 79960
rect 157748 79908 157754 79960
rect 157806 79908 157812 79960
rect 157444 79540 157472 79908
rect 157582 79880 157610 79908
rect 157536 79852 157610 79880
rect 157536 79688 157564 79852
rect 157766 79812 157794 79908
rect 157628 79784 157794 79812
rect 157518 79636 157524 79688
rect 157576 79636 157582 79688
rect 157518 79540 157524 79552
rect 157444 79512 157524 79540
rect 157518 79500 157524 79512
rect 157576 79500 157582 79552
rect 157024 79308 157380 79336
rect 157628 79336 157656 79784
rect 157858 79608 157886 79988
rect 158640 79988 158898 80016
rect 158208 79908 158214 79960
rect 158266 79948 158272 79960
rect 158266 79908 158300 79948
rect 158484 79908 158490 79960
rect 158542 79908 158548 79960
rect 158024 79840 158030 79892
rect 158082 79840 158088 79892
rect 157932 79772 157938 79824
rect 157990 79772 157996 79824
rect 157720 79580 157886 79608
rect 157720 79404 157748 79580
rect 157950 79552 157978 79772
rect 158042 79608 158070 79840
rect 158272 79688 158300 79908
rect 158392 79880 158398 79892
rect 158364 79840 158398 79880
rect 158450 79840 158456 79892
rect 158364 79688 158392 79840
rect 158502 79688 158530 79908
rect 158640 79688 158668 79988
rect 158870 79960 158898 79988
rect 160250 79988 160784 80016
rect 160250 79960 160278 79988
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 158852 79908 158858 79960
rect 158910 79908 158916 79960
rect 159036 79908 159042 79960
rect 159094 79948 159100 79960
rect 159094 79920 159266 79948
rect 159094 79908 159100 79920
rect 158778 79824 158806 79908
rect 159128 79880 159134 79892
rect 158916 79852 159134 79880
rect 158778 79784 158812 79824
rect 158806 79772 158812 79784
rect 158864 79772 158870 79824
rect 158916 79688 158944 79852
rect 159128 79840 159134 79852
rect 159186 79840 159192 79892
rect 159082 79704 159088 79756
rect 159140 79744 159146 79756
rect 159238 79744 159266 79920
rect 159588 79908 159594 79960
rect 159646 79908 159652 79960
rect 159680 79908 159686 79960
rect 159738 79948 159744 79960
rect 159738 79920 159864 79948
rect 159738 79908 159744 79920
rect 159496 79772 159502 79824
rect 159554 79772 159560 79824
rect 159140 79716 159266 79744
rect 159140 79704 159146 79716
rect 158254 79636 158260 79688
rect 158312 79636 158318 79688
rect 158346 79636 158352 79688
rect 158404 79636 158410 79688
rect 158502 79648 158536 79688
rect 158530 79636 158536 79648
rect 158588 79636 158594 79688
rect 158622 79636 158628 79688
rect 158680 79636 158686 79688
rect 158898 79636 158904 79688
rect 158956 79636 158962 79688
rect 159514 79620 159542 79772
rect 159606 79688 159634 79908
rect 159606 79648 159640 79688
rect 159634 79636 159640 79648
rect 159692 79636 159698 79688
rect 158438 79608 158444 79620
rect 158042 79580 158444 79608
rect 158438 79568 158444 79580
rect 158496 79568 158502 79620
rect 159514 79580 159548 79620
rect 159542 79568 159548 79580
rect 159600 79568 159606 79620
rect 159836 79552 159864 79920
rect 160048 79908 160054 79960
rect 160106 79908 160112 79960
rect 160232 79908 160238 79960
rect 160290 79908 160296 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 160066 79688 160094 79908
rect 160140 79840 160146 79892
rect 160198 79840 160204 79892
rect 160324 79840 160330 79892
rect 160382 79840 160388 79892
rect 160002 79636 160008 79688
rect 160060 79648 160094 79688
rect 160060 79636 160066 79648
rect 160158 79620 160186 79840
rect 160342 79756 160370 79840
rect 160278 79704 160284 79756
rect 160336 79716 160370 79756
rect 160336 79704 160342 79716
rect 160434 79676 160462 79908
rect 160618 79880 160646 79908
rect 160618 79852 160692 79880
rect 160554 79676 160560 79688
rect 160434 79648 160560 79676
rect 160554 79636 160560 79648
rect 160612 79636 160618 79688
rect 160094 79568 160100 79620
rect 160152 79580 160186 79620
rect 160152 79568 160158 79580
rect 160370 79568 160376 79620
rect 160428 79608 160434 79620
rect 160664 79608 160692 79852
rect 160756 79620 160784 79988
rect 162274 79988 162670 80016
rect 162274 79960 162302 79988
rect 160876 79908 160882 79960
rect 160934 79908 160940 79960
rect 160968 79908 160974 79960
rect 161026 79948 161032 79960
rect 161026 79908 161060 79948
rect 161152 79908 161158 79960
rect 161210 79908 161216 79960
rect 161704 79908 161710 79960
rect 161762 79908 161768 79960
rect 161980 79948 161986 79960
rect 161814 79920 161986 79948
rect 160428 79580 160692 79608
rect 160428 79568 160434 79580
rect 160738 79568 160744 79620
rect 160796 79568 160802 79620
rect 160894 79552 160922 79908
rect 161032 79688 161060 79908
rect 161170 79824 161198 79908
rect 161336 79840 161342 79892
rect 161394 79840 161400 79892
rect 161170 79784 161204 79824
rect 161198 79772 161204 79784
rect 161256 79772 161262 79824
rect 161354 79756 161382 79840
rect 161722 79824 161750 79908
rect 161658 79772 161664 79824
rect 161716 79784 161750 79824
rect 161716 79772 161722 79784
rect 161290 79704 161296 79756
rect 161348 79716 161382 79756
rect 161348 79704 161354 79716
rect 161014 79636 161020 79688
rect 161072 79636 161078 79688
rect 161814 79608 161842 79920
rect 161980 79908 161986 79920
rect 162038 79908 162044 79960
rect 162072 79908 162078 79960
rect 162130 79908 162136 79960
rect 162256 79908 162262 79960
rect 162314 79908 162320 79960
rect 161888 79840 161894 79892
rect 161946 79880 161952 79892
rect 162090 79880 162118 79908
rect 162532 79880 162538 79892
rect 161946 79840 161980 79880
rect 162090 79852 162256 79880
rect 161952 79688 161980 79840
rect 161934 79636 161940 79688
rect 161992 79636 161998 79688
rect 162026 79608 162032 79620
rect 161814 79580 162032 79608
rect 162026 79568 162032 79580
rect 162084 79568 162090 79620
rect 157886 79500 157892 79552
rect 157944 79512 157978 79552
rect 157944 79500 157950 79512
rect 159818 79500 159824 79552
rect 159876 79500 159882 79552
rect 160830 79500 160836 79552
rect 160888 79512 160922 79552
rect 160888 79500 160894 79512
rect 162118 79500 162124 79552
rect 162176 79540 162182 79552
rect 162228 79540 162256 79852
rect 162504 79840 162538 79880
rect 162590 79840 162596 79892
rect 162504 79552 162532 79840
rect 162642 79812 162670 79988
rect 164804 79988 166166 80016
rect 163268 79908 163274 79960
rect 163326 79908 163332 79960
rect 163452 79908 163458 79960
rect 163510 79908 163516 79960
rect 163820 79908 163826 79960
rect 163878 79948 163884 79960
rect 163878 79908 163912 79948
rect 162808 79840 162814 79892
rect 162866 79880 162872 79892
rect 162866 79840 162900 79880
rect 162992 79840 162998 79892
rect 163050 79840 163056 79892
rect 163176 79840 163182 79892
rect 163234 79840 163240 79892
rect 162596 79784 162670 79812
rect 162596 79688 162624 79784
rect 162872 79688 162900 79840
rect 162578 79636 162584 79688
rect 162636 79636 162642 79688
rect 162854 79636 162860 79688
rect 162912 79636 162918 79688
rect 162176 79512 162256 79540
rect 162176 79500 162182 79512
rect 162486 79500 162492 79552
rect 162544 79500 162550 79552
rect 163010 79484 163038 79840
rect 163194 79688 163222 79840
rect 163130 79636 163136 79688
rect 163188 79648 163222 79688
rect 163188 79636 163194 79648
rect 163130 79500 163136 79552
rect 163188 79540 163194 79552
rect 163286 79540 163314 79908
rect 163360 79840 163366 79892
rect 163418 79840 163424 79892
rect 163188 79512 163314 79540
rect 163188 79500 163194 79512
rect 157794 79432 157800 79484
rect 157852 79472 157858 79484
rect 158162 79472 158168 79484
rect 157852 79444 158168 79472
rect 157852 79432 157858 79444
rect 158162 79432 158168 79444
rect 158220 79432 158226 79484
rect 162946 79432 162952 79484
rect 163004 79444 163038 79484
rect 163004 79432 163010 79444
rect 157978 79404 157984 79416
rect 157720 79376 157984 79404
rect 157978 79364 157984 79376
rect 158036 79364 158042 79416
rect 158070 79364 158076 79416
rect 158128 79404 158134 79416
rect 162394 79404 162400 79416
rect 158128 79376 162400 79404
rect 158128 79364 158134 79376
rect 162394 79364 162400 79376
rect 162452 79364 162458 79416
rect 162762 79364 162768 79416
rect 162820 79404 162826 79416
rect 163378 79404 163406 79840
rect 163470 79540 163498 79908
rect 163728 79840 163734 79892
rect 163786 79840 163792 79892
rect 163636 79812 163642 79824
rect 163608 79772 163642 79812
rect 163694 79772 163700 79824
rect 163608 79620 163636 79772
rect 163746 79756 163774 79840
rect 163746 79716 163780 79756
rect 163774 79704 163780 79716
rect 163832 79704 163838 79756
rect 163590 79568 163596 79620
rect 163648 79568 163654 79620
rect 163682 79540 163688 79552
rect 163470 79512 163688 79540
rect 163682 79500 163688 79512
rect 163740 79500 163746 79552
rect 163498 79432 163504 79484
rect 163556 79472 163562 79484
rect 163884 79472 163912 79908
rect 164096 79880 164102 79892
rect 164068 79840 164102 79880
rect 164154 79840 164160 79892
rect 164464 79840 164470 79892
rect 164522 79840 164528 79892
rect 164068 79552 164096 79840
rect 164372 79812 164378 79824
rect 164160 79784 164378 79812
rect 164160 79756 164188 79784
rect 164372 79772 164378 79784
rect 164430 79772 164436 79824
rect 164142 79704 164148 79756
rect 164200 79704 164206 79756
rect 164482 79688 164510 79840
rect 164648 79772 164654 79824
rect 164706 79772 164712 79824
rect 164666 79688 164694 79772
rect 164418 79636 164424 79688
rect 164476 79648 164510 79688
rect 164476 79636 164482 79648
rect 164602 79636 164608 79688
rect 164660 79648 164694 79688
rect 164660 79636 164666 79648
rect 164804 79552 164832 79988
rect 166138 79960 166166 79988
rect 166230 79988 166442 80016
rect 165016 79908 165022 79960
rect 165074 79908 165080 79960
rect 165108 79908 165114 79960
rect 165166 79948 165172 79960
rect 165166 79920 165660 79948
rect 165166 79908 165172 79920
rect 164050 79500 164056 79552
rect 164108 79500 164114 79552
rect 164786 79500 164792 79552
rect 164844 79500 164850 79552
rect 165034 79540 165062 79908
rect 165292 79840 165298 79892
rect 165350 79840 165356 79892
rect 165200 79772 165206 79824
rect 165258 79772 165264 79824
rect 165218 79688 165246 79772
rect 165154 79636 165160 79688
rect 165212 79648 165246 79688
rect 165212 79636 165218 79648
rect 165310 79620 165338 79840
rect 165246 79568 165252 79620
rect 165304 79580 165338 79620
rect 165304 79568 165310 79580
rect 165632 79552 165660 79920
rect 165936 79908 165942 79960
rect 165994 79908 166000 79960
rect 166120 79908 166126 79960
rect 166178 79908 166184 79960
rect 165954 79824 165982 79908
rect 166028 79840 166034 79892
rect 166086 79840 166092 79892
rect 166230 79880 166258 79988
rect 166414 79960 166442 79988
rect 168530 79960 168558 80056
rect 168806 79988 169294 80016
rect 168806 79960 168834 79988
rect 166396 79908 166402 79960
rect 166454 79908 166460 79960
rect 166488 79908 166494 79960
rect 166546 79908 166552 79960
rect 166764 79908 166770 79960
rect 166822 79908 166828 79960
rect 167224 79948 167230 79960
rect 167058 79920 167230 79948
rect 166230 79852 166350 79880
rect 165752 79772 165758 79824
rect 165810 79772 165816 79824
rect 165890 79772 165896 79824
rect 165948 79784 165982 79824
rect 165948 79772 165954 79784
rect 165770 79620 165798 79772
rect 165770 79580 165804 79620
rect 165798 79568 165804 79580
rect 165856 79568 165862 79620
rect 165430 79540 165436 79552
rect 165034 79512 165436 79540
rect 165430 79500 165436 79512
rect 165488 79500 165494 79552
rect 165614 79500 165620 79552
rect 165672 79500 165678 79552
rect 163556 79444 163912 79472
rect 166046 79472 166074 79840
rect 166322 79676 166350 79852
rect 166506 79812 166534 79908
rect 166506 79784 166580 79812
rect 166442 79676 166448 79688
rect 166322 79648 166448 79676
rect 166442 79636 166448 79648
rect 166500 79636 166506 79688
rect 166350 79568 166356 79620
rect 166408 79608 166414 79620
rect 166552 79608 166580 79784
rect 166408 79580 166580 79608
rect 166782 79620 166810 79908
rect 166856 79840 166862 79892
rect 166914 79880 166920 79892
rect 166914 79840 166948 79880
rect 166782 79580 166816 79620
rect 166408 79568 166414 79580
rect 166810 79568 166816 79580
rect 166868 79568 166874 79620
rect 166920 79540 166948 79840
rect 167058 79620 167086 79920
rect 167224 79908 167230 79920
rect 167282 79908 167288 79960
rect 167500 79908 167506 79960
rect 167558 79908 167564 79960
rect 167868 79908 167874 79960
rect 167926 79908 167932 79960
rect 167960 79908 167966 79960
rect 168018 79948 168024 79960
rect 168018 79920 168328 79948
rect 168018 79908 168024 79920
rect 167132 79840 167138 79892
rect 167190 79840 167196 79892
rect 167408 79840 167414 79892
rect 167466 79840 167472 79892
rect 167518 79880 167546 79908
rect 167518 79852 167684 79880
rect 167150 79812 167178 79840
rect 167426 79812 167454 79840
rect 167150 79784 167316 79812
rect 167426 79784 167500 79812
rect 167058 79580 167092 79620
rect 167086 79568 167092 79580
rect 167144 79568 167150 79620
rect 167178 79540 167184 79552
rect 166920 79512 167184 79540
rect 167178 79500 167184 79512
rect 167236 79500 167242 79552
rect 166534 79472 166540 79484
rect 166046 79444 166540 79472
rect 163556 79432 163562 79444
rect 166534 79432 166540 79444
rect 166592 79432 166598 79484
rect 167288 79472 167316 79784
rect 167472 79756 167500 79784
rect 167454 79704 167460 79756
rect 167512 79704 167518 79756
rect 167656 79688 167684 79852
rect 167776 79840 167782 79892
rect 167834 79840 167840 79892
rect 167794 79756 167822 79840
rect 167886 79824 167914 79908
rect 167886 79784 167920 79824
rect 167914 79772 167920 79784
rect 167972 79772 167978 79824
rect 167794 79716 167828 79756
rect 167822 79704 167828 79716
rect 167880 79704 167886 79756
rect 168300 79688 168328 79920
rect 168512 79908 168518 79960
rect 168570 79908 168576 79960
rect 168788 79908 168794 79960
rect 168846 79908 168852 79960
rect 169064 79948 169070 79960
rect 169036 79908 169070 79948
rect 169122 79908 169128 79960
rect 167638 79636 167644 79688
rect 167696 79636 167702 79688
rect 168282 79636 168288 79688
rect 168340 79636 168346 79688
rect 169036 79620 169064 79908
rect 169018 79568 169024 79620
rect 169076 79568 169082 79620
rect 169266 79608 169294 79988
rect 170646 79988 170950 80016
rect 169340 79908 169346 79960
rect 169398 79948 169404 79960
rect 169398 79908 169432 79948
rect 169524 79908 169530 79960
rect 169582 79908 169588 79960
rect 169708 79908 169714 79960
rect 169766 79908 169772 79960
rect 170260 79908 170266 79960
rect 170318 79908 170324 79960
rect 170352 79908 170358 79960
rect 170410 79908 170416 79960
rect 169404 79688 169432 79908
rect 169542 79688 169570 79908
rect 169616 79840 169622 79892
rect 169674 79840 169680 79892
rect 169386 79636 169392 79688
rect 169444 79636 169450 79688
rect 169478 79636 169484 79688
rect 169536 79648 169570 79688
rect 169536 79636 169542 79648
rect 169634 79620 169662 79840
rect 169266 79580 169432 79608
rect 169404 79552 169432 79580
rect 169570 79568 169576 79620
rect 169628 79580 169662 79620
rect 169726 79608 169754 79908
rect 169892 79840 169898 79892
rect 169950 79880 169956 79892
rect 169950 79840 169984 79880
rect 170168 79840 170174 79892
rect 170226 79840 170232 79892
rect 169846 79608 169852 79620
rect 169726 79580 169852 79608
rect 169628 79568 169634 79580
rect 169846 79568 169852 79580
rect 169904 79568 169910 79620
rect 169386 79500 169392 79552
rect 169444 79500 169450 79552
rect 169956 79540 169984 79840
rect 170186 79756 170214 79840
rect 170122 79744 170128 79756
rect 169772 79512 169984 79540
rect 170048 79716 170128 79744
rect 169772 79484 169800 79512
rect 168742 79472 168748 79484
rect 167288 79444 168748 79472
rect 168742 79432 168748 79444
rect 168800 79432 168806 79484
rect 169754 79432 169760 79484
rect 169812 79432 169818 79484
rect 170048 79472 170076 79716
rect 170122 79704 170128 79716
rect 170180 79716 170214 79756
rect 170180 79704 170186 79716
rect 170278 79608 170306 79908
rect 170370 79824 170398 79908
rect 170646 79880 170674 79988
rect 170922 79960 170950 79988
rect 173038 79960 173066 80192
rect 177758 80180 177764 80192
rect 177816 80180 177822 80232
rect 177850 80180 177856 80232
rect 177908 80220 177914 80232
rect 178402 80220 178408 80232
rect 177908 80192 178408 80220
rect 177908 80180 177914 80192
rect 178402 80180 178408 80192
rect 178460 80180 178466 80232
rect 178586 80180 178592 80232
rect 178644 80220 178650 80232
rect 182542 80220 182548 80232
rect 178644 80192 182548 80220
rect 178644 80180 178650 80192
rect 182542 80180 182548 80192
rect 182600 80220 182606 80232
rect 238754 80220 238760 80232
rect 182600 80192 238760 80220
rect 182600 80180 182606 80192
rect 238754 80180 238760 80192
rect 238812 80180 238818 80232
rect 178310 80152 178316 80164
rect 173498 80124 178316 80152
rect 170720 79908 170726 79960
rect 170778 79908 170784 79960
rect 170812 79908 170818 79960
rect 170870 79908 170876 79960
rect 170904 79908 170910 79960
rect 170962 79908 170968 79960
rect 171824 79948 171830 79960
rect 171796 79908 171830 79948
rect 171882 79908 171888 79960
rect 172192 79908 172198 79960
rect 172250 79908 172256 79960
rect 172468 79908 172474 79960
rect 172526 79908 172532 79960
rect 173020 79908 173026 79960
rect 173078 79908 173084 79960
rect 170508 79852 170674 79880
rect 170370 79784 170404 79824
rect 170398 79772 170404 79784
rect 170456 79772 170462 79824
rect 170140 79580 170306 79608
rect 170140 79552 170168 79580
rect 170508 79552 170536 79852
rect 170628 79772 170634 79824
rect 170686 79772 170692 79824
rect 170646 79676 170674 79772
rect 170600 79648 170674 79676
rect 170600 79552 170628 79648
rect 170122 79500 170128 79552
rect 170180 79500 170186 79552
rect 170490 79500 170496 79552
rect 170548 79500 170554 79552
rect 170582 79500 170588 79552
rect 170640 79500 170646 79552
rect 170738 79540 170766 79908
rect 170830 79608 170858 79908
rect 171272 79840 171278 79892
rect 171330 79880 171336 79892
rect 171330 79852 171548 79880
rect 171330 79840 171336 79852
rect 171088 79772 171094 79824
rect 171146 79772 171152 79824
rect 171106 79676 171134 79772
rect 171520 79688 171548 79852
rect 171640 79840 171646 79892
rect 171698 79840 171704 79892
rect 171106 79648 171272 79676
rect 171134 79608 171140 79620
rect 170830 79580 171140 79608
rect 171134 79568 171140 79580
rect 171192 79568 171198 79620
rect 170950 79540 170956 79552
rect 170738 79512 170956 79540
rect 170950 79500 170956 79512
rect 171008 79500 171014 79552
rect 171042 79472 171048 79484
rect 170048 79444 171048 79472
rect 171042 79432 171048 79444
rect 171100 79432 171106 79484
rect 162820 79376 163406 79404
rect 162820 79364 162826 79376
rect 157702 79336 157708 79348
rect 157628 79308 157708 79336
rect 157024 79296 157030 79308
rect 157702 79296 157708 79308
rect 157760 79296 157766 79348
rect 158438 79296 158444 79348
rect 158496 79336 158502 79348
rect 164970 79336 164976 79348
rect 158496 79308 164976 79336
rect 158496 79296 158502 79308
rect 164970 79296 164976 79308
rect 165028 79296 165034 79348
rect 171244 79336 171272 79648
rect 171502 79636 171508 79688
rect 171560 79636 171566 79688
rect 171658 79472 171686 79840
rect 171796 79620 171824 79908
rect 172210 79744 172238 79908
rect 172284 79840 172290 79892
rect 172342 79880 172348 79892
rect 172342 79840 172376 79880
rect 172072 79716 172238 79744
rect 172072 79688 172100 79716
rect 172348 79688 172376 79840
rect 172486 79824 172514 79908
rect 172836 79840 172842 79892
rect 172894 79840 172900 79892
rect 172928 79840 172934 79892
rect 172986 79880 172992 79892
rect 173112 79880 173118 79892
rect 172986 79840 173020 79880
rect 172422 79772 172428 79824
rect 172480 79784 172514 79824
rect 172480 79772 172486 79784
rect 172652 79772 172658 79824
rect 172710 79772 172716 79824
rect 172670 79688 172698 79772
rect 172854 79688 172882 79840
rect 172992 79756 173020 79840
rect 173084 79840 173118 79880
rect 173170 79840 173176 79892
rect 173204 79840 173210 79892
rect 173262 79880 173268 79892
rect 173262 79840 173296 79880
rect 173084 79756 173112 79840
rect 172974 79704 172980 79756
rect 173032 79704 173038 79756
rect 173066 79704 173072 79756
rect 173124 79704 173130 79756
rect 173158 79704 173164 79756
rect 173216 79704 173222 79756
rect 172054 79636 172060 79688
rect 172112 79636 172118 79688
rect 172330 79636 172336 79688
rect 172388 79636 172394 79688
rect 172670 79648 172704 79688
rect 172698 79636 172704 79648
rect 172756 79636 172762 79688
rect 172854 79648 172888 79688
rect 172882 79636 172888 79648
rect 172940 79636 172946 79688
rect 173176 79620 173204 79704
rect 173268 79620 173296 79840
rect 173388 79812 173394 79824
rect 173360 79772 173394 79812
rect 173446 79772 173452 79824
rect 173360 79620 173388 79772
rect 171778 79568 171784 79620
rect 171836 79568 171842 79620
rect 173158 79568 173164 79620
rect 173216 79568 173222 79620
rect 173250 79568 173256 79620
rect 173308 79568 173314 79620
rect 173342 79568 173348 79620
rect 173400 79568 173406 79620
rect 171870 79500 171876 79552
rect 171928 79540 171934 79552
rect 173498 79540 173526 80124
rect 178310 80112 178316 80124
rect 178368 80112 178374 80164
rect 178420 80084 178448 80180
rect 185210 80112 185216 80164
rect 185268 80152 185274 80164
rect 302234 80152 302240 80164
rect 185268 80124 302240 80152
rect 185268 80112 185274 80124
rect 302234 80112 302240 80124
rect 302292 80112 302298 80164
rect 380894 80084 380900 80096
rect 178420 80056 380900 80084
rect 380894 80044 380900 80056
rect 380952 80044 380958 80096
rect 178586 80016 178592 80028
rect 173866 79988 178592 80016
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 171928 79512 173526 79540
rect 171928 79500 171934 79512
rect 172790 79472 172796 79484
rect 171658 79444 172796 79472
rect 172790 79432 172796 79444
rect 172848 79432 172854 79484
rect 173434 79432 173440 79484
rect 173492 79472 173498 79484
rect 173590 79472 173618 79908
rect 173664 79840 173670 79892
rect 173722 79880 173728 79892
rect 173722 79840 173756 79880
rect 173728 79756 173756 79840
rect 173710 79704 173716 79756
rect 173768 79704 173774 79756
rect 173866 79608 173894 79988
rect 178586 79976 178592 79988
rect 178644 79976 178650 80028
rect 174032 79908 174038 79960
rect 174090 79908 174096 79960
rect 174308 79908 174314 79960
rect 174366 79908 174372 79960
rect 174400 79908 174406 79960
rect 174458 79908 174464 79960
rect 174768 79908 174774 79960
rect 174826 79908 174832 79960
rect 175044 79908 175050 79960
rect 175102 79948 175108 79960
rect 175102 79908 175136 79948
rect 175228 79908 175234 79960
rect 175286 79908 175292 79960
rect 175412 79908 175418 79960
rect 175470 79908 175476 79960
rect 175504 79908 175510 79960
rect 175562 79948 175568 79960
rect 175562 79908 175596 79948
rect 175780 79908 175786 79960
rect 175838 79908 175844 79960
rect 175964 79948 175970 79960
rect 175936 79908 175970 79948
rect 176022 79908 176028 79960
rect 176056 79908 176062 79960
rect 176114 79908 176120 79960
rect 177666 79908 177672 79960
rect 177724 79948 177730 79960
rect 177850 79948 177856 79960
rect 177724 79920 177856 79948
rect 177724 79908 177730 79920
rect 177850 79908 177856 79920
rect 177908 79908 177914 79960
rect 174050 79880 174078 79908
rect 174050 79852 174262 79880
rect 173940 79772 173946 79824
rect 173998 79812 174004 79824
rect 173998 79772 174032 79812
rect 174004 79688 174032 79772
rect 173986 79636 173992 79688
rect 174044 79636 174050 79688
rect 174078 79608 174084 79620
rect 173866 79580 174084 79608
rect 174078 79568 174084 79580
rect 174136 79568 174142 79620
rect 174234 79540 174262 79852
rect 174326 79756 174354 79908
rect 174418 79812 174446 79908
rect 174584 79840 174590 79892
rect 174642 79840 174648 79892
rect 174418 79784 174492 79812
rect 174464 79756 174492 79784
rect 174602 79756 174630 79840
rect 174786 79824 174814 79908
rect 174722 79772 174728 79824
rect 174780 79784 174814 79824
rect 174780 79772 174786 79784
rect 174326 79716 174360 79756
rect 174354 79704 174360 79716
rect 174412 79704 174418 79756
rect 174446 79704 174452 79756
rect 174504 79704 174510 79756
rect 174538 79704 174544 79756
rect 174596 79716 174630 79756
rect 174596 79704 174602 79716
rect 174814 79636 174820 79688
rect 174872 79676 174878 79688
rect 174872 79648 175044 79676
rect 174872 79636 174878 79648
rect 175016 79620 175044 79648
rect 174998 79568 175004 79620
rect 175056 79568 175062 79620
rect 174814 79540 174820 79552
rect 174234 79512 174820 79540
rect 174814 79500 174820 79512
rect 174872 79500 174878 79552
rect 175108 79540 175136 79908
rect 175246 79744 175274 79908
rect 175430 79880 175458 79908
rect 175430 79852 175504 79880
rect 175476 79756 175504 79852
rect 175246 79716 175412 79744
rect 175182 79568 175188 79620
rect 175240 79608 175246 79620
rect 175384 79608 175412 79716
rect 175458 79704 175464 79756
rect 175516 79704 175522 79756
rect 175240 79580 175412 79608
rect 175240 79568 175246 79580
rect 175274 79540 175280 79552
rect 175108 79512 175280 79540
rect 175274 79500 175280 79512
rect 175332 79500 175338 79552
rect 175568 79540 175596 79908
rect 175688 79880 175694 79892
rect 175660 79840 175694 79880
rect 175746 79840 175752 79892
rect 175660 79620 175688 79840
rect 175798 79756 175826 79908
rect 175734 79704 175740 79756
rect 175792 79716 175826 79756
rect 175792 79704 175798 79716
rect 175936 79676 175964 79908
rect 176074 79824 176102 79908
rect 176240 79840 176246 79892
rect 176298 79880 176304 79892
rect 176516 79880 176522 79892
rect 176298 79852 176424 79880
rect 176298 79840 176304 79852
rect 176010 79772 176016 79824
rect 176068 79784 176102 79824
rect 176068 79772 176074 79784
rect 176010 79676 176016 79688
rect 175936 79648 176016 79676
rect 176010 79636 176016 79648
rect 176068 79636 176074 79688
rect 176396 79620 176424 79852
rect 176488 79840 176522 79880
rect 176574 79840 176580 79892
rect 176792 79840 176798 79892
rect 176850 79840 176856 79892
rect 176884 79840 176890 79892
rect 176942 79840 176948 79892
rect 177068 79840 177074 79892
rect 177126 79840 177132 79892
rect 175642 79568 175648 79620
rect 175700 79568 175706 79620
rect 176378 79568 176384 79620
rect 176436 79568 176442 79620
rect 175568 79512 175826 79540
rect 173492 79444 173618 79472
rect 175798 79472 175826 79512
rect 175918 79500 175924 79552
rect 175976 79540 175982 79552
rect 176488 79540 176516 79840
rect 176608 79772 176614 79824
rect 176666 79772 176672 79824
rect 176626 79620 176654 79772
rect 176562 79568 176568 79620
rect 176620 79580 176654 79620
rect 176810 79608 176838 79840
rect 176902 79688 176930 79840
rect 177086 79688 177114 79840
rect 176902 79648 176936 79688
rect 176930 79636 176936 79648
rect 176988 79636 176994 79688
rect 177022 79636 177028 79688
rect 177080 79648 177114 79688
rect 177080 79636 177086 79648
rect 177114 79608 177120 79620
rect 176810 79580 177120 79608
rect 176620 79568 176626 79580
rect 177114 79568 177120 79580
rect 177172 79568 177178 79620
rect 175976 79512 176516 79540
rect 175976 79500 175982 79512
rect 176102 79472 176108 79484
rect 175798 79444 176108 79472
rect 173492 79432 173498 79444
rect 176102 79432 176108 79444
rect 176160 79432 176166 79484
rect 176286 79432 176292 79484
rect 176344 79472 176350 79484
rect 182174 79472 182180 79484
rect 176344 79444 182180 79472
rect 176344 79432 176350 79444
rect 182174 79432 182180 79444
rect 182232 79432 182238 79484
rect 171778 79364 171784 79416
rect 171836 79404 171842 79416
rect 174170 79404 174176 79416
rect 171836 79376 174176 79404
rect 171836 79364 171842 79376
rect 174170 79364 174176 79376
rect 174228 79364 174234 79416
rect 174354 79364 174360 79416
rect 174412 79404 174418 79416
rect 174814 79404 174820 79416
rect 174412 79376 174820 79404
rect 174412 79364 174418 79376
rect 174814 79364 174820 79376
rect 174872 79364 174878 79416
rect 175274 79364 175280 79416
rect 175332 79404 175338 79416
rect 178126 79404 178132 79416
rect 175332 79376 178132 79404
rect 175332 79364 175338 79376
rect 178126 79364 178132 79376
rect 178184 79364 178190 79416
rect 178310 79364 178316 79416
rect 178368 79404 178374 79416
rect 194318 79404 194324 79416
rect 178368 79376 194324 79404
rect 178368 79364 178374 79376
rect 194318 79364 194324 79376
rect 194376 79364 194382 79416
rect 172146 79336 172152 79348
rect 171244 79308 172152 79336
rect 172146 79296 172152 79308
rect 172204 79296 172210 79348
rect 175090 79296 175096 79348
rect 175148 79336 175154 79348
rect 177482 79336 177488 79348
rect 175148 79308 177488 79336
rect 175148 79296 175154 79308
rect 177482 79296 177488 79308
rect 177540 79296 177546 79348
rect 177758 79296 177764 79348
rect 177816 79336 177822 79348
rect 196802 79336 196808 79348
rect 177816 79308 196808 79336
rect 177816 79296 177822 79308
rect 196802 79296 196808 79308
rect 196860 79296 196866 79348
rect 525794 79336 525800 79348
rect 200086 79308 525800 79336
rect 123352 79240 131252 79268
rect 123352 79228 123358 79240
rect 132402 79228 132408 79280
rect 132460 79268 132466 79280
rect 147122 79268 147128 79280
rect 132460 79240 147128 79268
rect 132460 79228 132466 79240
rect 147122 79228 147128 79240
rect 147180 79228 147186 79280
rect 147950 79228 147956 79280
rect 148008 79268 148014 79280
rect 148008 79240 154712 79268
rect 148008 79228 148014 79240
rect 122466 79160 122472 79212
rect 122524 79200 122530 79212
rect 147674 79200 147680 79212
rect 122524 79172 147680 79200
rect 122524 79160 122530 79172
rect 147674 79160 147680 79172
rect 147732 79200 147738 79212
rect 148226 79200 148232 79212
rect 147732 79172 148232 79200
rect 147732 79160 147738 79172
rect 148226 79160 148232 79172
rect 148284 79160 148290 79212
rect 151906 79160 151912 79212
rect 151964 79200 151970 79212
rect 152274 79200 152280 79212
rect 151964 79172 152280 79200
rect 151964 79160 151970 79172
rect 152274 79160 152280 79172
rect 152332 79160 152338 79212
rect 154684 79200 154712 79240
rect 159542 79228 159548 79280
rect 159600 79268 159606 79280
rect 170306 79268 170312 79280
rect 159600 79240 170312 79268
rect 159600 79228 159606 79240
rect 170306 79228 170312 79240
rect 170364 79228 170370 79280
rect 171410 79228 171416 79280
rect 171468 79268 171474 79280
rect 171870 79268 171876 79280
rect 171468 79240 171876 79268
rect 171468 79228 171474 79240
rect 171870 79228 171876 79240
rect 171928 79228 171934 79280
rect 173158 79228 173164 79280
rect 173216 79268 173222 79280
rect 199102 79268 199108 79280
rect 173216 79240 199108 79268
rect 173216 79228 173222 79240
rect 199102 79228 199108 79240
rect 199160 79268 199166 79280
rect 200086 79268 200114 79308
rect 525794 79296 525800 79308
rect 525852 79296 525858 79348
rect 199160 79240 200114 79268
rect 199160 79228 199166 79240
rect 170766 79200 170772 79212
rect 154684 79172 170772 79200
rect 170766 79160 170772 79172
rect 170824 79160 170830 79212
rect 171594 79160 171600 79212
rect 171652 79200 171658 79212
rect 172238 79200 172244 79212
rect 171652 79172 172244 79200
rect 171652 79160 171658 79172
rect 172238 79160 172244 79172
rect 172296 79160 172302 79212
rect 172330 79160 172336 79212
rect 172388 79200 172394 79212
rect 198090 79200 198096 79212
rect 172388 79172 198096 79200
rect 172388 79160 172394 79172
rect 198090 79160 198096 79172
rect 198148 79160 198154 79212
rect 118786 79092 118792 79144
rect 118844 79132 118850 79144
rect 145006 79132 145012 79144
rect 118844 79104 145012 79132
rect 118844 79092 118850 79104
rect 145006 79092 145012 79104
rect 145064 79092 145070 79144
rect 146662 79092 146668 79144
rect 146720 79132 146726 79144
rect 146720 79104 150940 79132
rect 146720 79092 146726 79104
rect 118970 79024 118976 79076
rect 119028 79064 119034 79076
rect 146294 79064 146300 79076
rect 119028 79036 146300 79064
rect 119028 79024 119034 79036
rect 146294 79024 146300 79036
rect 146352 79024 146358 79076
rect 147030 79024 147036 79076
rect 147088 79064 147094 79076
rect 147214 79064 147220 79076
rect 147088 79036 147220 79064
rect 147088 79024 147094 79036
rect 147214 79024 147220 79036
rect 147272 79024 147278 79076
rect 150912 79064 150940 79104
rect 150986 79092 150992 79144
rect 151044 79132 151050 79144
rect 159542 79132 159548 79144
rect 151044 79104 159548 79132
rect 151044 79092 151050 79104
rect 159542 79092 159548 79104
rect 159600 79092 159606 79144
rect 162210 79092 162216 79144
rect 162268 79132 162274 79144
rect 162578 79132 162584 79144
rect 162268 79104 162584 79132
rect 162268 79092 162274 79104
rect 162578 79092 162584 79104
rect 162636 79092 162642 79144
rect 164878 79092 164884 79144
rect 164936 79132 164942 79144
rect 165614 79132 165620 79144
rect 164936 79104 165620 79132
rect 164936 79092 164942 79104
rect 165614 79092 165620 79104
rect 165672 79132 165678 79144
rect 191190 79132 191196 79144
rect 165672 79104 173756 79132
rect 165672 79092 165678 79104
rect 158438 79064 158444 79076
rect 150912 79036 158444 79064
rect 158438 79024 158444 79036
rect 158496 79024 158502 79076
rect 159082 79024 159088 79076
rect 159140 79064 159146 79076
rect 159818 79064 159824 79076
rect 159140 79036 159824 79064
rect 159140 79024 159146 79036
rect 159818 79024 159824 79036
rect 159876 79024 159882 79076
rect 164970 79024 164976 79076
rect 165028 79064 165034 79076
rect 173618 79064 173624 79076
rect 165028 79036 173624 79064
rect 165028 79024 165034 79036
rect 173618 79024 173624 79036
rect 173676 79024 173682 79076
rect 173728 79064 173756 79104
rect 173912 79104 191196 79132
rect 173912 79064 173940 79104
rect 191190 79092 191196 79104
rect 191248 79092 191254 79144
rect 173728 79036 173940 79064
rect 174262 79024 174268 79076
rect 174320 79064 174326 79076
rect 203702 79064 203708 79076
rect 174320 79036 203708 79064
rect 174320 79024 174326 79036
rect 203702 79024 203708 79036
rect 203760 79024 203766 79076
rect 120626 78956 120632 79008
rect 120684 78996 120690 79008
rect 141694 78996 141700 79008
rect 120684 78968 141700 78996
rect 120684 78956 120690 78968
rect 141694 78956 141700 78968
rect 141752 78956 141758 79008
rect 146220 78968 148640 78996
rect 119338 78888 119344 78940
rect 119396 78928 119402 78940
rect 146220 78928 146248 78968
rect 119396 78900 146248 78928
rect 119396 78888 119402 78900
rect 146294 78888 146300 78940
rect 146352 78928 146358 78940
rect 147030 78928 147036 78940
rect 146352 78900 147036 78928
rect 146352 78888 146358 78900
rect 147030 78888 147036 78900
rect 147088 78888 147094 78940
rect 148612 78928 148640 78968
rect 148686 78956 148692 79008
rect 148744 78996 148750 79008
rect 161750 78996 161756 79008
rect 148744 78968 161756 78996
rect 148744 78956 148750 78968
rect 161750 78956 161756 78968
rect 161808 78996 161814 79008
rect 167454 78996 167460 79008
rect 161808 78968 167460 78996
rect 161808 78956 161814 78968
rect 167454 78956 167460 78968
rect 167512 78956 167518 79008
rect 172514 78956 172520 79008
rect 172572 78996 172578 79008
rect 174078 78996 174084 79008
rect 172572 78968 174084 78996
rect 172572 78956 172578 78968
rect 174078 78956 174084 78968
rect 174136 78956 174142 79008
rect 174722 78956 174728 79008
rect 174780 78996 174786 79008
rect 175090 78996 175096 79008
rect 174780 78968 175096 78996
rect 174780 78956 174786 78968
rect 175090 78956 175096 78968
rect 175148 78956 175154 79008
rect 175366 78956 175372 79008
rect 175424 78996 175430 79008
rect 206370 78996 206376 79008
rect 175424 78968 206376 78996
rect 175424 78956 175430 78968
rect 206370 78956 206376 78968
rect 206428 78956 206434 79008
rect 149054 78928 149060 78940
rect 148612 78900 149060 78928
rect 149054 78888 149060 78900
rect 149112 78928 149118 78940
rect 149974 78928 149980 78940
rect 149112 78900 149980 78928
rect 149112 78888 149118 78900
rect 149974 78888 149980 78900
rect 150032 78888 150038 78940
rect 164234 78888 164240 78940
rect 164292 78928 164298 78940
rect 165614 78928 165620 78940
rect 164292 78900 165620 78928
rect 164292 78888 164298 78900
rect 165614 78888 165620 78900
rect 165672 78888 165678 78940
rect 171226 78888 171232 78940
rect 171284 78928 171290 78940
rect 195422 78928 195428 78940
rect 171284 78900 195428 78928
rect 171284 78888 171290 78900
rect 195422 78888 195428 78900
rect 195480 78888 195486 78940
rect 196250 78888 196256 78940
rect 196308 78928 196314 78940
rect 196618 78928 196624 78940
rect 196308 78900 196624 78928
rect 196308 78888 196314 78900
rect 196618 78888 196624 78900
rect 196676 78928 196682 78940
rect 483014 78928 483020 78940
rect 196676 78900 483020 78928
rect 196676 78888 196682 78900
rect 483014 78888 483020 78900
rect 483072 78888 483078 78940
rect 117866 78820 117872 78872
rect 117924 78860 117930 78872
rect 149238 78860 149244 78872
rect 117924 78832 149244 78860
rect 117924 78820 117930 78832
rect 149238 78820 149244 78832
rect 149296 78820 149302 78872
rect 159634 78820 159640 78872
rect 159692 78860 159698 78872
rect 191374 78860 191380 78872
rect 159692 78832 191380 78860
rect 159692 78820 159698 78832
rect 191374 78820 191380 78832
rect 191432 78820 191438 78872
rect 198734 78820 198740 78872
rect 198792 78860 198798 78872
rect 199378 78860 199384 78872
rect 198792 78832 199384 78860
rect 198792 78820 198798 78832
rect 199378 78820 199384 78832
rect 199436 78860 199442 78872
rect 500954 78860 500960 78872
rect 199436 78832 500960 78860
rect 199436 78820 199442 78832
rect 500954 78820 500960 78832
rect 501012 78820 501018 78872
rect 132402 78752 132408 78804
rect 132460 78792 132466 78804
rect 137738 78792 137744 78804
rect 132460 78764 137744 78792
rect 132460 78752 132466 78764
rect 137738 78752 137744 78764
rect 137796 78752 137802 78804
rect 139670 78752 139676 78804
rect 139728 78792 139734 78804
rect 139854 78792 139860 78804
rect 139728 78764 139860 78792
rect 139728 78752 139734 78764
rect 139854 78752 139860 78764
rect 139912 78752 139918 78804
rect 141694 78752 141700 78804
rect 141752 78792 141758 78804
rect 147766 78792 147772 78804
rect 141752 78764 147772 78792
rect 141752 78752 141758 78764
rect 147766 78752 147772 78764
rect 147824 78752 147830 78804
rect 171962 78752 171968 78804
rect 172020 78792 172026 78804
rect 196710 78792 196716 78804
rect 172020 78764 196716 78792
rect 172020 78752 172026 78764
rect 196710 78752 196716 78764
rect 196768 78752 196774 78804
rect 196802 78752 196808 78804
rect 196860 78792 196866 78804
rect 523126 78792 523132 78804
rect 196860 78764 523132 78792
rect 196860 78752 196866 78764
rect 523126 78752 523132 78764
rect 523184 78752 523190 78804
rect 127434 78684 127440 78736
rect 127492 78724 127498 78736
rect 132494 78724 132500 78736
rect 127492 78696 132500 78724
rect 127492 78684 127498 78696
rect 132494 78684 132500 78696
rect 132552 78684 132558 78736
rect 133598 78684 133604 78736
rect 133656 78724 133662 78736
rect 133874 78724 133880 78736
rect 133656 78696 133880 78724
rect 133656 78684 133662 78696
rect 133874 78684 133880 78696
rect 133932 78684 133938 78736
rect 134518 78684 134524 78736
rect 134576 78724 134582 78736
rect 138474 78724 138480 78736
rect 134576 78696 138480 78724
rect 134576 78684 134582 78696
rect 138474 78684 138480 78696
rect 138532 78684 138538 78736
rect 144362 78684 144368 78736
rect 144420 78724 144426 78736
rect 150618 78724 150624 78736
rect 144420 78696 150624 78724
rect 144420 78684 144426 78696
rect 150618 78684 150624 78696
rect 150676 78724 150682 78736
rect 151170 78724 151176 78736
rect 150676 78696 151176 78724
rect 150676 78684 150682 78696
rect 151170 78684 151176 78696
rect 151228 78684 151234 78736
rect 162026 78684 162032 78736
rect 162084 78724 162090 78736
rect 162084 78696 172468 78724
rect 162084 78684 162090 78696
rect 102134 78616 102140 78668
rect 102192 78656 102198 78668
rect 102870 78656 102876 78668
rect 102192 78628 102876 78656
rect 102192 78616 102198 78628
rect 102870 78616 102876 78628
rect 102928 78656 102934 78668
rect 133966 78656 133972 78668
rect 102928 78628 133972 78656
rect 102928 78616 102934 78628
rect 133966 78616 133972 78628
rect 134024 78616 134030 78668
rect 138750 78616 138756 78668
rect 138808 78656 138814 78668
rect 139026 78656 139032 78668
rect 138808 78628 139032 78656
rect 138808 78616 138814 78628
rect 139026 78616 139032 78628
rect 139084 78616 139090 78668
rect 151262 78616 151268 78668
rect 151320 78656 151326 78668
rect 151630 78656 151636 78668
rect 151320 78628 151636 78656
rect 151320 78616 151326 78628
rect 151630 78616 151636 78628
rect 151688 78616 151694 78668
rect 151998 78616 152004 78668
rect 152056 78656 152062 78668
rect 153102 78656 153108 78668
rect 152056 78628 153108 78656
rect 152056 78616 152062 78628
rect 153102 78616 153108 78628
rect 153160 78616 153166 78668
rect 153930 78616 153936 78668
rect 153988 78656 153994 78668
rect 154482 78656 154488 78668
rect 153988 78628 154488 78656
rect 153988 78616 153994 78628
rect 154482 78616 154488 78628
rect 154540 78616 154546 78668
rect 163130 78616 163136 78668
rect 163188 78656 163194 78668
rect 163774 78656 163780 78668
rect 163188 78628 163780 78656
rect 163188 78616 163194 78628
rect 163774 78616 163780 78628
rect 163832 78616 163838 78668
rect 164326 78616 164332 78668
rect 164384 78656 164390 78668
rect 164510 78656 164516 78668
rect 164384 78628 164516 78656
rect 164384 78616 164390 78628
rect 164510 78616 164516 78628
rect 164568 78616 164574 78668
rect 172440 78656 172468 78696
rect 173342 78684 173348 78736
rect 173400 78724 173406 78736
rect 196526 78724 196532 78736
rect 173400 78696 196532 78724
rect 173400 78684 173406 78696
rect 196526 78684 196532 78696
rect 196584 78684 196590 78736
rect 199102 78684 199108 78736
rect 199160 78724 199166 78736
rect 199562 78724 199568 78736
rect 199160 78696 199568 78724
rect 199160 78684 199166 78696
rect 199562 78684 199568 78696
rect 199620 78724 199626 78736
rect 536834 78724 536840 78736
rect 199620 78696 536840 78724
rect 199620 78684 199626 78696
rect 536834 78684 536840 78696
rect 536892 78684 536898 78736
rect 172440 78628 176700 78656
rect 104250 78548 104256 78600
rect 104308 78588 104314 78600
rect 132586 78588 132592 78600
rect 104308 78560 132592 78588
rect 104308 78548 104314 78560
rect 132586 78548 132592 78560
rect 132644 78548 132650 78600
rect 132678 78548 132684 78600
rect 132736 78588 132742 78600
rect 142338 78588 142344 78600
rect 132736 78560 142344 78588
rect 132736 78548 132742 78560
rect 142338 78548 142344 78560
rect 142396 78548 142402 78600
rect 170766 78548 170772 78600
rect 170824 78588 170830 78600
rect 176286 78588 176292 78600
rect 170824 78560 176292 78588
rect 170824 78548 170830 78560
rect 176286 78548 176292 78560
rect 176344 78548 176350 78600
rect 176672 78588 176700 78628
rect 176746 78616 176752 78668
rect 176804 78656 176810 78668
rect 177206 78656 177212 78668
rect 176804 78628 177212 78656
rect 176804 78616 176810 78628
rect 177206 78616 177212 78628
rect 177264 78616 177270 78668
rect 177666 78588 177672 78600
rect 176672 78560 177672 78588
rect 177666 78548 177672 78560
rect 177724 78548 177730 78600
rect 178770 78548 178776 78600
rect 178828 78588 178834 78600
rect 178828 78560 200114 78588
rect 178828 78548 178834 78560
rect 123018 78480 123024 78532
rect 123076 78520 123082 78532
rect 131298 78520 131304 78532
rect 123076 78492 131304 78520
rect 123076 78480 123082 78492
rect 131298 78480 131304 78492
rect 131356 78520 131362 78532
rect 132402 78520 132408 78532
rect 131356 78492 132408 78520
rect 131356 78480 131362 78492
rect 132402 78480 132408 78492
rect 132460 78480 132466 78532
rect 132494 78480 132500 78532
rect 132552 78520 132558 78532
rect 132552 78492 136312 78520
rect 132552 78480 132558 78492
rect 107286 78452 107292 78464
rect 103486 78424 107292 78452
rect 46934 78344 46940 78396
rect 46992 78384 46998 78396
rect 103486 78384 103514 78424
rect 107286 78412 107292 78424
rect 107344 78452 107350 78464
rect 136174 78452 136180 78464
rect 107344 78424 136180 78452
rect 107344 78412 107350 78424
rect 136174 78412 136180 78424
rect 136232 78412 136238 78464
rect 136284 78452 136312 78492
rect 139762 78480 139768 78532
rect 139820 78520 139826 78532
rect 140130 78520 140136 78532
rect 139820 78492 140136 78520
rect 139820 78480 139826 78492
rect 140130 78480 140136 78492
rect 140188 78480 140194 78532
rect 170214 78480 170220 78532
rect 170272 78520 170278 78532
rect 196250 78520 196256 78532
rect 170272 78492 196256 78520
rect 170272 78480 170278 78492
rect 196250 78480 196256 78492
rect 196308 78480 196314 78532
rect 141878 78452 141884 78464
rect 136284 78424 141884 78452
rect 141878 78412 141884 78424
rect 141936 78412 141942 78464
rect 159542 78412 159548 78464
rect 159600 78452 159606 78464
rect 161934 78452 161940 78464
rect 159600 78424 161940 78452
rect 159600 78412 159606 78424
rect 161934 78412 161940 78424
rect 161992 78452 161998 78464
rect 162394 78452 162400 78464
rect 161992 78424 162400 78452
rect 161992 78412 161998 78424
rect 162394 78412 162400 78424
rect 162452 78412 162458 78464
rect 167178 78412 167184 78464
rect 167236 78452 167242 78464
rect 182910 78452 182916 78464
rect 167236 78424 182916 78452
rect 167236 78412 167242 78424
rect 182910 78412 182916 78424
rect 182968 78412 182974 78464
rect 46992 78356 103514 78384
rect 46992 78344 46998 78356
rect 122098 78344 122104 78396
rect 122156 78384 122162 78396
rect 149146 78384 149152 78396
rect 122156 78356 149152 78384
rect 122156 78344 122162 78356
rect 149146 78344 149152 78356
rect 149204 78344 149210 78396
rect 173250 78344 173256 78396
rect 173308 78384 173314 78396
rect 173802 78384 173808 78396
rect 173308 78356 173808 78384
rect 173308 78344 173314 78356
rect 173802 78344 173808 78356
rect 173860 78344 173866 78396
rect 173894 78344 173900 78396
rect 173952 78384 173958 78396
rect 174538 78384 174544 78396
rect 173952 78356 174544 78384
rect 173952 78344 173958 78356
rect 174538 78344 174544 78356
rect 174596 78344 174602 78396
rect 174722 78344 174728 78396
rect 174780 78384 174786 78396
rect 175274 78384 175280 78396
rect 174780 78356 175280 78384
rect 174780 78344 174786 78356
rect 175274 78344 175280 78356
rect 175332 78344 175338 78396
rect 175642 78344 175648 78396
rect 175700 78384 175706 78396
rect 176102 78384 176108 78396
rect 175700 78356 176108 78384
rect 175700 78344 175706 78356
rect 176102 78344 176108 78356
rect 176160 78344 176166 78396
rect 178494 78344 178500 78396
rect 178552 78384 178558 78396
rect 200086 78384 200114 78560
rect 203334 78384 203340 78396
rect 178552 78356 186314 78384
rect 200086 78356 203340 78384
rect 178552 78344 178558 78356
rect 57974 78276 57980 78328
rect 58032 78316 58038 78328
rect 107286 78316 107292 78328
rect 58032 78288 107292 78316
rect 58032 78276 58038 78288
rect 107286 78276 107292 78288
rect 107344 78276 107350 78328
rect 122006 78276 122012 78328
rect 122064 78316 122070 78328
rect 148318 78316 148324 78328
rect 122064 78288 148324 78316
rect 122064 78276 122070 78288
rect 148318 78276 148324 78288
rect 148376 78276 148382 78328
rect 169018 78276 169024 78328
rect 169076 78316 169082 78328
rect 186286 78316 186314 78356
rect 203334 78344 203340 78356
rect 203392 78384 203398 78396
rect 287698 78384 287704 78396
rect 203392 78356 287704 78384
rect 203392 78344 203398 78356
rect 287698 78344 287704 78356
rect 287756 78344 287762 78396
rect 255958 78316 255964 78328
rect 169076 78288 179552 78316
rect 186286 78288 255964 78316
rect 169076 78276 169082 78288
rect 106918 78248 106924 78260
rect 103486 78220 106924 78248
rect 20714 78140 20720 78192
rect 20772 78180 20778 78192
rect 102134 78180 102140 78192
rect 20772 78152 102140 78180
rect 20772 78140 20778 78152
rect 102134 78140 102140 78152
rect 102192 78140 102198 78192
rect 6914 78072 6920 78124
rect 6972 78112 6978 78124
rect 103486 78112 103514 78220
rect 106918 78208 106924 78220
rect 106976 78248 106982 78260
rect 126974 78248 126980 78260
rect 106976 78220 126980 78248
rect 106976 78208 106982 78220
rect 126974 78208 126980 78220
rect 127032 78208 127038 78260
rect 132310 78248 132316 78260
rect 127084 78220 132316 78248
rect 127084 78180 127112 78220
rect 132310 78208 132316 78220
rect 132368 78208 132374 78260
rect 146570 78208 146576 78260
rect 146628 78248 146634 78260
rect 179414 78248 179420 78260
rect 146628 78220 179420 78248
rect 146628 78208 146634 78220
rect 179414 78208 179420 78220
rect 179472 78208 179478 78260
rect 6972 78084 103514 78112
rect 113146 78152 127112 78180
rect 6972 78072 6978 78084
rect 2866 78004 2872 78056
rect 2924 78044 2930 78056
rect 104250 78044 104256 78056
rect 2924 78016 104256 78044
rect 2924 78004 2930 78016
rect 104250 78004 104256 78016
rect 104308 78004 104314 78056
rect 2774 77936 2780 77988
rect 2832 77976 2838 77988
rect 108390 77976 108396 77988
rect 2832 77948 108396 77976
rect 2832 77936 2838 77948
rect 108390 77936 108396 77948
rect 108448 77976 108454 77988
rect 113146 77976 113174 78152
rect 127158 78140 127164 78192
rect 127216 78180 127222 78192
rect 141050 78180 141056 78192
rect 127216 78152 141056 78180
rect 127216 78140 127222 78152
rect 141050 78140 141056 78152
rect 141108 78140 141114 78192
rect 141694 78140 141700 78192
rect 141752 78180 141758 78192
rect 142890 78180 142896 78192
rect 141752 78152 142896 78180
rect 141752 78140 141758 78152
rect 142890 78140 142896 78152
rect 142948 78140 142954 78192
rect 171870 78140 171876 78192
rect 171928 78180 171934 78192
rect 172330 78180 172336 78192
rect 171928 78152 172336 78180
rect 171928 78140 171934 78152
rect 172330 78140 172336 78152
rect 172388 78140 172394 78192
rect 175274 78140 175280 78192
rect 175332 78180 175338 78192
rect 176194 78180 176200 78192
rect 175332 78152 176200 78180
rect 175332 78140 175338 78152
rect 176194 78140 176200 78152
rect 176252 78140 176258 78192
rect 179524 78180 179552 78288
rect 255958 78276 255964 78288
rect 256016 78276 256022 78328
rect 192570 78208 192576 78260
rect 192628 78248 192634 78260
rect 324314 78248 324320 78260
rect 192628 78220 324320 78248
rect 192628 78208 192634 78220
rect 324314 78208 324320 78220
rect 324372 78208 324378 78260
rect 337378 78180 337384 78192
rect 179524 78152 337384 78180
rect 337378 78140 337384 78152
rect 337436 78140 337442 78192
rect 123202 78072 123208 78124
rect 123260 78112 123266 78124
rect 146110 78112 146116 78124
rect 123260 78084 146116 78112
rect 123260 78072 123266 78084
rect 146110 78072 146116 78084
rect 146168 78072 146174 78124
rect 162946 78072 162952 78124
rect 163004 78112 163010 78124
rect 393314 78112 393320 78124
rect 163004 78084 393320 78112
rect 163004 78072 163010 78084
rect 393314 78072 393320 78084
rect 393372 78072 393378 78124
rect 113634 78004 113640 78056
rect 113692 78044 113698 78056
rect 130654 78044 130660 78056
rect 113692 78016 130660 78044
rect 113692 78004 113698 78016
rect 130654 78004 130660 78016
rect 130712 78004 130718 78056
rect 137278 78044 137284 78056
rect 130948 78016 137284 78044
rect 108448 77948 113174 77976
rect 108448 77936 108454 77948
rect 113726 77936 113732 77988
rect 113784 77976 113790 77988
rect 123018 77976 123024 77988
rect 113784 77948 123024 77976
rect 113784 77936 113790 77948
rect 123018 77936 123024 77948
rect 123076 77936 123082 77988
rect 129826 77976 129832 77988
rect 123312 77948 129832 77976
rect 115106 77800 115112 77852
rect 115164 77840 115170 77852
rect 123312 77840 123340 77948
rect 129826 77936 129832 77948
rect 129884 77976 129890 77988
rect 130948 77976 130976 78016
rect 137278 78004 137284 78016
rect 137336 78004 137342 78056
rect 139118 78004 139124 78056
rect 139176 78044 139182 78056
rect 139394 78044 139400 78056
rect 139176 78016 139400 78044
rect 139176 78004 139182 78016
rect 139394 78004 139400 78016
rect 139452 78004 139458 78056
rect 164786 78004 164792 78056
rect 164844 78044 164850 78056
rect 165522 78044 165528 78056
rect 164844 78016 165528 78044
rect 164844 78004 164850 78016
rect 165522 78004 165528 78016
rect 165580 78004 165586 78056
rect 169570 78004 169576 78056
rect 169628 78044 169634 78056
rect 400858 78044 400864 78056
rect 169628 78016 400864 78044
rect 169628 78004 169634 78016
rect 400858 78004 400864 78016
rect 400916 78004 400922 78056
rect 129884 77948 130976 77976
rect 129884 77936 129890 77948
rect 131574 77936 131580 77988
rect 131632 77976 131638 77988
rect 142430 77976 142436 77988
rect 131632 77948 142436 77976
rect 131632 77936 131638 77948
rect 142430 77936 142436 77948
rect 142488 77936 142494 77988
rect 163406 77936 163412 77988
rect 163464 77976 163470 77988
rect 400214 77976 400220 77988
rect 163464 77948 400220 77976
rect 163464 77936 163470 77948
rect 400214 77936 400220 77948
rect 400272 77936 400278 77988
rect 123386 77868 123392 77920
rect 123444 77908 123450 77920
rect 142614 77908 142620 77920
rect 123444 77880 142620 77908
rect 123444 77868 123450 77880
rect 142614 77868 142620 77880
rect 142672 77908 142678 77920
rect 142982 77908 142988 77920
rect 142672 77880 142988 77908
rect 142672 77868 142678 77880
rect 142982 77868 142988 77880
rect 143040 77868 143046 77920
rect 166626 77868 166632 77920
rect 166684 77908 166690 77920
rect 181622 77908 181628 77920
rect 166684 77880 181628 77908
rect 166684 77868 166690 77880
rect 181622 77868 181628 77880
rect 181680 77868 181686 77920
rect 115164 77812 123340 77840
rect 115164 77800 115170 77812
rect 130654 77800 130660 77852
rect 130712 77840 130718 77852
rect 132862 77840 132868 77852
rect 130712 77812 132868 77840
rect 130712 77800 130718 77812
rect 132862 77800 132868 77812
rect 132920 77800 132926 77852
rect 134150 77800 134156 77852
rect 134208 77840 134214 77852
rect 134426 77840 134432 77852
rect 134208 77812 134432 77840
rect 134208 77800 134214 77812
rect 134426 77800 134432 77812
rect 134484 77800 134490 77852
rect 135990 77800 135996 77852
rect 136048 77840 136054 77852
rect 136450 77840 136456 77852
rect 136048 77812 136456 77840
rect 136048 77800 136054 77812
rect 136450 77800 136456 77812
rect 136508 77800 136514 77852
rect 136818 77800 136824 77852
rect 136876 77840 136882 77852
rect 137186 77840 137192 77852
rect 136876 77812 137192 77840
rect 136876 77800 136882 77812
rect 137186 77800 137192 77812
rect 137244 77800 137250 77852
rect 142430 77800 142436 77852
rect 142488 77840 142494 77852
rect 143442 77840 143448 77852
rect 142488 77812 143448 77840
rect 142488 77800 142494 77812
rect 143442 77800 143448 77812
rect 143500 77800 143506 77852
rect 165798 77800 165804 77852
rect 165856 77840 165862 77852
rect 180702 77840 180708 77852
rect 165856 77812 180708 77840
rect 165856 77800 165862 77812
rect 180702 77800 180708 77812
rect 180760 77800 180766 77852
rect 107286 77732 107292 77784
rect 107344 77772 107350 77784
rect 136082 77772 136088 77784
rect 107344 77744 136088 77772
rect 107344 77732 107350 77744
rect 136082 77732 136088 77744
rect 136140 77732 136146 77784
rect 137830 77732 137836 77784
rect 137888 77772 137894 77784
rect 143718 77772 143724 77784
rect 137888 77744 143724 77772
rect 137888 77732 137894 77744
rect 143718 77732 143724 77744
rect 143776 77772 143782 77784
rect 144362 77772 144368 77784
rect 143776 77744 144368 77772
rect 143776 77732 143782 77744
rect 144362 77732 144368 77744
rect 144420 77732 144426 77784
rect 153470 77732 153476 77784
rect 153528 77772 153534 77784
rect 154390 77772 154396 77784
rect 153528 77744 154396 77772
rect 153528 77732 153534 77744
rect 154390 77732 154396 77744
rect 154448 77732 154454 77784
rect 164602 77732 164608 77784
rect 164660 77772 164666 77784
rect 178770 77772 178776 77784
rect 164660 77744 178776 77772
rect 164660 77732 164666 77744
rect 178770 77732 178776 77744
rect 178828 77732 178834 77784
rect 132954 77664 132960 77716
rect 133012 77704 133018 77716
rect 141694 77704 141700 77716
rect 133012 77676 141700 77704
rect 133012 77664 133018 77676
rect 141694 77664 141700 77676
rect 141752 77664 141758 77716
rect 157610 77664 157616 77716
rect 157668 77704 157674 77716
rect 192570 77704 192576 77716
rect 157668 77676 192576 77704
rect 157668 77664 157674 77676
rect 192570 77664 192576 77676
rect 192628 77664 192634 77716
rect 131022 77596 131028 77648
rect 131080 77636 131086 77648
rect 144914 77636 144920 77648
rect 131080 77608 144920 77636
rect 131080 77596 131086 77608
rect 144914 77596 144920 77608
rect 144972 77596 144978 77648
rect 148318 77596 148324 77648
rect 148376 77636 148382 77648
rect 148502 77636 148508 77648
rect 148376 77608 148508 77636
rect 148376 77596 148382 77608
rect 148502 77596 148508 77608
rect 148560 77596 148566 77648
rect 164602 77596 164608 77648
rect 164660 77636 164666 77648
rect 164878 77636 164884 77648
rect 164660 77608 164884 77636
rect 164660 77596 164666 77608
rect 164878 77596 164884 77608
rect 164936 77596 164942 77648
rect 165154 77596 165160 77648
rect 165212 77636 165218 77648
rect 180150 77636 180156 77648
rect 165212 77608 180156 77636
rect 165212 77596 165218 77608
rect 180150 77596 180156 77608
rect 180208 77596 180214 77648
rect 176010 77528 176016 77580
rect 176068 77568 176074 77580
rect 176378 77568 176384 77580
rect 176068 77540 176384 77568
rect 176068 77528 176074 77540
rect 176378 77528 176384 77540
rect 176436 77528 176442 77580
rect 176838 77528 176844 77580
rect 176896 77568 176902 77580
rect 177114 77568 177120 77580
rect 176896 77540 177120 77568
rect 176896 77528 176902 77540
rect 177114 77528 177120 77540
rect 177172 77528 177178 77580
rect 140958 77460 140964 77512
rect 141016 77500 141022 77512
rect 141326 77500 141332 77512
rect 141016 77472 141332 77500
rect 141016 77460 141022 77472
rect 141326 77460 141332 77472
rect 141384 77460 141390 77512
rect 146110 77460 146116 77512
rect 146168 77500 146174 77512
rect 148318 77500 148324 77512
rect 146168 77472 148324 77500
rect 146168 77460 146174 77472
rect 148318 77460 148324 77472
rect 148376 77460 148382 77512
rect 162946 77460 162952 77512
rect 163004 77500 163010 77512
rect 163314 77500 163320 77512
rect 163004 77472 163320 77500
rect 163004 77460 163010 77472
rect 163314 77460 163320 77472
rect 163372 77460 163378 77512
rect 170306 77460 170312 77512
rect 170364 77500 170370 77512
rect 178862 77500 178868 77512
rect 170364 77472 178868 77500
rect 170364 77460 170370 77472
rect 178862 77460 178868 77472
rect 178920 77460 178926 77512
rect 173618 77392 173624 77444
rect 173676 77432 173682 77444
rect 178034 77432 178040 77444
rect 173676 77404 178040 77432
rect 173676 77392 173682 77404
rect 178034 77392 178040 77404
rect 178092 77392 178098 77444
rect 160646 77324 160652 77376
rect 160704 77364 160710 77376
rect 163314 77364 163320 77376
rect 160704 77336 163320 77364
rect 160704 77324 160710 77336
rect 163314 77324 163320 77336
rect 163372 77324 163378 77376
rect 151538 77256 151544 77308
rect 151596 77296 151602 77308
rect 151596 77268 151676 77296
rect 151596 77256 151602 77268
rect 112622 77188 112628 77240
rect 112680 77228 112686 77240
rect 146294 77228 146300 77240
rect 112680 77200 146300 77228
rect 112680 77188 112686 77200
rect 146294 77188 146300 77200
rect 146352 77188 146358 77240
rect 151446 77188 151452 77240
rect 151504 77228 151510 77240
rect 151648 77228 151676 77268
rect 163222 77256 163228 77308
rect 163280 77296 163286 77308
rect 166258 77296 166264 77308
rect 163280 77268 166264 77296
rect 163280 77256 163286 77268
rect 166258 77256 166264 77268
rect 166316 77256 166322 77308
rect 171318 77256 171324 77308
rect 171376 77296 171382 77308
rect 171686 77296 171692 77308
rect 171376 77268 171692 77296
rect 171376 77256 171382 77268
rect 171686 77256 171692 77268
rect 171744 77256 171750 77308
rect 172514 77256 172520 77308
rect 172572 77296 172578 77308
rect 173342 77296 173348 77308
rect 172572 77268 173348 77296
rect 172572 77256 172578 77268
rect 173342 77256 173348 77268
rect 173400 77256 173406 77308
rect 151504 77200 151676 77228
rect 151504 77188 151510 77200
rect 161566 77188 161572 77240
rect 161624 77228 161630 77240
rect 196710 77228 196716 77240
rect 161624 77200 196716 77228
rect 161624 77188 161630 77200
rect 196710 77188 196716 77200
rect 196768 77188 196774 77240
rect 102778 77160 102784 77172
rect 84166 77132 102784 77160
rect 72418 76780 72424 76832
rect 72476 76820 72482 76832
rect 84166 76820 84194 77132
rect 102778 77120 102784 77132
rect 102836 77160 102842 77172
rect 137462 77160 137468 77172
rect 102836 77132 137468 77160
rect 102836 77120 102842 77132
rect 137462 77120 137468 77132
rect 137520 77120 137526 77172
rect 163038 77120 163044 77172
rect 163096 77160 163102 77172
rect 197814 77160 197820 77172
rect 163096 77132 197820 77160
rect 163096 77120 163102 77132
rect 197814 77120 197820 77132
rect 197872 77160 197878 77172
rect 198182 77160 198188 77172
rect 197872 77132 198188 77160
rect 197872 77120 197878 77132
rect 198182 77120 198188 77132
rect 198240 77120 198246 77172
rect 114554 77052 114560 77104
rect 114612 77092 114618 77104
rect 115198 77092 115204 77104
rect 114612 77064 115204 77092
rect 114612 77052 114618 77064
rect 115198 77052 115204 77064
rect 115256 77052 115262 77104
rect 115658 77052 115664 77104
rect 115716 77092 115722 77104
rect 115716 77064 138014 77092
rect 115716 77052 115722 77064
rect 100754 76984 100760 77036
rect 100812 77024 100818 77036
rect 101582 77024 101588 77036
rect 100812 76996 101588 77024
rect 100812 76984 100818 76996
rect 101582 76984 101588 76996
rect 101640 77024 101646 77036
rect 134978 77024 134984 77036
rect 101640 76996 134984 77024
rect 101640 76984 101646 76996
rect 134978 76984 134984 76996
rect 135036 76984 135042 77036
rect 135346 76984 135352 77036
rect 135404 77024 135410 77036
rect 135622 77024 135628 77036
rect 135404 76996 135628 77024
rect 135404 76984 135410 76996
rect 135622 76984 135628 76996
rect 135680 76984 135686 77036
rect 137986 77024 138014 77064
rect 159726 77052 159732 77104
rect 159784 77092 159790 77104
rect 193582 77092 193588 77104
rect 159784 77064 193588 77092
rect 159784 77052 159790 77064
rect 193582 77052 193588 77064
rect 193640 77052 193646 77104
rect 148410 77024 148416 77036
rect 137986 76996 148416 77024
rect 148410 76984 148416 76996
rect 148468 76984 148474 77036
rect 155494 76984 155500 77036
rect 155552 77024 155558 77036
rect 155552 76996 161244 77024
rect 155552 76984 155558 76996
rect 117038 76916 117044 76968
rect 117096 76956 117102 76968
rect 148870 76956 148876 76968
rect 117096 76928 148876 76956
rect 117096 76916 117102 76928
rect 148870 76916 148876 76928
rect 148928 76916 148934 76968
rect 155954 76916 155960 76968
rect 156012 76956 156018 76968
rect 156874 76956 156880 76968
rect 156012 76928 156880 76956
rect 156012 76916 156018 76928
rect 156874 76916 156880 76928
rect 156932 76916 156938 76968
rect 161216 76956 161244 76996
rect 162118 76984 162124 77036
rect 162176 77024 162182 77036
rect 162762 77024 162768 77036
rect 162176 76996 162768 77024
rect 162176 76984 162182 76996
rect 162762 76984 162768 76996
rect 162820 77024 162826 77036
rect 191098 77024 191104 77036
rect 162820 76996 191104 77024
rect 162820 76984 162826 76996
rect 191098 76984 191104 76996
rect 191156 76984 191162 77036
rect 177758 76956 177764 76968
rect 161216 76928 177764 76956
rect 177758 76916 177764 76928
rect 177816 76916 177822 76968
rect 177942 76916 177948 76968
rect 178000 76956 178006 76968
rect 180058 76956 180064 76968
rect 178000 76928 180064 76956
rect 178000 76916 178006 76928
rect 180058 76916 180064 76928
rect 180116 76916 180122 76968
rect 188982 76916 188988 76968
rect 189040 76956 189046 76968
rect 189166 76956 189172 76968
rect 189040 76928 189172 76956
rect 189040 76916 189046 76928
rect 189166 76916 189172 76928
rect 189224 76916 189230 76968
rect 105722 76888 105728 76900
rect 72476 76792 84194 76820
rect 103486 76860 105728 76888
rect 72476 76780 72482 76792
rect 64138 76712 64144 76764
rect 64196 76752 64202 76764
rect 103486 76752 103514 76860
rect 105722 76848 105728 76860
rect 105780 76888 105786 76900
rect 136910 76888 136916 76900
rect 105780 76860 136916 76888
rect 105780 76848 105786 76860
rect 136910 76848 136916 76860
rect 136968 76848 136974 76900
rect 145282 76848 145288 76900
rect 145340 76888 145346 76900
rect 146202 76888 146208 76900
rect 145340 76860 146208 76888
rect 145340 76848 145346 76860
rect 146202 76848 146208 76860
rect 146260 76848 146266 76900
rect 151078 76848 151084 76900
rect 151136 76888 151142 76900
rect 211798 76888 211804 76900
rect 151136 76860 211804 76888
rect 151136 76848 151142 76860
rect 211798 76848 211804 76860
rect 211856 76848 211862 76900
rect 119706 76780 119712 76832
rect 119764 76820 119770 76832
rect 151446 76820 151452 76832
rect 119764 76792 151452 76820
rect 119764 76780 119770 76792
rect 151446 76780 151452 76792
rect 151504 76820 151510 76832
rect 224218 76820 224224 76832
rect 151504 76792 224224 76820
rect 151504 76780 151510 76792
rect 224218 76780 224224 76792
rect 224276 76780 224282 76832
rect 64196 76724 103514 76752
rect 64196 76712 64202 76724
rect 111334 76712 111340 76764
rect 111392 76752 111398 76764
rect 141050 76752 141056 76764
rect 111392 76724 141056 76752
rect 111392 76712 111398 76724
rect 141050 76712 141056 76724
rect 141108 76752 141114 76764
rect 141418 76752 141424 76764
rect 141108 76724 141424 76752
rect 141108 76712 141114 76724
rect 141418 76712 141424 76724
rect 141476 76712 141482 76764
rect 143166 76712 143172 76764
rect 143224 76752 143230 76764
rect 143442 76752 143448 76764
rect 143224 76724 143448 76752
rect 143224 76712 143230 76724
rect 143442 76712 143448 76724
rect 143500 76712 143506 76764
rect 149146 76712 149152 76764
rect 149204 76752 149210 76764
rect 149790 76752 149796 76764
rect 149204 76724 149796 76752
rect 149204 76712 149210 76724
rect 149790 76712 149796 76724
rect 149848 76712 149854 76764
rect 152642 76712 152648 76764
rect 152700 76752 152706 76764
rect 260834 76752 260840 76764
rect 152700 76724 260840 76752
rect 152700 76712 152706 76724
rect 260834 76712 260840 76724
rect 260892 76712 260898 76764
rect 34514 76644 34520 76696
rect 34572 76684 34578 76696
rect 100754 76684 100760 76696
rect 34572 76656 100760 76684
rect 34572 76644 34578 76656
rect 100754 76644 100760 76656
rect 100812 76644 100818 76696
rect 115198 76644 115204 76696
rect 115256 76684 115262 76696
rect 127158 76684 127164 76696
rect 115256 76656 127164 76684
rect 115256 76644 115262 76656
rect 127158 76644 127164 76656
rect 127216 76644 127222 76696
rect 153194 76644 153200 76696
rect 153252 76684 153258 76696
rect 153470 76684 153476 76696
rect 153252 76656 153476 76684
rect 153252 76644 153258 76656
rect 153470 76644 153476 76656
rect 153528 76644 153534 76696
rect 155218 76644 155224 76696
rect 155276 76684 155282 76696
rect 171778 76684 171784 76696
rect 155276 76656 171784 76684
rect 155276 76644 155282 76656
rect 171778 76644 171784 76656
rect 171836 76644 171842 76696
rect 181438 76684 181444 76696
rect 171888 76656 181444 76684
rect 52454 76576 52460 76628
rect 52512 76616 52518 76628
rect 135346 76616 135352 76628
rect 52512 76588 135352 76616
rect 52512 76576 52518 76588
rect 135346 76576 135352 76588
rect 135404 76576 135410 76628
rect 149514 76576 149520 76628
rect 149572 76616 149578 76628
rect 149974 76616 149980 76628
rect 149572 76588 149980 76616
rect 149572 76576 149578 76588
rect 149974 76576 149980 76588
rect 150032 76576 150038 76628
rect 168466 76576 168472 76628
rect 168524 76616 168530 76628
rect 169294 76616 169300 76628
rect 168524 76588 169300 76616
rect 168524 76576 168530 76588
rect 169294 76576 169300 76588
rect 169352 76576 169358 76628
rect 35894 76508 35900 76560
rect 35952 76548 35958 76560
rect 134242 76548 134248 76560
rect 35952 76520 134248 76548
rect 35952 76508 35958 76520
rect 134242 76508 134248 76520
rect 134300 76508 134306 76560
rect 147122 76508 147128 76560
rect 147180 76548 147186 76560
rect 171888 76548 171916 76656
rect 181438 76644 181444 76656
rect 181496 76644 181502 76696
rect 193582 76644 193588 76696
rect 193640 76684 193646 76696
rect 194042 76684 194048 76696
rect 193640 76656 194048 76684
rect 193640 76644 193646 76656
rect 194042 76644 194048 76656
rect 194100 76684 194106 76696
rect 353294 76684 353300 76696
rect 194100 76656 353300 76684
rect 194100 76644 194106 76656
rect 353294 76644 353300 76656
rect 353352 76644 353358 76696
rect 187694 76616 187700 76628
rect 147180 76520 171916 76548
rect 173590 76588 187700 76616
rect 147180 76508 147186 76520
rect 112530 76440 112536 76492
rect 112588 76480 112594 76492
rect 138290 76480 138296 76492
rect 112588 76452 138296 76480
rect 112588 76440 112594 76452
rect 138290 76440 138296 76452
rect 138348 76440 138354 76492
rect 170858 76440 170864 76492
rect 170916 76480 170922 76492
rect 173590 76480 173618 76588
rect 187694 76576 187700 76588
rect 187752 76576 187758 76628
rect 196710 76576 196716 76628
rect 196768 76616 196774 76628
rect 373994 76616 374000 76628
rect 196768 76588 374000 76616
rect 196768 76576 196774 76588
rect 373994 76576 374000 76588
rect 374052 76576 374058 76628
rect 174538 76508 174544 76560
rect 174596 76548 174602 76560
rect 174722 76548 174728 76560
rect 174596 76520 174728 76548
rect 174596 76508 174602 76520
rect 174722 76508 174728 76520
rect 174780 76508 174786 76560
rect 186682 76548 186688 76560
rect 179386 76520 186688 76548
rect 170916 76452 173618 76480
rect 170916 76440 170922 76452
rect 170674 76372 170680 76424
rect 170732 76412 170738 76424
rect 179386 76412 179414 76520
rect 186682 76508 186688 76520
rect 186740 76508 186746 76560
rect 197814 76508 197820 76560
rect 197872 76548 197878 76560
rect 391934 76548 391940 76560
rect 197872 76520 391940 76548
rect 197872 76508 197878 76520
rect 391934 76508 391940 76520
rect 391992 76508 391998 76560
rect 170732 76384 179414 76412
rect 180536 76452 183554 76480
rect 170732 76372 170738 76384
rect 131850 76304 131856 76356
rect 131908 76344 131914 76356
rect 140590 76344 140596 76356
rect 131908 76316 140596 76344
rect 131908 76304 131914 76316
rect 140590 76304 140596 76316
rect 140648 76304 140654 76356
rect 145466 76304 145472 76356
rect 145524 76344 145530 76356
rect 145926 76344 145932 76356
rect 145524 76316 145932 76344
rect 145524 76304 145530 76316
rect 145926 76304 145932 76316
rect 145984 76304 145990 76356
rect 170766 76304 170772 76356
rect 170824 76344 170830 76356
rect 180536 76344 180564 76452
rect 183526 76412 183554 76452
rect 187326 76412 187332 76424
rect 183526 76384 187332 76412
rect 187326 76372 187332 76384
rect 187384 76372 187390 76424
rect 170824 76316 180564 76344
rect 170824 76304 170830 76316
rect 180702 76304 180708 76356
rect 180760 76344 180766 76356
rect 200758 76344 200764 76356
rect 180760 76316 200764 76344
rect 180760 76304 180766 76316
rect 200758 76304 200764 76316
rect 200816 76304 200822 76356
rect 177022 76168 177028 76220
rect 177080 76208 177086 76220
rect 177942 76208 177948 76220
rect 177080 76180 177948 76208
rect 177080 76168 177086 76180
rect 177942 76168 177948 76180
rect 178000 76168 178006 76220
rect 170122 76100 170128 76152
rect 170180 76140 170186 76152
rect 170674 76140 170680 76152
rect 170180 76112 170680 76140
rect 170180 76100 170186 76112
rect 170674 76100 170680 76112
rect 170732 76100 170738 76152
rect 124858 76032 124864 76084
rect 124916 76072 124922 76084
rect 125594 76072 125600 76084
rect 124916 76044 125600 76072
rect 124916 76032 124922 76044
rect 125594 76032 125600 76044
rect 125652 76032 125658 76084
rect 171226 76032 171232 76084
rect 171284 76072 171290 76084
rect 171594 76072 171600 76084
rect 171284 76044 171600 76072
rect 171284 76032 171290 76044
rect 171594 76032 171600 76044
rect 171652 76032 171658 76084
rect 172790 76032 172796 76084
rect 172848 76072 172854 76084
rect 177206 76072 177212 76084
rect 172848 76044 177212 76072
rect 172848 76032 172854 76044
rect 177206 76032 177212 76044
rect 177264 76032 177270 76084
rect 171778 75964 171784 76016
rect 171836 76004 171842 76016
rect 179874 76004 179880 76016
rect 171836 75976 179880 76004
rect 171836 75964 171842 75976
rect 179874 75964 179880 75976
rect 179932 76004 179938 76016
rect 289814 76004 289820 76016
rect 179932 75976 289820 76004
rect 179932 75964 179938 75976
rect 289814 75964 289820 75976
rect 289872 75964 289878 76016
rect 167914 75896 167920 75948
rect 167972 75936 167978 75948
rect 168282 75936 168288 75948
rect 167972 75908 168288 75936
rect 167972 75896 167978 75908
rect 168282 75896 168288 75908
rect 168340 75896 168346 75948
rect 168926 75896 168932 75948
rect 168984 75936 168990 75948
rect 169570 75936 169576 75948
rect 168984 75908 169576 75936
rect 168984 75896 168990 75908
rect 169570 75896 169576 75908
rect 169628 75896 169634 75948
rect 169846 75896 169852 75948
rect 169904 75936 169910 75948
rect 170582 75936 170588 75948
rect 169904 75908 170588 75936
rect 169904 75896 169910 75908
rect 170582 75896 170588 75908
rect 170640 75896 170646 75948
rect 177758 75896 177764 75948
rect 177816 75936 177822 75948
rect 181346 75936 181352 75948
rect 177816 75908 181352 75936
rect 177816 75896 177822 75908
rect 181346 75896 181352 75908
rect 181404 75936 181410 75948
rect 296714 75936 296720 75948
rect 181404 75908 296720 75936
rect 181404 75896 181410 75908
rect 296714 75896 296720 75908
rect 296772 75896 296778 75948
rect 111518 75828 111524 75880
rect 111576 75868 111582 75880
rect 145466 75868 145472 75880
rect 111576 75840 145472 75868
rect 111576 75828 111582 75840
rect 145466 75828 145472 75840
rect 145524 75828 145530 75880
rect 167546 75828 167552 75880
rect 167604 75868 167610 75880
rect 202322 75868 202328 75880
rect 167604 75840 202328 75868
rect 167604 75828 167610 75840
rect 202322 75828 202328 75840
rect 202380 75828 202386 75880
rect 115382 75760 115388 75812
rect 115440 75800 115446 75812
rect 115440 75772 140774 75800
rect 115440 75760 115446 75772
rect 96614 75692 96620 75744
rect 96672 75732 96678 75744
rect 105814 75732 105820 75744
rect 96672 75704 105820 75732
rect 96672 75692 96678 75704
rect 105814 75692 105820 75704
rect 105872 75732 105878 75744
rect 139670 75732 139676 75744
rect 105872 75704 139676 75732
rect 105872 75692 105878 75704
rect 139670 75692 139676 75704
rect 139728 75692 139734 75744
rect 130746 75624 130752 75676
rect 130804 75664 130810 75676
rect 131022 75664 131028 75676
rect 130804 75636 131028 75664
rect 130804 75624 130810 75636
rect 131022 75624 131028 75636
rect 131080 75624 131086 75676
rect 134242 75624 134248 75676
rect 134300 75664 134306 75676
rect 134702 75664 134708 75676
rect 134300 75636 134708 75664
rect 134300 75624 134306 75636
rect 134702 75624 134708 75636
rect 134760 75624 134766 75676
rect 135438 75624 135444 75676
rect 135496 75664 135502 75676
rect 136450 75664 136456 75676
rect 135496 75636 136456 75664
rect 135496 75624 135502 75636
rect 136450 75624 136456 75636
rect 136508 75624 136514 75676
rect 107010 75556 107016 75608
rect 107068 75596 107074 75608
rect 139118 75596 139124 75608
rect 107068 75568 139124 75596
rect 107068 75556 107074 75568
rect 139118 75556 139124 75568
rect 139176 75556 139182 75608
rect 140746 75596 140774 75772
rect 156414 75760 156420 75812
rect 156472 75800 156478 75812
rect 156874 75800 156880 75812
rect 156472 75772 156880 75800
rect 156472 75760 156478 75772
rect 156874 75760 156880 75772
rect 156932 75760 156938 75812
rect 161658 75760 161664 75812
rect 161716 75800 161722 75812
rect 162762 75800 162768 75812
rect 161716 75772 162768 75800
rect 161716 75760 161722 75772
rect 162762 75760 162768 75772
rect 162820 75800 162826 75812
rect 196342 75800 196348 75812
rect 162820 75772 196348 75800
rect 162820 75760 162826 75772
rect 196342 75760 196348 75772
rect 196400 75760 196406 75812
rect 146294 75692 146300 75744
rect 146352 75732 146358 75744
rect 180794 75732 180800 75744
rect 146352 75704 180800 75732
rect 146352 75692 146358 75704
rect 180794 75692 180800 75704
rect 180852 75692 180858 75744
rect 146754 75624 146760 75676
rect 146812 75664 146818 75676
rect 185026 75664 185032 75676
rect 146812 75636 185032 75664
rect 146812 75624 146818 75636
rect 185026 75624 185032 75636
rect 185084 75624 185090 75676
rect 140746 75568 147766 75596
rect 117222 75488 117228 75540
rect 117280 75528 117286 75540
rect 145374 75528 145380 75540
rect 117280 75500 145380 75528
rect 117280 75488 117286 75500
rect 145374 75488 145380 75500
rect 145432 75488 145438 75540
rect 147738 75528 147766 75568
rect 147858 75556 147864 75608
rect 147916 75596 147922 75608
rect 198734 75596 198740 75608
rect 147916 75568 198740 75596
rect 147916 75556 147922 75568
rect 198734 75556 198740 75568
rect 198792 75556 198798 75608
rect 147738 75500 148364 75528
rect 121178 75420 121184 75472
rect 121236 75460 121242 75472
rect 148134 75460 148140 75472
rect 121236 75432 148140 75460
rect 121236 75420 121242 75432
rect 148134 75420 148140 75432
rect 148192 75420 148198 75472
rect 148336 75460 148364 75500
rect 150158 75488 150164 75540
rect 150216 75528 150222 75540
rect 216674 75528 216680 75540
rect 150216 75500 216680 75528
rect 150216 75488 150222 75500
rect 216674 75488 216680 75500
rect 216732 75488 216738 75540
rect 149606 75460 149612 75472
rect 148336 75432 149612 75460
rect 149606 75420 149612 75432
rect 149664 75460 149670 75472
rect 223574 75460 223580 75472
rect 149664 75432 223580 75460
rect 149664 75420 149670 75432
rect 223574 75420 223580 75432
rect 223632 75420 223638 75472
rect 122742 75352 122748 75404
rect 122800 75392 122806 75404
rect 149882 75392 149888 75404
rect 122800 75364 149888 75392
rect 122800 75352 122806 75364
rect 149882 75352 149888 75364
rect 149940 75352 149946 75404
rect 165706 75352 165712 75404
rect 165764 75392 165770 75404
rect 165982 75392 165988 75404
rect 165764 75364 165988 75392
rect 165764 75352 165770 75364
rect 165982 75352 165988 75364
rect 166040 75352 166046 75404
rect 167546 75352 167552 75404
rect 167604 75392 167610 75404
rect 168006 75392 168012 75404
rect 167604 75364 168012 75392
rect 167604 75352 167610 75364
rect 168006 75352 168012 75364
rect 168064 75352 168070 75404
rect 171502 75352 171508 75404
rect 171560 75392 171566 75404
rect 171560 75364 172100 75392
rect 171560 75352 171566 75364
rect 118602 75284 118608 75336
rect 118660 75324 118666 75336
rect 145558 75324 145564 75336
rect 118660 75296 145564 75324
rect 118660 75284 118666 75296
rect 145558 75284 145564 75296
rect 145616 75284 145622 75336
rect 156046 75284 156052 75336
rect 156104 75324 156110 75336
rect 156782 75324 156788 75336
rect 156104 75296 156788 75324
rect 156104 75284 156110 75296
rect 156782 75284 156788 75296
rect 156840 75284 156846 75336
rect 160462 75284 160468 75336
rect 160520 75324 160526 75336
rect 162026 75324 162032 75336
rect 160520 75296 162032 75324
rect 160520 75284 160526 75296
rect 162026 75284 162032 75296
rect 162084 75284 162090 75336
rect 166074 75284 166080 75336
rect 166132 75324 166138 75336
rect 171962 75324 171968 75336
rect 166132 75296 171968 75324
rect 166132 75284 166138 75296
rect 171962 75284 171968 75296
rect 172020 75284 172026 75336
rect 172072 75324 172100 75364
rect 174170 75352 174176 75404
rect 174228 75392 174234 75404
rect 504358 75392 504364 75404
rect 174228 75364 504364 75392
rect 174228 75352 174234 75364
rect 504358 75352 504364 75364
rect 504416 75352 504422 75404
rect 454678 75324 454684 75336
rect 172072 75296 454684 75324
rect 454678 75284 454684 75296
rect 454736 75284 454742 75336
rect 81434 75216 81440 75268
rect 81492 75256 81498 75268
rect 138658 75256 138664 75268
rect 81492 75228 138664 75256
rect 81492 75216 81498 75228
rect 138658 75216 138664 75228
rect 138716 75216 138722 75268
rect 145374 75216 145380 75268
rect 145432 75256 145438 75268
rect 145742 75256 145748 75268
rect 145432 75228 145748 75256
rect 145432 75216 145438 75228
rect 145742 75216 145748 75228
rect 145800 75216 145806 75268
rect 166994 75216 167000 75268
rect 167052 75256 167058 75268
rect 168098 75256 168104 75268
rect 167052 75228 168104 75256
rect 167052 75216 167058 75228
rect 168098 75216 168104 75228
rect 168156 75216 168162 75268
rect 172882 75216 172888 75268
rect 172940 75256 172946 75268
rect 173710 75256 173716 75268
rect 172940 75228 173716 75256
rect 172940 75216 172946 75228
rect 173710 75216 173716 75228
rect 173768 75216 173774 75268
rect 174354 75216 174360 75268
rect 174412 75256 174418 75268
rect 511258 75256 511264 75268
rect 174412 75228 511264 75256
rect 174412 75216 174418 75228
rect 511258 75216 511264 75228
rect 511316 75216 511322 75268
rect 67634 75148 67640 75200
rect 67692 75188 67698 75200
rect 132586 75188 132592 75200
rect 67692 75160 132592 75188
rect 67692 75148 67698 75160
rect 132586 75148 132592 75160
rect 132644 75148 132650 75200
rect 132678 75148 132684 75200
rect 132736 75188 132742 75200
rect 133782 75188 133788 75200
rect 132736 75160 133788 75188
rect 132736 75148 132742 75160
rect 133782 75148 133788 75160
rect 133840 75148 133846 75200
rect 135806 75148 135812 75200
rect 135864 75188 135870 75200
rect 136542 75188 136548 75200
rect 135864 75160 136548 75188
rect 135864 75148 135870 75160
rect 136542 75148 136548 75160
rect 136600 75148 136606 75200
rect 136634 75148 136640 75200
rect 136692 75188 136698 75200
rect 137186 75188 137192 75200
rect 136692 75160 137192 75188
rect 136692 75148 136698 75160
rect 137186 75148 137192 75160
rect 137244 75148 137250 75200
rect 168650 75148 168656 75200
rect 168708 75188 168714 75200
rect 169110 75188 169116 75200
rect 168708 75160 169116 75188
rect 168708 75148 168714 75160
rect 169110 75148 169116 75160
rect 169168 75148 169174 75200
rect 172974 75148 172980 75200
rect 173032 75188 173038 75200
rect 521654 75188 521660 75200
rect 173032 75160 521660 75188
rect 173032 75148 173038 75160
rect 521654 75148 521660 75160
rect 521712 75148 521718 75200
rect 115934 75080 115940 75132
rect 115992 75120 115998 75132
rect 116486 75120 116492 75132
rect 115992 75092 116492 75120
rect 115992 75080 115998 75092
rect 116486 75080 116492 75092
rect 116544 75120 116550 75132
rect 141326 75120 141332 75132
rect 116544 75092 141332 75120
rect 116544 75080 116550 75092
rect 141326 75080 141332 75092
rect 141384 75080 141390 75132
rect 157518 75080 157524 75132
rect 157576 75120 157582 75132
rect 189902 75120 189908 75132
rect 157576 75092 189908 75120
rect 157576 75080 157582 75092
rect 189902 75080 189908 75092
rect 189960 75080 189966 75132
rect 114462 75012 114468 75064
rect 114520 75052 114526 75064
rect 147214 75052 147220 75064
rect 114520 75024 147220 75052
rect 114520 75012 114526 75024
rect 147214 75012 147220 75024
rect 147272 75012 147278 75064
rect 159818 75012 159824 75064
rect 159876 75052 159882 75064
rect 160002 75052 160008 75064
rect 159876 75024 160008 75052
rect 159876 75012 159882 75024
rect 160002 75012 160008 75024
rect 160060 75012 160066 75064
rect 164786 75012 164792 75064
rect 164844 75052 164850 75064
rect 192478 75052 192484 75064
rect 164844 75024 192484 75052
rect 164844 75012 164850 75024
rect 192478 75012 192484 75024
rect 192536 75012 192542 75064
rect 134334 74944 134340 74996
rect 134392 74984 134398 74996
rect 135162 74984 135168 74996
rect 134392 74956 135168 74984
rect 134392 74944 134398 74956
rect 135162 74944 135168 74956
rect 135220 74944 135226 74996
rect 135438 74944 135444 74996
rect 135496 74984 135502 74996
rect 136266 74984 136272 74996
rect 135496 74956 136272 74984
rect 135496 74944 135502 74956
rect 136266 74944 136272 74956
rect 136324 74944 136330 74996
rect 173710 74944 173716 74996
rect 173768 74984 173774 74996
rect 198366 74984 198372 74996
rect 173768 74956 198372 74984
rect 173768 74944 173774 74956
rect 198366 74944 198372 74956
rect 198424 74944 198430 74996
rect 132586 74876 132592 74928
rect 132644 74916 132650 74928
rect 137646 74916 137652 74928
rect 132644 74888 137652 74916
rect 132644 74876 132650 74888
rect 137646 74876 137652 74888
rect 137704 74876 137710 74928
rect 158806 74876 158812 74928
rect 158864 74916 158870 74928
rect 159818 74916 159824 74928
rect 158864 74888 159824 74916
rect 158864 74876 158870 74888
rect 159818 74876 159824 74888
rect 159876 74876 159882 74928
rect 176838 74876 176844 74928
rect 176896 74916 176902 74928
rect 177758 74916 177764 74928
rect 176896 74888 177764 74916
rect 176896 74876 176902 74888
rect 177758 74876 177764 74888
rect 177816 74876 177822 74928
rect 129918 74672 129924 74724
rect 129976 74712 129982 74724
rect 142154 74712 142160 74724
rect 129976 74684 142160 74712
rect 129976 74672 129982 74684
rect 142154 74672 142160 74684
rect 142212 74672 142218 74724
rect 158898 74604 158904 74656
rect 158956 74644 158962 74656
rect 159450 74644 159456 74656
rect 158956 74616 159456 74644
rect 158956 74604 158962 74616
rect 159450 74604 159456 74616
rect 159508 74604 159514 74656
rect 168558 74604 168564 74656
rect 168616 74644 168622 74656
rect 169202 74644 169208 74656
rect 168616 74616 169208 74644
rect 168616 74604 168622 74616
rect 169202 74604 169208 74616
rect 169260 74604 169266 74656
rect 111150 74468 111156 74520
rect 111208 74508 111214 74520
rect 143534 74508 143540 74520
rect 111208 74480 143540 74508
rect 111208 74468 111214 74480
rect 143534 74468 143540 74480
rect 143592 74468 143598 74520
rect 143718 74468 143724 74520
rect 143776 74508 143782 74520
rect 144086 74508 144092 74520
rect 143776 74480 144092 74508
rect 143776 74468 143782 74480
rect 144086 74468 144092 74480
rect 144144 74468 144150 74520
rect 145006 74468 145012 74520
rect 145064 74508 145070 74520
rect 145374 74508 145380 74520
rect 145064 74480 145380 74508
rect 145064 74468 145070 74480
rect 145374 74468 145380 74480
rect 145432 74468 145438 74520
rect 161014 74468 161020 74520
rect 161072 74508 161078 74520
rect 161474 74508 161480 74520
rect 161072 74480 161480 74508
rect 161072 74468 161078 74480
rect 161474 74468 161480 74480
rect 161532 74468 161538 74520
rect 165890 74468 165896 74520
rect 165948 74508 165954 74520
rect 166810 74508 166816 74520
rect 165948 74480 166816 74508
rect 165948 74468 165954 74480
rect 166810 74468 166816 74480
rect 166868 74508 166874 74520
rect 200850 74508 200856 74520
rect 166868 74480 200856 74508
rect 166868 74468 166874 74480
rect 200850 74468 200856 74480
rect 200908 74468 200914 74520
rect 111702 74400 111708 74452
rect 111760 74440 111766 74452
rect 144270 74440 144276 74452
rect 111760 74412 144276 74440
rect 111760 74400 111766 74412
rect 144270 74400 144276 74412
rect 144328 74400 144334 74452
rect 168742 74400 168748 74452
rect 168800 74440 168806 74452
rect 202046 74440 202052 74452
rect 168800 74412 202052 74440
rect 168800 74400 168806 74412
rect 202046 74400 202052 74412
rect 202104 74400 202110 74452
rect 120350 74332 120356 74384
rect 120408 74372 120414 74384
rect 152090 74372 152096 74384
rect 120408 74344 152096 74372
rect 120408 74332 120414 74344
rect 152090 74332 152096 74344
rect 152148 74332 152154 74384
rect 160554 74332 160560 74384
rect 160612 74372 160618 74384
rect 161290 74372 161296 74384
rect 160612 74344 161296 74372
rect 160612 74332 160618 74344
rect 161290 74332 161296 74344
rect 161348 74372 161354 74384
rect 193858 74372 193864 74384
rect 161348 74344 193864 74372
rect 161348 74332 161354 74344
rect 193858 74332 193864 74344
rect 193916 74332 193922 74384
rect 108298 74264 108304 74316
rect 108356 74304 108362 74316
rect 140682 74304 140688 74316
rect 108356 74276 140688 74304
rect 108356 74264 108362 74276
rect 140682 74264 140688 74276
rect 140740 74264 140746 74316
rect 150250 74264 150256 74316
rect 150308 74304 150314 74316
rect 203610 74304 203616 74316
rect 150308 74276 203616 74304
rect 150308 74264 150314 74276
rect 203610 74264 203616 74276
rect 203668 74264 203674 74316
rect 114094 74196 114100 74248
rect 114152 74236 114158 74248
rect 145006 74236 145012 74248
rect 114152 74208 145012 74236
rect 114152 74196 114158 74208
rect 145006 74196 145012 74208
rect 145064 74196 145070 74248
rect 150894 74196 150900 74248
rect 150952 74236 150958 74248
rect 237374 74236 237380 74248
rect 150952 74208 237380 74236
rect 150952 74196 150958 74208
rect 237374 74196 237380 74208
rect 237432 74196 237438 74248
rect 112714 74128 112720 74180
rect 112772 74168 112778 74180
rect 143718 74168 143724 74180
rect 112772 74140 143724 74168
rect 112772 74128 112778 74140
rect 143718 74128 143724 74140
rect 143776 74128 143782 74180
rect 151722 74128 151728 74180
rect 151780 74168 151786 74180
rect 247678 74168 247684 74180
rect 151780 74140 247684 74168
rect 151780 74128 151786 74140
rect 247678 74128 247684 74140
rect 247736 74128 247742 74180
rect 117958 74060 117964 74112
rect 118016 74100 118022 74112
rect 148042 74100 148048 74112
rect 118016 74072 148048 74100
rect 118016 74060 118022 74072
rect 148042 74060 148048 74072
rect 148100 74060 148106 74112
rect 154206 74060 154212 74112
rect 154264 74100 154270 74112
rect 284294 74100 284300 74112
rect 154264 74072 284300 74100
rect 154264 74060 154270 74072
rect 284294 74060 284300 74072
rect 284352 74060 284358 74112
rect 112990 73992 112996 74044
rect 113048 74032 113054 74044
rect 142430 74032 142436 74044
rect 113048 74004 142436 74032
rect 113048 73992 113054 74004
rect 142430 73992 142436 74004
rect 142488 73992 142494 74044
rect 157518 73992 157524 74044
rect 157576 74032 157582 74044
rect 158254 74032 158260 74044
rect 157576 74004 158260 74032
rect 157576 73992 157582 74004
rect 158254 73992 158260 74004
rect 158312 73992 158318 74044
rect 159358 73992 159364 74044
rect 159416 74032 159422 74044
rect 347774 74032 347780 74044
rect 159416 74004 347780 74032
rect 159416 73992 159422 74004
rect 347774 73992 347780 74004
rect 347832 73992 347838 74044
rect 113450 73924 113456 73976
rect 113508 73964 113514 73976
rect 138566 73964 138572 73976
rect 113508 73936 138572 73964
rect 113508 73924 113514 73936
rect 138566 73924 138572 73936
rect 138624 73924 138630 73976
rect 141602 73924 141608 73976
rect 141660 73964 141666 73976
rect 141970 73964 141976 73976
rect 141660 73936 141976 73964
rect 141660 73924 141666 73936
rect 141970 73924 141976 73936
rect 142028 73924 142034 73976
rect 152182 73924 152188 73976
rect 152240 73964 152246 73976
rect 255314 73964 255320 73976
rect 152240 73936 255320 73964
rect 152240 73924 152246 73936
rect 255314 73924 255320 73936
rect 255372 73924 255378 73976
rect 255958 73924 255964 73976
rect 256016 73964 256022 73976
rect 456794 73964 456800 73976
rect 256016 73936 456800 73964
rect 256016 73924 256022 73936
rect 456794 73924 456800 73936
rect 456852 73924 456858 73976
rect 95234 73856 95240 73908
rect 95292 73896 95298 73908
rect 140038 73896 140044 73908
rect 95292 73868 140044 73896
rect 95292 73856 95298 73868
rect 140038 73856 140044 73868
rect 140096 73856 140102 73908
rect 157334 73856 157340 73908
rect 157392 73896 157398 73908
rect 158346 73896 158352 73908
rect 157392 73868 158352 73896
rect 157392 73856 157398 73868
rect 158346 73856 158352 73868
rect 158404 73856 158410 73908
rect 172422 73856 172428 73908
rect 172480 73896 172486 73908
rect 190178 73896 190184 73908
rect 172480 73868 190184 73896
rect 172480 73856 172486 73868
rect 190178 73856 190184 73868
rect 190236 73856 190242 73908
rect 202046 73856 202052 73908
rect 202104 73896 202110 73908
rect 446398 73896 446404 73908
rect 202104 73868 446404 73896
rect 202104 73856 202110 73868
rect 446398 73856 446404 73868
rect 446456 73856 446462 73908
rect 54478 73788 54484 73840
rect 54536 73828 54542 73840
rect 107378 73828 107384 73840
rect 54536 73800 107384 73828
rect 54536 73788 54542 73800
rect 107378 73788 107384 73800
rect 107436 73788 107442 73840
rect 115198 73788 115204 73840
rect 115256 73828 115262 73840
rect 138382 73828 138388 73840
rect 115256 73800 138388 73828
rect 115256 73788 115262 73800
rect 138382 73788 138388 73800
rect 138440 73788 138446 73840
rect 143534 73788 143540 73840
rect 143592 73828 143598 73840
rect 144178 73828 144184 73840
rect 143592 73800 144184 73828
rect 143592 73788 143598 73800
rect 144178 73788 144184 73800
rect 144236 73828 144242 73840
rect 152182 73828 152188 73840
rect 144236 73800 152188 73828
rect 144236 73788 144242 73800
rect 152182 73788 152188 73800
rect 152240 73788 152246 73840
rect 152918 73788 152924 73840
rect 152976 73828 152982 73840
rect 261478 73828 261484 73840
rect 152976 73800 261484 73828
rect 152976 73788 152982 73800
rect 261478 73788 261484 73800
rect 261536 73788 261542 73840
rect 264238 73788 264244 73840
rect 264296 73828 264302 73840
rect 518894 73828 518900 73840
rect 264296 73800 518900 73828
rect 264296 73788 264302 73800
rect 518894 73788 518900 73800
rect 518952 73788 518958 73840
rect 117682 73720 117688 73772
rect 117740 73760 117746 73772
rect 129734 73760 129740 73772
rect 117740 73732 129740 73760
rect 117740 73720 117746 73732
rect 129734 73720 129740 73732
rect 129792 73760 129798 73772
rect 132954 73760 132960 73772
rect 129792 73732 132960 73760
rect 129792 73720 129798 73732
rect 132954 73720 132960 73732
rect 133012 73720 133018 73772
rect 176194 73720 176200 73772
rect 176252 73760 176258 73772
rect 204622 73760 204628 73772
rect 176252 73732 204628 73760
rect 176252 73720 176258 73732
rect 204622 73720 204628 73732
rect 204680 73720 204686 73772
rect 169386 73652 169392 73704
rect 169444 73692 169450 73704
rect 180242 73692 180248 73704
rect 169444 73664 180248 73692
rect 169444 73652 169450 73664
rect 180242 73652 180248 73664
rect 180300 73652 180306 73704
rect 107378 73584 107384 73636
rect 107436 73624 107442 73636
rect 136358 73624 136364 73636
rect 107436 73596 136364 73624
rect 107436 73584 107442 73596
rect 136358 73584 136364 73596
rect 136416 73584 136422 73636
rect 158990 73244 158996 73296
rect 159048 73284 159054 73296
rect 159174 73284 159180 73296
rect 159048 73256 159180 73284
rect 159048 73244 159054 73256
rect 159174 73244 159180 73256
rect 159232 73244 159238 73296
rect 107654 73176 107660 73228
rect 107712 73216 107718 73228
rect 108298 73216 108304 73228
rect 107712 73188 108304 73216
rect 107712 73176 107718 73188
rect 108298 73176 108304 73188
rect 108356 73176 108362 73228
rect 124950 73176 124956 73228
rect 125008 73216 125014 73228
rect 125686 73216 125692 73228
rect 125008 73188 125692 73216
rect 125008 73176 125014 73188
rect 125686 73176 125692 73188
rect 125744 73176 125750 73228
rect 142448 73188 143212 73216
rect 105906 73108 105912 73160
rect 105964 73148 105970 73160
rect 139578 73148 139584 73160
rect 105964 73120 139584 73148
rect 105964 73108 105970 73120
rect 139578 73108 139584 73120
rect 139636 73148 139642 73160
rect 140498 73148 140504 73160
rect 139636 73120 140504 73148
rect 139636 73108 139642 73120
rect 140498 73108 140504 73120
rect 140556 73108 140562 73160
rect 142448 73148 142476 73188
rect 142172 73120 142476 73148
rect 143184 73148 143212 73188
rect 146662 73148 146668 73160
rect 143184 73120 146668 73148
rect 114278 73040 114284 73092
rect 114336 73080 114342 73092
rect 142172 73080 142200 73120
rect 146662 73108 146668 73120
rect 146720 73108 146726 73160
rect 164694 73108 164700 73160
rect 164752 73148 164758 73160
rect 165246 73148 165252 73160
rect 164752 73120 165252 73148
rect 164752 73108 164758 73120
rect 165246 73108 165252 73120
rect 165304 73148 165310 73160
rect 199470 73148 199476 73160
rect 165304 73120 199476 73148
rect 165304 73108 165310 73120
rect 199470 73108 199476 73120
rect 199528 73108 199534 73160
rect 327718 73108 327724 73160
rect 327776 73148 327782 73160
rect 579982 73148 579988 73160
rect 327776 73120 579988 73148
rect 327776 73108 327782 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 114336 73052 142200 73080
rect 114336 73040 114342 73052
rect 142246 73040 142252 73092
rect 142304 73080 142310 73092
rect 143442 73080 143448 73092
rect 142304 73052 143448 73080
rect 142304 73040 142310 73052
rect 143442 73040 143448 73052
rect 143500 73040 143506 73092
rect 157058 73040 157064 73092
rect 157116 73080 157122 73092
rect 191006 73080 191012 73092
rect 157116 73052 191012 73080
rect 157116 73040 157122 73052
rect 191006 73040 191012 73052
rect 191064 73040 191070 73092
rect 121270 72972 121276 73024
rect 121328 73012 121334 73024
rect 153746 73012 153752 73024
rect 121328 72984 138014 73012
rect 121328 72972 121334 72984
rect 100202 72904 100208 72956
rect 100260 72944 100266 72956
rect 133598 72944 133604 72956
rect 100260 72916 133604 72944
rect 100260 72904 100266 72916
rect 133598 72904 133604 72916
rect 133656 72904 133662 72956
rect 137986 72944 138014 72984
rect 142264 72984 153752 73012
rect 142264 72944 142292 72984
rect 153746 72972 153752 72984
rect 153804 72972 153810 73024
rect 156506 72972 156512 73024
rect 156564 73012 156570 73024
rect 187050 73012 187056 73024
rect 156564 72984 187056 73012
rect 156564 72972 156570 72984
rect 187050 72972 187056 72984
rect 187108 73012 187114 73024
rect 187602 73012 187608 73024
rect 187108 72984 187608 73012
rect 187108 72972 187114 72984
rect 187602 72972 187608 72984
rect 187660 72972 187666 73024
rect 137986 72916 142292 72944
rect 154850 72904 154856 72956
rect 154908 72944 154914 72956
rect 242158 72944 242164 72956
rect 154908 72916 242164 72944
rect 154908 72904 154914 72916
rect 242158 72904 242164 72916
rect 242216 72904 242222 72956
rect 122650 72836 122656 72888
rect 122708 72876 122714 72888
rect 154022 72876 154028 72888
rect 122708 72848 154028 72876
rect 122708 72836 122714 72848
rect 154022 72836 154028 72848
rect 154080 72836 154086 72888
rect 160094 72836 160100 72888
rect 160152 72876 160158 72888
rect 160738 72876 160744 72888
rect 160152 72848 160744 72876
rect 160152 72836 160158 72848
rect 160738 72836 160744 72848
rect 160796 72876 160802 72888
rect 189810 72876 189816 72888
rect 160796 72848 189816 72876
rect 160796 72836 160802 72848
rect 189810 72836 189816 72848
rect 189868 72836 189874 72888
rect 191006 72836 191012 72888
rect 191064 72876 191070 72888
rect 301498 72876 301504 72888
rect 191064 72848 301504 72876
rect 191064 72836 191070 72848
rect 301498 72836 301504 72848
rect 301556 72836 301562 72888
rect 104342 72768 104348 72820
rect 104400 72808 104406 72820
rect 135254 72808 135260 72820
rect 104400 72780 135260 72808
rect 104400 72768 104406 72780
rect 135254 72768 135260 72780
rect 135312 72768 135318 72820
rect 187602 72768 187608 72820
rect 187660 72808 187666 72820
rect 304994 72808 305000 72820
rect 187660 72780 305000 72808
rect 187660 72768 187666 72780
rect 304994 72768 305000 72780
rect 305052 72768 305058 72820
rect 111426 72700 111432 72752
rect 111484 72740 111490 72752
rect 142890 72740 142896 72752
rect 111484 72712 142896 72740
rect 111484 72700 111490 72712
rect 142890 72700 142896 72712
rect 142948 72700 142954 72752
rect 156966 72700 156972 72752
rect 157024 72740 157030 72752
rect 311158 72740 311164 72752
rect 157024 72712 311164 72740
rect 157024 72700 157030 72712
rect 311158 72700 311164 72712
rect 311216 72700 311222 72752
rect 111610 72632 111616 72684
rect 111668 72672 111674 72684
rect 142246 72672 142252 72684
rect 111668 72644 142252 72672
rect 111668 72632 111674 72644
rect 142246 72632 142252 72644
rect 142304 72632 142310 72684
rect 157426 72632 157432 72684
rect 157484 72672 157490 72684
rect 318794 72672 318800 72684
rect 157484 72644 318800 72672
rect 157484 72632 157490 72644
rect 318794 72632 318800 72644
rect 318852 72632 318858 72684
rect 70394 72564 70400 72616
rect 70452 72604 70458 72616
rect 137922 72604 137928 72616
rect 70452 72576 137928 72604
rect 70452 72564 70458 72576
rect 137922 72564 137928 72576
rect 137980 72564 137986 72616
rect 153286 72564 153292 72616
rect 153344 72604 153350 72616
rect 153654 72604 153660 72616
rect 153344 72576 153660 72604
rect 153344 72564 153350 72576
rect 153654 72564 153660 72576
rect 153712 72564 153718 72616
rect 157702 72564 157708 72616
rect 157760 72604 157766 72616
rect 324958 72604 324964 72616
rect 157760 72576 324964 72604
rect 157760 72564 157766 72576
rect 324958 72564 324964 72576
rect 325016 72564 325022 72616
rect 21358 72496 21364 72548
rect 21416 72536 21422 72548
rect 100202 72536 100208 72548
rect 21416 72508 100208 72536
rect 21416 72496 21422 72508
rect 100202 72496 100208 72508
rect 100260 72496 100266 72548
rect 112898 72496 112904 72548
rect 112956 72536 112962 72548
rect 142522 72536 142528 72548
rect 112956 72508 142528 72536
rect 112956 72496 112962 72508
rect 142522 72496 142528 72508
rect 142580 72496 142586 72548
rect 157794 72496 157800 72548
rect 157852 72536 157858 72548
rect 332594 72536 332600 72548
rect 157852 72508 332600 72536
rect 157852 72496 157858 72508
rect 332594 72496 332600 72508
rect 332652 72496 332658 72548
rect 45554 72428 45560 72480
rect 45612 72468 45618 72480
rect 135530 72468 135536 72480
rect 45612 72440 135536 72468
rect 45612 72428 45618 72440
rect 135530 72428 135536 72440
rect 135588 72428 135594 72480
rect 145650 72428 145656 72480
rect 145708 72468 145714 72480
rect 156322 72468 156328 72480
rect 145708 72440 156328 72468
rect 145708 72428 145714 72440
rect 156322 72428 156328 72440
rect 156380 72428 156386 72480
rect 167454 72428 167460 72480
rect 167512 72468 167518 72480
rect 375374 72468 375380 72480
rect 167512 72440 375380 72468
rect 167512 72428 167518 72440
rect 375374 72428 375380 72440
rect 375432 72428 375438 72480
rect 119798 72360 119804 72412
rect 119856 72400 119862 72412
rect 141510 72400 141516 72412
rect 119856 72372 141516 72400
rect 119856 72360 119862 72372
rect 141510 72360 141516 72372
rect 141568 72360 141574 72412
rect 146662 72360 146668 72412
rect 146720 72400 146726 72412
rect 147398 72400 147404 72412
rect 146720 72372 147404 72400
rect 146720 72360 146726 72372
rect 147398 72360 147404 72372
rect 147456 72360 147462 72412
rect 162210 72360 162216 72412
rect 162268 72400 162274 72412
rect 190086 72400 190092 72412
rect 162268 72372 190092 72400
rect 162268 72360 162274 72372
rect 190086 72360 190092 72372
rect 190144 72360 190150 72412
rect 121362 72292 121368 72344
rect 121420 72332 121426 72344
rect 129918 72332 129924 72344
rect 121420 72304 129924 72332
rect 121420 72292 121426 72304
rect 129918 72292 129924 72304
rect 129976 72292 129982 72344
rect 135254 72292 135260 72344
rect 135312 72332 135318 72344
rect 135530 72332 135536 72344
rect 135312 72304 135536 72332
rect 135312 72292 135318 72304
rect 135530 72292 135536 72304
rect 135588 72292 135594 72344
rect 160002 72292 160008 72344
rect 160060 72332 160066 72344
rect 187234 72332 187240 72344
rect 160060 72304 187240 72332
rect 160060 72292 160066 72304
rect 187234 72292 187240 72304
rect 187292 72292 187298 72344
rect 174906 72224 174912 72276
rect 174964 72264 174970 72276
rect 205910 72264 205916 72276
rect 174964 72236 205916 72264
rect 174964 72224 174970 72236
rect 205910 72224 205916 72236
rect 205968 72224 205974 72276
rect 164234 72156 164240 72208
rect 164292 72196 164298 72208
rect 165522 72196 165528 72208
rect 164292 72168 165528 72196
rect 164292 72156 164298 72168
rect 165522 72156 165528 72168
rect 165580 72196 165586 72208
rect 195514 72196 195520 72208
rect 165580 72168 195520 72196
rect 165580 72156 165586 72168
rect 195514 72156 195520 72168
rect 195572 72156 195578 72208
rect 148042 72088 148048 72140
rect 148100 72128 148106 72140
rect 148778 72128 148784 72140
rect 148100 72100 148784 72128
rect 148100 72088 148106 72100
rect 148778 72088 148784 72100
rect 148836 72088 148842 72140
rect 152090 72088 152096 72140
rect 152148 72128 152154 72140
rect 152826 72128 152832 72140
rect 152148 72100 152832 72128
rect 152148 72088 152154 72100
rect 152826 72088 152832 72100
rect 152884 72088 152890 72140
rect 164234 72020 164240 72072
rect 164292 72060 164298 72072
rect 164602 72060 164608 72072
rect 164292 72032 164608 72060
rect 164292 72020 164298 72032
rect 164602 72020 164608 72032
rect 164660 72020 164666 72072
rect 161842 71952 161848 72004
rect 161900 71992 161906 72004
rect 162394 71992 162400 72004
rect 161900 71964 162400 71992
rect 161900 71952 161906 71964
rect 162394 71952 162400 71964
rect 162452 71952 162458 72004
rect 166350 71816 166356 71868
rect 166408 71856 166414 71868
rect 166902 71856 166908 71868
rect 166408 71828 166908 71856
rect 166408 71816 166414 71828
rect 166902 71816 166908 71828
rect 166960 71816 166966 71868
rect 118694 71748 118700 71800
rect 118752 71788 118758 71800
rect 119798 71788 119804 71800
rect 118752 71760 119804 71788
rect 118752 71748 118758 71760
rect 119798 71748 119804 71760
rect 119856 71748 119862 71800
rect 163958 71748 163964 71800
rect 164016 71788 164022 71800
rect 164016 71760 166994 71788
rect 164016 71748 164022 71760
rect 117590 71680 117596 71732
rect 117648 71720 117654 71732
rect 151814 71720 151820 71732
rect 117648 71692 151820 71720
rect 117648 71680 117654 71692
rect 151814 71680 151820 71692
rect 151872 71680 151878 71732
rect 164326 71680 164332 71732
rect 164384 71720 164390 71732
rect 165430 71720 165436 71732
rect 164384 71692 165436 71720
rect 164384 71680 164390 71692
rect 165430 71680 165436 71692
rect 165488 71680 165494 71732
rect 165982 71680 165988 71732
rect 166040 71720 166046 71732
rect 166350 71720 166356 71732
rect 166040 71692 166356 71720
rect 166040 71680 166046 71692
rect 166350 71680 166356 71692
rect 166408 71680 166414 71732
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 8938 71652 8944 71664
rect 3568 71624 8944 71652
rect 3568 71612 3574 71624
rect 8938 71612 8944 71624
rect 8996 71612 9002 71664
rect 120810 71612 120816 71664
rect 120868 71652 120874 71664
rect 154574 71652 154580 71664
rect 120868 71624 154580 71652
rect 120868 71612 120874 71624
rect 154574 71612 154580 71624
rect 154632 71652 154638 71664
rect 155218 71652 155224 71664
rect 154632 71624 155224 71652
rect 154632 71612 154638 71624
rect 155218 71612 155224 71624
rect 155276 71612 155282 71664
rect 166966 71652 166994 71760
rect 182174 71680 182180 71732
rect 182232 71720 182238 71732
rect 192110 71720 192116 71732
rect 182232 71692 192116 71720
rect 182232 71680 182238 71692
rect 192110 71680 192116 71692
rect 192168 71680 192174 71732
rect 197998 71652 198004 71664
rect 166966 71624 198004 71652
rect 197998 71612 198004 71624
rect 198056 71612 198062 71664
rect 100110 71544 100116 71596
rect 100168 71584 100174 71596
rect 134610 71584 134616 71596
rect 100168 71556 134616 71584
rect 100168 71544 100174 71556
rect 134610 71544 134616 71556
rect 134668 71544 134674 71596
rect 138566 71544 138572 71596
rect 138624 71584 138630 71596
rect 139302 71584 139308 71596
rect 138624 71556 139308 71584
rect 138624 71544 138630 71556
rect 139302 71544 139308 71556
rect 139360 71544 139366 71596
rect 141510 71544 141516 71596
rect 141568 71584 141574 71596
rect 142890 71584 142896 71596
rect 141568 71556 142896 71584
rect 141568 71544 141574 71556
rect 142890 71544 142896 71556
rect 142948 71544 142954 71596
rect 165154 71544 165160 71596
rect 165212 71584 165218 71596
rect 165614 71584 165620 71596
rect 165212 71556 165620 71584
rect 165212 71544 165218 71556
rect 165614 71544 165620 71556
rect 165672 71584 165678 71596
rect 199286 71584 199292 71596
rect 165672 71556 199292 71584
rect 165672 71544 165678 71556
rect 199286 71544 199292 71556
rect 199344 71544 199350 71596
rect 118142 71476 118148 71528
rect 118200 71516 118206 71528
rect 150802 71516 150808 71528
rect 118200 71488 150808 71516
rect 118200 71476 118206 71488
rect 150802 71476 150808 71488
rect 150860 71476 150866 71528
rect 196986 71516 196992 71528
rect 165540 71488 196992 71516
rect 120442 71408 120448 71460
rect 120500 71448 120506 71460
rect 120500 71420 138014 71448
rect 120500 71408 120506 71420
rect 104434 71340 104440 71392
rect 104492 71380 104498 71392
rect 134150 71380 134156 71392
rect 104492 71352 134156 71380
rect 104492 71340 104498 71352
rect 134150 71340 134156 71352
rect 134208 71380 134214 71392
rect 134794 71380 134800 71392
rect 134208 71352 134800 71380
rect 134208 71340 134214 71352
rect 134794 71340 134800 71352
rect 134852 71340 134858 71392
rect 137986 71380 138014 71420
rect 142338 71408 142344 71460
rect 142396 71448 142402 71460
rect 143166 71448 143172 71460
rect 142396 71420 143172 71448
rect 142396 71408 142402 71420
rect 143166 71408 143172 71420
rect 143224 71408 143230 71460
rect 151814 71408 151820 71460
rect 151872 71448 151878 71460
rect 152734 71448 152740 71460
rect 151872 71420 152740 71448
rect 151872 71408 151878 71420
rect 152734 71408 152740 71420
rect 152792 71408 152798 71460
rect 163682 71408 163688 71460
rect 163740 71448 163746 71460
rect 163958 71448 163964 71460
rect 163740 71420 163964 71448
rect 163740 71408 163746 71420
rect 163958 71408 163964 71420
rect 164016 71448 164022 71460
rect 165540 71448 165568 71488
rect 196986 71476 196992 71488
rect 197044 71476 197050 71528
rect 192294 71448 192300 71460
rect 164016 71420 165568 71448
rect 166966 71420 192300 71448
rect 164016 71408 164022 71420
rect 153562 71380 153568 71392
rect 137986 71352 153568 71380
rect 153562 71340 153568 71352
rect 153620 71340 153626 71392
rect 161014 71340 161020 71392
rect 161072 71380 161078 71392
rect 166966 71380 166994 71420
rect 192294 71408 192300 71420
rect 192352 71408 192358 71460
rect 161072 71352 166994 71380
rect 161072 71340 161078 71352
rect 169478 71340 169484 71392
rect 169536 71380 169542 71392
rect 196434 71380 196440 71392
rect 169536 71352 196440 71380
rect 169536 71340 169542 71352
rect 196434 71340 196440 71352
rect 196492 71340 196498 71392
rect 108574 71272 108580 71324
rect 108632 71312 108638 71324
rect 121454 71312 121460 71324
rect 108632 71284 121460 71312
rect 108632 71272 108638 71284
rect 121454 71272 121460 71284
rect 121512 71272 121518 71324
rect 123110 71272 123116 71324
rect 123168 71312 123174 71324
rect 152550 71312 152556 71324
rect 123168 71284 152556 71312
rect 123168 71272 123174 71284
rect 152550 71272 152556 71284
rect 152608 71272 152614 71324
rect 161382 71272 161388 71324
rect 161440 71312 161446 71324
rect 187142 71312 187148 71324
rect 161440 71284 187148 71312
rect 161440 71272 161446 71284
rect 187142 71272 187148 71284
rect 187200 71272 187206 71324
rect 108850 71204 108856 71256
rect 108908 71244 108914 71256
rect 138382 71244 138388 71256
rect 108908 71216 138388 71244
rect 108908 71204 108914 71216
rect 138382 71204 138388 71216
rect 138440 71244 138446 71256
rect 139026 71244 139032 71256
rect 138440 71216 139032 71244
rect 138440 71204 138446 71216
rect 139026 71204 139032 71216
rect 139084 71204 139090 71256
rect 162394 71204 162400 71256
rect 162452 71244 162458 71256
rect 188338 71244 188344 71256
rect 162452 71216 188344 71244
rect 162452 71204 162458 71216
rect 188338 71204 188344 71216
rect 188396 71204 188402 71256
rect 113358 71136 113364 71188
rect 113416 71176 113422 71188
rect 142338 71176 142344 71188
rect 113416 71148 142344 71176
rect 113416 71136 113422 71148
rect 142338 71136 142344 71148
rect 142396 71136 142402 71188
rect 153562 71136 153568 71188
rect 153620 71176 153626 71188
rect 153930 71176 153936 71188
rect 153620 71148 153936 71176
rect 153620 71136 153626 71148
rect 153930 71136 153936 71148
rect 153988 71136 153994 71188
rect 165430 71136 165436 71188
rect 165488 71176 165494 71188
rect 186958 71176 186964 71188
rect 165488 71148 186964 71176
rect 165488 71136 165494 71148
rect 186958 71136 186964 71148
rect 187016 71136 187022 71188
rect 115290 71068 115296 71120
rect 115348 71108 115354 71120
rect 138566 71108 138572 71120
rect 115348 71080 138572 71108
rect 115348 71068 115354 71080
rect 138566 71068 138572 71080
rect 138624 71068 138630 71120
rect 148870 71068 148876 71120
rect 148928 71108 148934 71120
rect 148928 71080 157334 71108
rect 148928 71068 148934 71080
rect 27614 71000 27620 71052
rect 27672 71040 27678 71052
rect 100110 71040 100116 71052
rect 27672 71012 100116 71040
rect 27672 71000 27678 71012
rect 100110 71000 100116 71012
rect 100168 71000 100174 71052
rect 102778 71000 102784 71052
rect 102836 71040 102842 71052
rect 106826 71040 106832 71052
rect 102836 71012 106832 71040
rect 102836 71000 102842 71012
rect 106826 71000 106832 71012
rect 106884 71000 106890 71052
rect 116118 71000 116124 71052
rect 116176 71040 116182 71052
rect 136910 71040 136916 71052
rect 116176 71012 136916 71040
rect 116176 71000 116182 71012
rect 136910 71000 136916 71012
rect 136968 71040 136974 71052
rect 142798 71040 142804 71052
rect 136968 71012 142804 71040
rect 136968 71000 136974 71012
rect 142798 71000 142804 71012
rect 142856 71000 142862 71052
rect 153562 71000 153568 71052
rect 153620 71040 153626 71052
rect 154114 71040 154120 71052
rect 153620 71012 154120 71040
rect 153620 71000 153626 71012
rect 154114 71000 154120 71012
rect 154172 71000 154178 71052
rect 157306 71040 157334 71080
rect 184198 71040 184204 71052
rect 157306 71012 184204 71040
rect 184198 71000 184204 71012
rect 184256 71000 184262 71052
rect 192110 71000 192116 71052
rect 192168 71040 192174 71052
rect 192846 71040 192852 71052
rect 192168 71012 192852 71040
rect 192168 71000 192174 71012
rect 192846 71000 192852 71012
rect 192904 71040 192910 71052
rect 200114 71040 200120 71052
rect 192904 71012 200120 71040
rect 192904 71000 192910 71012
rect 200114 71000 200120 71012
rect 200172 71000 200178 71052
rect 121454 70932 121460 70984
rect 121512 70972 121518 70984
rect 142062 70972 142068 70984
rect 121512 70944 142068 70972
rect 121512 70932 121518 70944
rect 142062 70932 142068 70944
rect 142120 70932 142126 70984
rect 142430 70864 142436 70916
rect 142488 70904 142494 70916
rect 142798 70904 142804 70916
rect 142488 70876 142804 70904
rect 142488 70864 142494 70876
rect 142798 70864 142804 70876
rect 142856 70864 142862 70916
rect 150802 70864 150808 70916
rect 150860 70904 150866 70916
rect 151262 70904 151268 70916
rect 150860 70876 151268 70904
rect 150860 70864 150866 70876
rect 151262 70864 151268 70876
rect 151320 70864 151326 70916
rect 166350 70864 166356 70916
rect 166408 70904 166414 70916
rect 200022 70904 200028 70916
rect 166408 70876 200028 70904
rect 166408 70864 166414 70876
rect 200022 70864 200028 70876
rect 200080 70864 200086 70916
rect 187602 70456 187608 70508
rect 187660 70496 187666 70508
rect 480254 70496 480260 70508
rect 187660 70468 480260 70496
rect 187660 70456 187666 70468
rect 480254 70456 480260 70468
rect 480312 70456 480318 70508
rect 190362 70388 190368 70440
rect 190420 70428 190426 70440
rect 531314 70428 531320 70440
rect 190420 70400 531320 70428
rect 190420 70388 190426 70400
rect 531314 70388 531320 70400
rect 531372 70388 531378 70440
rect 116762 70320 116768 70372
rect 116820 70360 116826 70372
rect 151078 70360 151084 70372
rect 116820 70332 151084 70360
rect 116820 70320 116826 70332
rect 151078 70320 151084 70332
rect 151136 70320 151142 70372
rect 168098 70320 168104 70372
rect 168156 70360 168162 70372
rect 202230 70360 202236 70372
rect 168156 70332 202236 70360
rect 168156 70320 168162 70332
rect 202230 70320 202236 70332
rect 202288 70320 202294 70372
rect 120994 70252 121000 70304
rect 121052 70292 121058 70304
rect 154666 70292 154672 70304
rect 121052 70264 154672 70292
rect 121052 70252 121058 70264
rect 154666 70252 154672 70264
rect 154724 70292 154730 70304
rect 155402 70292 155408 70304
rect 154724 70264 155408 70292
rect 154724 70252 154730 70264
rect 155402 70252 155408 70264
rect 155460 70252 155466 70304
rect 166534 70252 166540 70304
rect 166592 70292 166598 70304
rect 166718 70292 166724 70304
rect 166592 70264 166724 70292
rect 166592 70252 166598 70264
rect 166718 70252 166724 70264
rect 166776 70252 166782 70304
rect 169570 70252 169576 70304
rect 169628 70292 169634 70304
rect 203518 70292 203524 70304
rect 169628 70264 203524 70292
rect 169628 70252 169634 70264
rect 203518 70252 203524 70264
rect 203576 70252 203582 70304
rect 117498 70184 117504 70236
rect 117556 70224 117562 70236
rect 152274 70224 152280 70236
rect 117556 70196 152280 70224
rect 117556 70184 117562 70196
rect 152274 70184 152280 70196
rect 152332 70224 152338 70236
rect 152550 70224 152556 70236
rect 152332 70196 152556 70224
rect 152332 70184 152338 70196
rect 152550 70184 152556 70196
rect 152608 70184 152614 70236
rect 168282 70184 168288 70236
rect 168340 70224 168346 70236
rect 198274 70224 198280 70236
rect 168340 70196 198280 70224
rect 168340 70184 168346 70196
rect 198274 70184 198280 70196
rect 198332 70184 198338 70236
rect 105998 70116 106004 70168
rect 106056 70156 106062 70168
rect 140222 70156 140228 70168
rect 106056 70128 140228 70156
rect 106056 70116 106062 70128
rect 140222 70116 140228 70128
rect 140280 70116 140286 70168
rect 165890 70116 165896 70168
rect 165948 70156 165954 70168
rect 166718 70156 166724 70168
rect 165948 70128 166724 70156
rect 165948 70116 165954 70128
rect 166718 70116 166724 70128
rect 166776 70156 166782 70168
rect 194134 70156 194140 70168
rect 166776 70128 194140 70156
rect 166776 70116 166782 70128
rect 194134 70116 194140 70128
rect 194192 70116 194198 70168
rect 122190 70048 122196 70100
rect 122248 70088 122254 70100
rect 154942 70088 154948 70100
rect 122248 70060 154948 70088
rect 122248 70048 122254 70060
rect 154942 70048 154948 70060
rect 155000 70088 155006 70100
rect 155310 70088 155316 70100
rect 155000 70060 155316 70088
rect 155000 70048 155006 70060
rect 155310 70048 155316 70060
rect 155368 70048 155374 70100
rect 166902 70048 166908 70100
rect 166960 70088 166966 70100
rect 192570 70088 192576 70100
rect 166960 70060 192576 70088
rect 166960 70048 166966 70060
rect 192570 70048 192576 70060
rect 192628 70048 192634 70100
rect 102134 69980 102140 70032
rect 102192 70020 102198 70032
rect 102962 70020 102968 70032
rect 102192 69992 102968 70020
rect 102192 69980 102198 69992
rect 102962 69980 102968 69992
rect 103020 70020 103026 70032
rect 136542 70020 136548 70032
rect 103020 69992 136548 70020
rect 103020 69980 103026 69992
rect 136542 69980 136548 69992
rect 136600 69980 136606 70032
rect 171962 69980 171968 70032
rect 172020 70020 172026 70032
rect 192754 70020 192760 70032
rect 172020 69992 192760 70020
rect 172020 69980 172026 69992
rect 192754 69980 192760 69992
rect 192812 69980 192818 70032
rect 103514 69912 103520 69964
rect 103572 69952 103578 69964
rect 105998 69952 106004 69964
rect 103572 69924 106004 69952
rect 103572 69912 103578 69924
rect 105998 69912 106004 69924
rect 106056 69912 106062 69964
rect 110230 69912 110236 69964
rect 110288 69952 110294 69964
rect 142614 69952 142620 69964
rect 110288 69924 142620 69952
rect 110288 69912 110294 69924
rect 142614 69912 142620 69924
rect 142672 69912 142678 69964
rect 175826 69912 175832 69964
rect 175884 69952 175890 69964
rect 199562 69952 199568 69964
rect 175884 69924 199568 69952
rect 175884 69912 175890 69924
rect 199562 69912 199568 69924
rect 199620 69912 199626 69964
rect 89714 69844 89720 69896
rect 89772 69884 89778 69896
rect 107010 69884 107016 69896
rect 89772 69856 107016 69884
rect 89772 69844 89778 69856
rect 107010 69844 107016 69856
rect 107068 69844 107074 69896
rect 110322 69844 110328 69896
rect 110380 69884 110386 69896
rect 142430 69884 142436 69896
rect 110380 69856 142436 69884
rect 110380 69844 110386 69856
rect 142430 69844 142436 69856
rect 142488 69884 142494 69896
rect 142706 69884 142712 69896
rect 142488 69856 142712 69884
rect 142488 69844 142494 69856
rect 142706 69844 142712 69856
rect 142764 69844 142770 69896
rect 147030 69844 147036 69896
rect 147088 69884 147094 69896
rect 179414 69884 179420 69896
rect 147088 69856 179420 69884
rect 147088 69844 147094 69856
rect 179414 69844 179420 69856
rect 179472 69844 179478 69896
rect 46198 69776 46204 69828
rect 46256 69816 46262 69828
rect 103330 69816 103336 69828
rect 46256 69788 103336 69816
rect 46256 69776 46262 69788
rect 103330 69776 103336 69788
rect 103388 69816 103394 69828
rect 134702 69816 134708 69828
rect 103388 69788 134708 69816
rect 103388 69776 103394 69788
rect 134702 69776 134708 69788
rect 134760 69776 134766 69828
rect 147858 69776 147864 69828
rect 147916 69816 147922 69828
rect 196618 69816 196624 69828
rect 147916 69788 196624 69816
rect 147916 69776 147922 69788
rect 196618 69776 196624 69788
rect 196676 69776 196682 69828
rect 41414 69708 41420 69760
rect 41472 69748 41478 69760
rect 102134 69748 102140 69760
rect 41472 69720 102140 69748
rect 41472 69708 41478 69720
rect 102134 69708 102140 69720
rect 102192 69708 102198 69760
rect 122558 69708 122564 69760
rect 122616 69748 122622 69760
rect 153286 69748 153292 69760
rect 122616 69720 153292 69748
rect 122616 69708 122622 69720
rect 153286 69708 153292 69720
rect 153344 69748 153350 69760
rect 153838 69748 153844 69760
rect 153344 69720 153844 69748
rect 153344 69708 153350 69720
rect 153838 69708 153844 69720
rect 153896 69708 153902 69760
rect 160186 69708 160192 69760
rect 160244 69748 160250 69760
rect 354674 69748 354680 69760
rect 160244 69720 354680 69748
rect 160244 69708 160250 69720
rect 354674 69708 354680 69720
rect 354732 69708 354738 69760
rect 18598 69640 18604 69692
rect 18656 69680 18662 69692
rect 103422 69680 103428 69692
rect 18656 69652 103428 69680
rect 18656 69640 18662 69652
rect 103422 69640 103428 69652
rect 103480 69680 103486 69692
rect 103480 69640 103514 69680
rect 113542 69640 113548 69692
rect 113600 69680 113606 69692
rect 142154 69680 142160 69692
rect 113600 69652 142160 69680
rect 113600 69640 113606 69652
rect 142154 69640 142160 69652
rect 142212 69680 142218 69692
rect 142982 69680 142988 69692
rect 142212 69652 142988 69680
rect 142212 69640 142218 69652
rect 142982 69640 142988 69652
rect 143040 69640 143046 69692
rect 143718 69640 143724 69692
rect 143776 69680 143782 69692
rect 147030 69680 147036 69692
rect 143776 69652 147036 69680
rect 143776 69640 143782 69652
rect 147030 69640 147036 69652
rect 147088 69640 147094 69692
rect 147214 69640 147220 69692
rect 147272 69680 147278 69692
rect 182818 69680 182824 69692
rect 147272 69652 182824 69680
rect 147272 69640 147278 69652
rect 182818 69640 182824 69652
rect 182876 69640 182882 69692
rect 192754 69640 192760 69692
rect 192812 69680 192818 69692
rect 430574 69680 430580 69692
rect 192812 69652 430580 69680
rect 192812 69640 192818 69652
rect 430574 69640 430580 69652
rect 430632 69640 430638 69692
rect 103486 69544 103514 69640
rect 116302 69572 116308 69624
rect 116360 69612 116366 69624
rect 128446 69612 128452 69624
rect 116360 69584 128452 69612
rect 116360 69572 116366 69584
rect 128446 69572 128452 69584
rect 128504 69612 128510 69624
rect 141602 69612 141608 69624
rect 128504 69584 141608 69612
rect 128504 69572 128510 69584
rect 141602 69572 141608 69584
rect 141660 69572 141666 69624
rect 166534 69572 166540 69624
rect 166592 69612 166598 69624
rect 188430 69612 188436 69624
rect 166592 69584 188436 69612
rect 166592 69572 166598 69584
rect 188430 69572 188436 69584
rect 188488 69572 188494 69624
rect 133690 69544 133696 69556
rect 103486 69516 133696 69544
rect 133690 69504 133696 69516
rect 133748 69504 133754 69556
rect 199562 69028 199568 69080
rect 199620 69068 199626 69080
rect 561674 69068 561680 69080
rect 199620 69040 561680 69068
rect 199620 69028 199626 69040
rect 561674 69028 561680 69040
rect 561732 69028 561738 69080
rect 109034 68960 109040 69012
rect 109092 69000 109098 69012
rect 110966 69000 110972 69012
rect 109092 68972 110972 69000
rect 109092 68960 109098 68972
rect 110966 68960 110972 68972
rect 111024 68960 111030 69012
rect 135438 69000 135444 69012
rect 113146 68972 135444 69000
rect 104526 68892 104532 68944
rect 104584 68932 104590 68944
rect 104802 68932 104808 68944
rect 104584 68904 104808 68932
rect 104584 68892 104590 68904
rect 104802 68892 104808 68904
rect 104860 68932 104866 68944
rect 113146 68932 113174 68972
rect 135438 68960 135444 68972
rect 135496 68960 135502 69012
rect 145374 68960 145380 69012
rect 145432 69000 145438 69012
rect 147122 69000 147128 69012
rect 145432 68972 147128 69000
rect 145432 68960 145438 68972
rect 147122 68960 147128 68972
rect 147180 68960 147186 69012
rect 164326 68960 164332 69012
rect 164384 69000 164390 69012
rect 199102 69000 199108 69012
rect 164384 68972 199108 69000
rect 164384 68960 164390 68972
rect 199102 68960 199108 68972
rect 199160 69000 199166 69012
rect 199654 69000 199660 69012
rect 199160 68972 199660 69000
rect 199160 68960 199166 68972
rect 199654 68960 199660 68972
rect 199712 68960 199718 69012
rect 104860 68904 113174 68932
rect 104860 68892 104866 68904
rect 161474 68892 161480 68944
rect 161532 68932 161538 68944
rect 195238 68932 195244 68944
rect 161532 68904 195244 68932
rect 161532 68892 161538 68904
rect 195238 68892 195244 68904
rect 195296 68892 195302 68944
rect 180334 68824 180340 68876
rect 180392 68864 180398 68876
rect 182174 68864 182180 68876
rect 180392 68836 182180 68864
rect 180392 68824 180398 68836
rect 182174 68824 182180 68836
rect 182232 68824 182238 68876
rect 196250 68864 196256 68876
rect 190426 68836 196256 68864
rect 176746 68756 176752 68808
rect 176804 68796 176810 68808
rect 190426 68796 190454 68836
rect 196250 68824 196256 68836
rect 196308 68824 196314 68876
rect 176804 68768 190454 68796
rect 176804 68756 176810 68768
rect 195238 68416 195244 68468
rect 195296 68456 195302 68468
rect 367094 68456 367100 68468
rect 195296 68428 367100 68456
rect 195296 68416 195302 68428
rect 367094 68416 367100 68428
rect 367152 68416 367158 68468
rect 199102 68348 199108 68400
rect 199160 68388 199166 68400
rect 412634 68388 412640 68400
rect 199160 68360 412640 68388
rect 199160 68348 199166 68360
rect 412634 68348 412640 68360
rect 412692 68348 412698 68400
rect 48314 68280 48320 68332
rect 48372 68320 48378 68332
rect 104802 68320 104808 68332
rect 48372 68292 104808 68320
rect 48372 68280 48378 68292
rect 104802 68280 104808 68292
rect 104860 68280 104866 68332
rect 167730 68280 167736 68332
rect 167788 68320 167794 68332
rect 453298 68320 453304 68332
rect 167788 68292 453304 68320
rect 167788 68280 167794 68292
rect 453298 68280 453304 68292
rect 453356 68280 453362 68332
rect 196250 67600 196256 67652
rect 196308 67640 196314 67652
rect 574738 67640 574744 67652
rect 196308 67612 574744 67640
rect 196308 67600 196314 67612
rect 574738 67600 574744 67612
rect 574796 67600 574802 67652
rect 110046 67532 110052 67584
rect 110104 67572 110110 67584
rect 143994 67572 144000 67584
rect 110104 67544 144000 67572
rect 110104 67532 110110 67544
rect 143994 67532 144000 67544
rect 144052 67532 144058 67584
rect 155126 67532 155132 67584
rect 155184 67572 155190 67584
rect 189258 67572 189264 67584
rect 155184 67544 189264 67572
rect 155184 67532 155190 67544
rect 189258 67532 189264 67544
rect 189316 67532 189322 67584
rect 108942 67464 108948 67516
rect 109000 67504 109006 67516
rect 135438 67504 135444 67516
rect 109000 67476 135444 67504
rect 109000 67464 109006 67476
rect 135438 67464 135444 67476
rect 135496 67504 135502 67516
rect 135806 67504 135812 67516
rect 135496 67476 135812 67504
rect 135496 67464 135502 67476
rect 135806 67464 135812 67476
rect 135864 67464 135870 67516
rect 163038 67464 163044 67516
rect 163096 67504 163102 67516
rect 195146 67504 195152 67516
rect 163096 67476 195152 67504
rect 163096 67464 163102 67476
rect 195146 67464 195152 67476
rect 195204 67464 195210 67516
rect 175642 67396 175648 67448
rect 175700 67436 175706 67448
rect 200850 67436 200856 67448
rect 175700 67408 200856 67436
rect 175700 67396 175706 67408
rect 200850 67396 200856 67408
rect 200908 67436 200914 67448
rect 201402 67436 201408 67448
rect 200908 67408 201408 67436
rect 200908 67396 200914 67408
rect 201402 67396 201408 67408
rect 201460 67396 201466 67448
rect 78674 67056 78680 67108
rect 78732 67096 78738 67108
rect 108482 67096 108488 67108
rect 78732 67068 108488 67096
rect 78732 67056 78738 67068
rect 108482 67056 108488 67068
rect 108540 67056 108546 67108
rect 120074 67056 120080 67108
rect 120132 67096 120138 67108
rect 141970 67096 141976 67108
rect 120132 67068 141976 67096
rect 120132 67056 120138 67068
rect 141970 67056 141976 67068
rect 142028 67056 142034 67108
rect 75914 66988 75920 67040
rect 75972 67028 75978 67040
rect 107102 67028 107108 67040
rect 75972 67000 107108 67028
rect 75972 66988 75978 67000
rect 107102 66988 107108 67000
rect 107160 66988 107166 67040
rect 113174 66988 113180 67040
rect 113232 67028 113238 67040
rect 141050 67028 141056 67040
rect 113232 67000 141056 67028
rect 113232 66988 113238 67000
rect 141050 66988 141056 67000
rect 141108 66988 141114 67040
rect 150618 66988 150624 67040
rect 150676 67028 150682 67040
rect 242894 67028 242900 67040
rect 150676 67000 242900 67028
rect 150676 66988 150682 67000
rect 242894 66988 242900 67000
rect 242952 66988 242958 67040
rect 80054 66920 80060 66972
rect 80112 66960 80118 66972
rect 113450 66960 113456 66972
rect 80112 66932 113456 66960
rect 80112 66920 80118 66932
rect 113450 66920 113456 66932
rect 113508 66920 113514 66972
rect 117314 66920 117320 66972
rect 117372 66960 117378 66972
rect 140958 66960 140964 66972
rect 117372 66932 140964 66960
rect 117372 66920 117378 66932
rect 140958 66920 140964 66932
rect 141016 66920 141022 66972
rect 189258 66920 189264 66972
rect 189316 66960 189322 66972
rect 295334 66960 295340 66972
rect 189316 66932 295340 66960
rect 189316 66920 189322 66932
rect 295334 66920 295340 66932
rect 295392 66920 295398 66972
rect 60734 66852 60740 66904
rect 60792 66892 60798 66904
rect 137278 66892 137284 66904
rect 60792 66864 137284 66892
rect 60792 66852 60798 66864
rect 137278 66852 137284 66864
rect 137336 66852 137342 66904
rect 195146 66852 195152 66904
rect 195204 66892 195210 66904
rect 402974 66892 402980 66904
rect 195204 66864 402980 66892
rect 195204 66852 195210 66864
rect 402974 66852 402980 66864
rect 403032 66852 403038 66904
rect 140774 66240 140780 66292
rect 140832 66280 140838 66292
rect 142154 66280 142160 66292
rect 140832 66252 142160 66280
rect 140832 66240 140838 66252
rect 142154 66240 142160 66252
rect 142212 66240 142218 66292
rect 201402 66240 201408 66292
rect 201460 66280 201466 66292
rect 557534 66280 557540 66292
rect 201460 66252 557540 66280
rect 201460 66240 201466 66252
rect 557534 66240 557540 66252
rect 557592 66240 557598 66292
rect 102134 66172 102140 66224
rect 102192 66212 102198 66224
rect 103238 66212 103244 66224
rect 102192 66184 103244 66212
rect 102192 66172 102198 66184
rect 103238 66172 103244 66184
rect 103296 66212 103302 66224
rect 137186 66212 137192 66224
rect 103296 66184 137192 66212
rect 103296 66172 103302 66184
rect 137186 66172 137192 66184
rect 137244 66172 137250 66224
rect 144362 66172 144368 66224
rect 144420 66212 144426 66224
rect 147214 66212 147220 66224
rect 144420 66184 147220 66212
rect 144420 66172 144426 66184
rect 147214 66172 147220 66184
rect 147272 66172 147278 66224
rect 159174 66172 159180 66224
rect 159232 66212 159238 66224
rect 192018 66212 192024 66224
rect 159232 66184 192024 66212
rect 159232 66172 159238 66184
rect 192018 66172 192024 66184
rect 192076 66212 192082 66224
rect 193122 66212 193128 66224
rect 192076 66184 193128 66212
rect 192076 66172 192082 66184
rect 193122 66172 193128 66184
rect 193180 66172 193186 66224
rect 109126 66104 109132 66156
rect 109184 66144 109190 66156
rect 109954 66144 109960 66156
rect 109184 66116 109960 66144
rect 109184 66104 109190 66116
rect 109954 66104 109960 66116
rect 110012 66144 110018 66156
rect 139946 66144 139952 66156
rect 110012 66116 139952 66144
rect 110012 66104 110018 66116
rect 139946 66104 139952 66116
rect 140004 66104 140010 66156
rect 173158 66104 173164 66156
rect 173216 66144 173222 66156
rect 194042 66144 194048 66156
rect 173216 66116 194048 66144
rect 173216 66104 173222 66116
rect 194042 66104 194048 66116
rect 194100 66144 194106 66156
rect 194502 66144 194508 66156
rect 194100 66116 194508 66144
rect 194100 66104 194106 66116
rect 194502 66104 194508 66116
rect 194560 66104 194566 66156
rect 104802 66036 104808 66088
rect 104860 66076 104866 66088
rect 134334 66076 134340 66088
rect 104860 66048 134340 66076
rect 104860 66036 104866 66048
rect 134334 66036 134340 66048
rect 134392 66036 134398 66088
rect 116578 66008 116584 66020
rect 113146 65980 116584 66008
rect 97994 65696 98000 65748
rect 98052 65736 98058 65748
rect 109126 65736 109132 65748
rect 98052 65708 109132 65736
rect 98052 65696 98058 65708
rect 109126 65696 109132 65708
rect 109184 65696 109190 65748
rect 93118 65628 93124 65680
rect 93176 65668 93182 65680
rect 113146 65668 113174 65980
rect 116578 65968 116584 65980
rect 116636 66008 116642 66020
rect 139854 66008 139860 66020
rect 116636 65980 139860 66008
rect 116636 65968 116642 65980
rect 139854 65968 139860 65980
rect 139912 65968 139918 66020
rect 93176 65640 113174 65668
rect 93176 65628 93182 65640
rect 148410 65628 148416 65680
rect 148468 65668 148474 65680
rect 207014 65668 207020 65680
rect 148468 65640 207020 65668
rect 148468 65628 148474 65640
rect 207014 65628 207020 65640
rect 207072 65628 207078 65680
rect 57238 65560 57244 65612
rect 57296 65600 57302 65612
rect 102134 65600 102140 65612
rect 57296 65572 102140 65600
rect 57296 65560 57302 65572
rect 102134 65560 102140 65572
rect 102192 65560 102198 65612
rect 153746 65560 153752 65612
rect 153804 65600 153810 65612
rect 274634 65600 274640 65612
rect 153804 65572 274640 65600
rect 153804 65560 153810 65572
rect 274634 65560 274640 65572
rect 274692 65560 274698 65612
rect 35986 65492 35992 65544
rect 36044 65532 36050 65544
rect 104802 65532 104808 65544
rect 36044 65504 104808 65532
rect 36044 65492 36050 65504
rect 104802 65492 104808 65504
rect 104860 65492 104866 65544
rect 146386 65492 146392 65544
rect 146444 65532 146450 65544
rect 183554 65532 183560 65544
rect 146444 65504 183560 65532
rect 146444 65492 146450 65504
rect 183554 65492 183560 65504
rect 183612 65492 183618 65544
rect 193122 65492 193128 65544
rect 193180 65532 193186 65544
rect 346394 65532 346400 65544
rect 193180 65504 346400 65532
rect 193180 65492 193186 65504
rect 346394 65492 346400 65504
rect 346452 65492 346458 65544
rect 142246 64988 142252 65000
rect 142172 64960 142252 64988
rect 139394 64880 139400 64932
rect 139452 64920 139458 64932
rect 142172 64920 142200 64960
rect 142246 64948 142252 64960
rect 142304 64948 142310 65000
rect 139452 64892 142200 64920
rect 139452 64880 139458 64892
rect 194502 64880 194508 64932
rect 194560 64920 194566 64932
rect 529934 64920 529940 64932
rect 194560 64892 529940 64920
rect 194560 64880 194566 64892
rect 529934 64880 529940 64892
rect 529992 64880 529998 64932
rect 106182 64812 106188 64864
rect 106240 64852 106246 64864
rect 137094 64852 137100 64864
rect 106240 64824 137100 64852
rect 106240 64812 106246 64824
rect 137094 64812 137100 64824
rect 137152 64812 137158 64864
rect 160186 64812 160192 64864
rect 160244 64852 160250 64864
rect 194870 64852 194876 64864
rect 160244 64824 194876 64852
rect 160244 64812 160250 64824
rect 194870 64812 194876 64824
rect 194928 64812 194934 64864
rect 168650 64744 168656 64796
rect 168708 64784 168714 64796
rect 203242 64784 203248 64796
rect 168708 64756 203248 64784
rect 168708 64744 168714 64756
rect 203242 64744 203248 64756
rect 203300 64744 203306 64796
rect 149882 64268 149888 64320
rect 149940 64308 149946 64320
rect 224954 64308 224960 64320
rect 149940 64280 224960 64308
rect 149940 64268 149946 64280
rect 224954 64268 224960 64280
rect 225012 64268 225018 64320
rect 62114 64200 62120 64252
rect 62172 64240 62178 64252
rect 106182 64240 106188 64252
rect 62172 64212 106188 64240
rect 62172 64200 62178 64212
rect 106182 64200 106188 64212
rect 106240 64200 106246 64252
rect 194870 64200 194876 64252
rect 194928 64240 194934 64252
rect 358814 64240 358820 64252
rect 194928 64212 358820 64240
rect 194928 64200 194934 64212
rect 358814 64200 358820 64212
rect 358872 64200 358878 64252
rect 4154 64132 4160 64184
rect 4212 64172 4218 64184
rect 133414 64172 133420 64184
rect 4212 64144 133420 64172
rect 4212 64132 4218 64144
rect 133414 64132 133420 64144
rect 133472 64132 133478 64184
rect 147398 64132 147404 64184
rect 147456 64172 147462 64184
rect 187694 64172 187700 64184
rect 147456 64144 187700 64172
rect 147456 64132 147462 64144
rect 187694 64132 187700 64144
rect 187752 64132 187758 64184
rect 203242 64132 203248 64184
rect 203300 64172 203306 64184
rect 472618 64172 472624 64184
rect 203300 64144 472624 64172
rect 203300 64132 203306 64144
rect 472618 64132 472624 64144
rect 472676 64132 472682 64184
rect 104618 63452 104624 63504
rect 104676 63492 104682 63504
rect 132770 63492 132776 63504
rect 104676 63464 132776 63492
rect 104676 63452 104682 63464
rect 132770 63452 132776 63464
rect 132828 63452 132834 63504
rect 159082 63452 159088 63504
rect 159140 63492 159146 63504
rect 193490 63492 193496 63504
rect 159140 63464 193496 63492
rect 159140 63452 159146 63464
rect 193490 63452 193496 63464
rect 193548 63452 193554 63504
rect 75178 62908 75184 62960
rect 75236 62948 75242 62960
rect 104158 62948 104164 62960
rect 75236 62920 104164 62948
rect 75236 62908 75242 62920
rect 104158 62908 104164 62920
rect 104216 62908 104222 62960
rect 88334 62840 88340 62892
rect 88392 62880 88398 62892
rect 139210 62880 139216 62892
rect 88392 62852 139216 62880
rect 88392 62840 88398 62852
rect 139210 62840 139216 62852
rect 139268 62840 139274 62892
rect 178862 62840 178868 62892
rect 178920 62880 178926 62892
rect 227714 62880 227720 62892
rect 178920 62852 227720 62880
rect 178920 62840 178926 62852
rect 227714 62840 227720 62852
rect 227772 62840 227778 62892
rect 10318 62772 10324 62824
rect 10376 62812 10382 62824
rect 104618 62812 104624 62824
rect 10376 62784 104624 62812
rect 10376 62772 10382 62784
rect 104618 62772 104624 62784
rect 104676 62772 104682 62824
rect 193490 62772 193496 62824
rect 193548 62812 193554 62824
rect 340874 62812 340880 62824
rect 193548 62784 340880 62812
rect 193548 62772 193554 62784
rect 340874 62772 340880 62784
rect 340932 62772 340938 62824
rect 197446 62160 197452 62212
rect 197504 62200 197510 62212
rect 197722 62200 197728 62212
rect 197504 62172 197728 62200
rect 197504 62160 197510 62172
rect 197722 62160 197728 62172
rect 197780 62160 197786 62212
rect 104526 62024 104532 62076
rect 104584 62064 104590 62076
rect 104710 62064 104716 62076
rect 104584 62036 104716 62064
rect 104584 62024 104590 62036
rect 104710 62024 104716 62036
rect 104768 62064 104774 62076
rect 135990 62064 135996 62076
rect 104768 62036 135996 62064
rect 104768 62024 104774 62036
rect 135990 62024 135996 62036
rect 136048 62024 136054 62076
rect 162946 62024 162952 62076
rect 163004 62064 163010 62076
rect 197446 62064 197452 62076
rect 163004 62036 197452 62064
rect 163004 62024 163010 62036
rect 197446 62024 197452 62036
rect 197504 62064 197510 62076
rect 197630 62064 197636 62076
rect 197504 62036 197636 62064
rect 197504 62024 197510 62036
rect 197630 62024 197636 62036
rect 197688 62024 197694 62076
rect 167178 61956 167184 62008
rect 167236 61996 167242 62008
rect 199010 61996 199016 62008
rect 167236 61968 199016 61996
rect 167236 61956 167242 61968
rect 199010 61956 199016 61968
rect 199068 61956 199074 62008
rect 52546 61412 52552 61464
rect 52604 61452 52610 61464
rect 104526 61452 104532 61464
rect 52604 61424 104532 61452
rect 52604 61412 52610 61424
rect 104526 61412 104532 61424
rect 104584 61412 104590 61464
rect 197446 61412 197452 61464
rect 197504 61452 197510 61464
rect 394694 61452 394700 61464
rect 197504 61424 394700 61452
rect 197504 61412 197510 61424
rect 394694 61412 394700 61424
rect 394752 61412 394758 61464
rect 42794 61344 42800 61396
rect 42852 61384 42858 61396
rect 135714 61384 135720 61396
rect 42852 61356 135720 61384
rect 42852 61344 42858 61356
rect 135714 61344 135720 61356
rect 135772 61344 135778 61396
rect 199010 61344 199016 61396
rect 199068 61384 199074 61396
rect 459554 61384 459560 61396
rect 199068 61356 459560 61384
rect 199068 61344 199074 61356
rect 459554 61344 459560 61356
rect 459612 61344 459618 61396
rect 135254 61208 135260 61260
rect 135312 61248 135318 61260
rect 142522 61248 142528 61260
rect 135312 61220 142528 61248
rect 135312 61208 135318 61220
rect 142522 61208 142528 61220
rect 142580 61208 142586 61260
rect 99374 60664 99380 60716
rect 99432 60704 99438 60716
rect 100386 60704 100392 60716
rect 99432 60676 100392 60704
rect 99432 60664 99438 60676
rect 100386 60664 100392 60676
rect 100444 60704 100450 60716
rect 134426 60704 134432 60716
rect 100444 60676 134432 60704
rect 100444 60664 100450 60676
rect 134426 60664 134432 60676
rect 134484 60664 134490 60716
rect 162854 60664 162860 60716
rect 162912 60704 162918 60716
rect 197446 60704 197452 60716
rect 162912 60676 197452 60704
rect 162912 60664 162918 60676
rect 197446 60664 197452 60676
rect 197504 60704 197510 60716
rect 197722 60704 197728 60716
rect 197504 60676 197728 60704
rect 197504 60664 197510 60676
rect 197722 60664 197728 60676
rect 197780 60664 197786 60716
rect 99466 60596 99472 60648
rect 99524 60636 99530 60648
rect 100570 60636 100576 60648
rect 99524 60608 100576 60636
rect 99524 60596 99530 60608
rect 100570 60596 100576 60608
rect 100628 60636 100634 60648
rect 132678 60636 132684 60648
rect 100628 60608 132684 60636
rect 100628 60596 100634 60608
rect 132678 60596 132684 60608
rect 132736 60596 132742 60648
rect 166258 60596 166264 60648
rect 166316 60636 166322 60648
rect 194226 60636 194232 60648
rect 166316 60608 194232 60636
rect 166316 60596 166322 60608
rect 194226 60596 194232 60608
rect 194284 60636 194290 60648
rect 194502 60636 194508 60648
rect 194284 60608 194508 60636
rect 194284 60596 194290 60608
rect 194502 60596 194508 60608
rect 194560 60596 194566 60648
rect 107470 60528 107476 60580
rect 107528 60568 107534 60580
rect 137370 60568 137376 60580
rect 107528 60540 137376 60568
rect 107528 60528 107534 60540
rect 137370 60528 137376 60540
rect 137428 60528 137434 60580
rect 69014 60120 69020 60172
rect 69072 60160 69078 60172
rect 107470 60160 107476 60172
rect 69072 60132 107476 60160
rect 69072 60120 69078 60132
rect 107470 60120 107476 60132
rect 107528 60120 107534 60172
rect 23474 60052 23480 60104
rect 23532 60092 23538 60104
rect 99374 60092 99380 60104
rect 23532 60064 99380 60092
rect 23532 60052 23538 60064
rect 99374 60052 99380 60064
rect 99432 60052 99438 60104
rect 197446 60052 197452 60104
rect 197504 60092 197510 60104
rect 398834 60092 398840 60104
rect 197504 60064 398840 60092
rect 197504 60052 197510 60064
rect 398834 60052 398840 60064
rect 398892 60052 398898 60104
rect 17954 59984 17960 60036
rect 18012 60024 18018 60036
rect 99466 60024 99472 60036
rect 18012 59996 99472 60024
rect 18012 59984 18018 59996
rect 99466 59984 99472 59996
rect 99524 59984 99530 60036
rect 147306 59984 147312 60036
rect 147364 60024 147370 60036
rect 186314 60024 186320 60036
rect 147364 59996 186320 60024
rect 147364 59984 147370 59996
rect 186314 59984 186320 59996
rect 186372 59984 186378 60036
rect 194502 59984 194508 60036
rect 194560 60024 194566 60036
rect 396074 60024 396080 60036
rect 194560 59996 396080 60024
rect 194560 59984 194566 59996
rect 396074 59984 396080 59996
rect 396132 59984 396138 60036
rect 110506 59304 110512 59356
rect 110564 59344 110570 59356
rect 114922 59344 114928 59356
rect 110564 59316 114928 59344
rect 110564 59304 110570 59316
rect 114922 59304 114928 59316
rect 114980 59304 114986 59356
rect 144270 59304 144276 59356
rect 144328 59344 144334 59356
rect 148410 59344 148416 59356
rect 144328 59316 148416 59344
rect 144328 59304 144334 59316
rect 148410 59304 148416 59316
rect 148468 59304 148474 59356
rect 167086 59304 167092 59356
rect 167144 59344 167150 59356
rect 201954 59344 201960 59356
rect 167144 59316 201960 59344
rect 167144 59304 167150 59316
rect 201954 59304 201960 59316
rect 202012 59344 202018 59356
rect 202782 59344 202788 59356
rect 202012 59316 202788 59344
rect 202012 59304 202018 59316
rect 202782 59304 202788 59316
rect 202840 59304 202846 59356
rect 148962 58760 148968 58812
rect 149020 58800 149026 58812
rect 209866 58800 209872 58812
rect 149020 58772 209872 58800
rect 149020 58760 149026 58772
rect 209866 58760 209872 58772
rect 209924 58760 209930 58812
rect 202782 58692 202788 58744
rect 202840 58732 202846 58744
rect 448514 58732 448520 58744
rect 202840 58704 448520 58732
rect 202840 58692 202846 58704
rect 448514 58692 448520 58704
rect 448572 58692 448578 58744
rect 169938 58624 169944 58676
rect 169996 58664 170002 58676
rect 489914 58664 489920 58676
rect 169996 58636 489920 58664
rect 169996 58624 170002 58636
rect 489914 58624 489920 58636
rect 489972 58624 489978 58676
rect 168558 57876 168564 57928
rect 168616 57916 168622 57928
rect 203426 57916 203432 57928
rect 168616 57888 203432 57916
rect 168616 57876 168622 57888
rect 203426 57876 203432 57888
rect 203484 57916 203490 57928
rect 204162 57916 204168 57928
rect 203484 57888 204168 57916
rect 203484 57876 203490 57888
rect 204162 57876 204168 57888
rect 204220 57876 204226 57928
rect 158990 57808 158996 57860
rect 159048 57848 159054 57860
rect 193306 57848 193312 57860
rect 159048 57820 193312 57848
rect 159048 57808 159054 57820
rect 193306 57808 193312 57820
rect 193364 57848 193370 57860
rect 194502 57848 194508 57860
rect 193364 57820 194508 57848
rect 193364 57808 193370 57820
rect 194502 57808 194508 57820
rect 194560 57808 194566 57860
rect 151262 57332 151268 57384
rect 151320 57372 151326 57384
rect 235994 57372 236000 57384
rect 151320 57344 236000 57372
rect 151320 57332 151326 57344
rect 235994 57332 236000 57344
rect 236052 57332 236058 57384
rect 194502 57264 194508 57316
rect 194560 57304 194566 57316
rect 345014 57304 345020 57316
rect 194560 57276 345020 57304
rect 194560 57264 194566 57276
rect 345014 57264 345020 57276
rect 345072 57264 345078 57316
rect 77386 57196 77392 57248
rect 77444 57236 77450 57248
rect 112530 57236 112536 57248
rect 77444 57208 112536 57236
rect 77444 57196 77450 57208
rect 112530 57196 112536 57208
rect 112588 57196 112594 57248
rect 147766 57196 147772 57248
rect 147824 57236 147830 57248
rect 197446 57236 197452 57248
rect 147824 57208 197452 57236
rect 147824 57196 147830 57208
rect 197446 57196 197452 57208
rect 197504 57196 197510 57248
rect 204162 57196 204168 57248
rect 204220 57236 204226 57248
rect 473446 57236 473452 57248
rect 204220 57208 473452 57236
rect 204220 57196 204226 57208
rect 473446 57196 473452 57208
rect 473504 57196 473510 57248
rect 99374 56516 99380 56568
rect 99432 56556 99438 56568
rect 100662 56556 100668 56568
rect 99432 56528 100668 56556
rect 99432 56516 99438 56528
rect 100662 56516 100668 56528
rect 100720 56556 100726 56568
rect 133598 56556 133604 56568
rect 100720 56528 133604 56556
rect 100720 56516 100726 56528
rect 133598 56516 133604 56528
rect 133656 56516 133662 56568
rect 167822 56516 167828 56568
rect 167880 56556 167886 56568
rect 201862 56556 201868 56568
rect 167880 56528 201868 56556
rect 167880 56516 167886 56528
rect 201862 56516 201868 56528
rect 201920 56556 201926 56568
rect 202782 56556 202788 56568
rect 201920 56528 202788 56556
rect 201920 56516 201926 56528
rect 202782 56516 202788 56528
rect 202840 56516 202846 56568
rect 158898 56448 158904 56500
rect 158956 56488 158962 56500
rect 193398 56488 193404 56500
rect 158956 56460 193404 56488
rect 158956 56448 158962 56460
rect 193398 56448 193404 56460
rect 193456 56488 193462 56500
rect 194502 56488 194508 56500
rect 193456 56460 194508 56488
rect 193456 56448 193462 56460
rect 194502 56448 194508 56460
rect 194560 56448 194566 56500
rect 176930 56380 176936 56432
rect 176988 56420 176994 56432
rect 200666 56420 200672 56432
rect 176988 56392 200672 56420
rect 176988 56380 176994 56392
rect 200666 56380 200672 56392
rect 200724 56420 200730 56432
rect 201402 56420 201408 56432
rect 200724 56392 201408 56420
rect 200724 56380 200730 56392
rect 201402 56380 201408 56392
rect 201460 56380 201466 56432
rect 63494 55904 63500 55956
rect 63552 55944 63558 55956
rect 136818 55944 136824 55956
rect 63552 55916 136824 55944
rect 63552 55904 63558 55916
rect 136818 55904 136824 55916
rect 136876 55904 136882 55956
rect 194502 55904 194508 55956
rect 194560 55944 194566 55956
rect 349154 55944 349160 55956
rect 194560 55916 349160 55944
rect 194560 55904 194566 55916
rect 349154 55904 349160 55916
rect 349212 55904 349218 55956
rect 12434 55836 12440 55888
rect 12492 55876 12498 55888
rect 99374 55876 99380 55888
rect 12492 55848 99380 55876
rect 12492 55836 12498 55848
rect 99374 55836 99380 55848
rect 99432 55836 99438 55888
rect 145742 55836 145748 55888
rect 145800 55876 145806 55888
rect 162118 55876 162124 55888
rect 145800 55848 162124 55876
rect 145800 55836 145806 55848
rect 162118 55836 162124 55848
rect 162176 55836 162182 55888
rect 202782 55836 202788 55888
rect 202840 55876 202846 55888
rect 450538 55876 450544 55888
rect 202840 55848 450544 55876
rect 202840 55836 202846 55848
rect 450538 55836 450544 55848
rect 450596 55836 450602 55888
rect 138658 55224 138664 55276
rect 138716 55264 138722 55276
rect 142246 55264 142252 55276
rect 138716 55236 142252 55264
rect 138716 55224 138722 55236
rect 142246 55224 142252 55236
rect 142304 55224 142310 55276
rect 201402 55224 201408 55276
rect 201460 55264 201466 55276
rect 560938 55264 560944 55276
rect 201460 55236 560944 55264
rect 201460 55224 201466 55236
rect 560938 55224 560944 55236
rect 560996 55224 561002 55276
rect 169018 55156 169024 55208
rect 169076 55196 169082 55208
rect 203058 55196 203064 55208
rect 169076 55168 203064 55196
rect 169076 55156 169082 55168
rect 203058 55156 203064 55168
rect 203116 55156 203122 55208
rect 152826 54612 152832 54664
rect 152884 54652 152890 54664
rect 253934 54652 253940 54664
rect 152884 54624 253940 54652
rect 152884 54612 152890 54624
rect 253934 54612 253940 54624
rect 253992 54612 253998 54664
rect 84194 54544 84200 54596
rect 84252 54584 84258 54596
rect 115198 54584 115204 54596
rect 84252 54556 115204 54584
rect 84252 54544 84258 54556
rect 115198 54544 115204 54556
rect 115256 54544 115262 54596
rect 158070 54544 158076 54596
rect 158128 54584 158134 54596
rect 333974 54584 333980 54596
rect 158128 54556 333980 54584
rect 158128 54544 158134 54556
rect 333974 54544 333980 54556
rect 334032 54544 334038 54596
rect 99374 54476 99380 54528
rect 99432 54516 99438 54528
rect 139762 54516 139768 54528
rect 99432 54488 139768 54516
rect 99432 54476 99438 54488
rect 139762 54476 139768 54488
rect 139820 54476 139826 54528
rect 203058 54476 203064 54528
rect 203116 54516 203122 54528
rect 468478 54516 468484 54528
rect 203116 54488 468484 54516
rect 203116 54476 203122 54488
rect 468478 54476 468484 54488
rect 468536 54476 468542 54528
rect 100478 53728 100484 53780
rect 100536 53768 100542 53780
rect 133046 53768 133052 53780
rect 100536 53740 133052 53768
rect 100536 53728 100542 53740
rect 133046 53728 133052 53740
rect 133104 53728 133110 53780
rect 147674 53116 147680 53168
rect 147732 53156 147738 53168
rect 204254 53156 204260 53168
rect 147732 53128 204260 53156
rect 147732 53116 147738 53128
rect 204254 53116 204260 53128
rect 204312 53116 204318 53168
rect 9674 53048 9680 53100
rect 9732 53088 9738 53100
rect 100478 53088 100484 53100
rect 9732 53060 100484 53088
rect 9732 53048 9738 53060
rect 100478 53048 100484 53060
rect 100536 53048 100542 53100
rect 176102 53048 176108 53100
rect 176160 53088 176166 53100
rect 556154 53088 556160 53100
rect 176160 53060 556160 53088
rect 176160 53048 176166 53060
rect 556154 53048 556160 53060
rect 556212 53048 556218 53100
rect 143810 52844 143816 52896
rect 143868 52884 143874 52896
rect 148502 52884 148508 52896
rect 143868 52856 148508 52884
rect 143868 52844 143874 52856
rect 148502 52844 148508 52856
rect 148560 52844 148566 52896
rect 168374 52368 168380 52420
rect 168432 52408 168438 52420
rect 201494 52408 201500 52420
rect 168432 52380 201500 52408
rect 168432 52368 168438 52380
rect 201494 52368 201500 52380
rect 201552 52408 201558 52420
rect 202782 52408 202788 52420
rect 201552 52380 202788 52408
rect 201552 52368 201558 52380
rect 202782 52368 202788 52380
rect 202840 52368 202846 52420
rect 149790 51824 149796 51876
rect 149848 51864 149854 51876
rect 215294 51864 215300 51876
rect 149848 51836 215300 51864
rect 149848 51824 149854 51836
rect 215294 51824 215300 51836
rect 215352 51824 215358 51876
rect 202782 51756 202788 51808
rect 202840 51796 202846 51808
rect 464338 51796 464344 51808
rect 202840 51768 464344 51796
rect 202840 51756 202846 51768
rect 464338 51756 464344 51768
rect 464396 51756 464402 51808
rect 176654 51688 176660 51740
rect 176712 51728 176718 51740
rect 578234 51728 578240 51740
rect 176712 51700 578240 51728
rect 176712 51688 176718 51700
rect 578234 51688 578240 51700
rect 578292 51688 578298 51740
rect 100754 51008 100760 51060
rect 100812 51048 100818 51060
rect 101858 51048 101864 51060
rect 100812 51020 101864 51048
rect 100812 51008 100818 51020
rect 101858 51008 101864 51020
rect 101916 51048 101922 51060
rect 134242 51048 134248 51060
rect 101916 51020 134248 51048
rect 101916 51008 101922 51020
rect 134242 51008 134248 51020
rect 134300 51008 134306 51060
rect 93946 50396 93952 50448
rect 94004 50436 94010 50448
rect 105538 50436 105544 50448
rect 94004 50408 105544 50436
rect 94004 50396 94010 50408
rect 105538 50396 105544 50408
rect 105596 50396 105602 50448
rect 30374 50328 30380 50380
rect 30432 50368 30438 50380
rect 100754 50368 100760 50380
rect 30432 50340 100760 50368
rect 30432 50328 30438 50340
rect 100754 50328 100760 50340
rect 100812 50328 100818 50380
rect 155586 50328 155592 50380
rect 155644 50368 155650 50380
rect 293954 50368 293960 50380
rect 155644 50340 293960 50368
rect 155644 50328 155650 50340
rect 293954 50328 293960 50340
rect 294012 50328 294018 50380
rect 148778 49104 148784 49156
rect 148836 49144 148842 49156
rect 201494 49144 201500 49156
rect 148836 49116 201500 49144
rect 148836 49104 148842 49116
rect 201494 49104 201500 49116
rect 201552 49104 201558 49156
rect 149974 49036 149980 49088
rect 150032 49076 150038 49088
rect 218146 49076 218152 49088
rect 150032 49048 218152 49076
rect 150032 49036 150038 49048
rect 218146 49036 218152 49048
rect 218204 49036 218210 49088
rect 170674 48968 170680 49020
rect 170732 49008 170738 49020
rect 486418 49008 486424 49020
rect 170732 48980 486424 49008
rect 170732 48968 170738 48980
rect 486418 48968 486424 48980
rect 486476 48968 486482 49020
rect 149238 47676 149244 47728
rect 149296 47716 149302 47728
rect 222194 47716 222200 47728
rect 149296 47688 222200 47716
rect 149296 47676 149302 47688
rect 222194 47676 222200 47688
rect 222252 47676 222258 47728
rect 151906 47608 151912 47660
rect 151964 47648 151970 47660
rect 267734 47648 267740 47660
rect 151964 47620 267740 47648
rect 151964 47608 151970 47620
rect 267734 47608 267740 47620
rect 267792 47608 267798 47660
rect 144178 47540 144184 47592
rect 144236 47580 144242 47592
rect 149238 47580 149244 47592
rect 144236 47552 149244 47580
rect 144236 47540 144242 47552
rect 149238 47540 149244 47552
rect 149296 47540 149302 47592
rect 173894 47540 173900 47592
rect 173952 47580 173958 47592
rect 542354 47580 542360 47592
rect 173952 47552 542360 47580
rect 173952 47540 173958 47552
rect 542354 47540 542360 47552
rect 542412 47540 542418 47592
rect 155402 46316 155408 46368
rect 155460 46356 155466 46368
rect 285674 46356 285680 46368
rect 155460 46328 285680 46356
rect 155460 46316 155466 46328
rect 285674 46316 285680 46328
rect 285732 46316 285738 46368
rect 165062 46248 165068 46300
rect 165120 46288 165126 46300
rect 418154 46288 418160 46300
rect 165120 46260 418160 46288
rect 165120 46248 165126 46260
rect 418154 46248 418160 46260
rect 418212 46248 418218 46300
rect 145190 46180 145196 46232
rect 145248 46220 145254 46232
rect 168374 46220 168380 46232
rect 145248 46192 168380 46220
rect 145248 46180 145254 46192
rect 168374 46180 168380 46192
rect 168432 46180 168438 46232
rect 169202 46180 169208 46232
rect 169260 46220 169266 46232
rect 463694 46220 463700 46232
rect 169260 46192 463700 46220
rect 169260 46180 169266 46192
rect 463694 46180 463700 46192
rect 463752 46180 463758 46232
rect 148686 44888 148692 44940
rect 148744 44928 148750 44940
rect 201586 44928 201592 44940
rect 148744 44900 201592 44928
rect 148744 44888 148750 44900
rect 201586 44888 201592 44900
rect 201644 44888 201650 44940
rect 60826 44820 60832 44872
rect 60884 44860 60890 44872
rect 136634 44860 136640 44872
rect 60884 44832 136640 44860
rect 60884 44820 60890 44832
rect 136634 44820 136640 44832
rect 136692 44820 136698 44872
rect 154298 44820 154304 44872
rect 154356 44860 154362 44872
rect 273254 44860 273260 44872
rect 154356 44832 273260 44860
rect 154356 44820 154362 44832
rect 273254 44820 273260 44832
rect 273312 44820 273318 44872
rect 146110 43596 146116 43648
rect 146168 43636 146174 43648
rect 166994 43636 167000 43648
rect 146168 43608 167000 43636
rect 146168 43596 146174 43608
rect 166994 43596 167000 43608
rect 167052 43596 167058 43648
rect 151170 43528 151176 43580
rect 151228 43568 151234 43580
rect 233234 43568 233240 43580
rect 151228 43540 233240 43568
rect 151228 43528 151234 43540
rect 233234 43528 233240 43540
rect 233292 43528 233298 43580
rect 162026 43460 162032 43512
rect 162084 43500 162090 43512
rect 361574 43500 361580 43512
rect 162084 43472 361580 43500
rect 162084 43460 162090 43472
rect 361574 43460 361580 43472
rect 361632 43460 361638 43512
rect 74534 43392 74540 43444
rect 74592 43432 74598 43444
rect 112438 43432 112444 43444
rect 74592 43404 112444 43432
rect 74592 43392 74598 43404
rect 112438 43392 112444 43404
rect 112496 43392 112502 43444
rect 164878 43392 164884 43444
rect 164936 43432 164942 43444
rect 426434 43432 426440 43444
rect 164936 43404 426440 43432
rect 164936 43392 164942 43404
rect 426434 43392 426440 43404
rect 426492 43392 426498 43444
rect 155310 42236 155316 42288
rect 155368 42276 155374 42288
rect 292666 42276 292672 42288
rect 155368 42248 292672 42276
rect 155368 42236 155374 42248
rect 292666 42236 292672 42248
rect 292724 42236 292730 42288
rect 156966 42168 156972 42220
rect 157024 42208 157030 42220
rect 307846 42208 307852 42220
rect 157024 42180 307852 42208
rect 157024 42168 157030 42180
rect 307846 42168 307852 42180
rect 307904 42168 307910 42220
rect 171502 42100 171508 42152
rect 171560 42140 171566 42152
rect 498286 42140 498292 42152
rect 171560 42112 498292 42140
rect 171560 42100 171566 42112
rect 498286 42100 498292 42112
rect 498344 42100 498350 42152
rect 174814 42032 174820 42084
rect 174872 42072 174878 42084
rect 538858 42072 538864 42084
rect 174872 42044 538864 42072
rect 174872 42032 174878 42044
rect 538858 42032 538864 42044
rect 538916 42032 538922 42084
rect 138014 41624 138020 41676
rect 138072 41664 138078 41676
rect 142614 41664 142620 41676
rect 138072 41636 142620 41664
rect 138072 41624 138078 41636
rect 142614 41624 142620 41636
rect 142672 41624 142678 41676
rect 154390 40944 154396 40996
rect 154448 40984 154454 40996
rect 276014 40984 276020 40996
rect 154448 40956 276020 40984
rect 154448 40944 154454 40956
rect 276014 40944 276020 40956
rect 276072 40944 276078 40996
rect 158254 40876 158260 40928
rect 158312 40916 158318 40928
rect 322934 40916 322940 40928
rect 158312 40888 322940 40916
rect 158312 40876 158318 40888
rect 322934 40876 322940 40888
rect 322992 40876 322998 40928
rect 166350 40808 166356 40860
rect 166408 40848 166414 40860
rect 427814 40848 427820 40860
rect 166408 40820 427820 40848
rect 166408 40808 166414 40820
rect 427814 40808 427820 40820
rect 427872 40808 427878 40860
rect 173434 40740 173440 40792
rect 173492 40780 173498 40792
rect 516134 40780 516140 40792
rect 173492 40752 516140 40780
rect 173492 40740 173498 40752
rect 516134 40740 516140 40752
rect 516192 40740 516198 40792
rect 13814 40672 13820 40724
rect 13872 40712 13878 40724
rect 132862 40712 132868 40724
rect 13872 40684 132868 40712
rect 13872 40672 13878 40684
rect 132862 40672 132868 40684
rect 132920 40672 132926 40724
rect 177298 40672 177304 40724
rect 177356 40712 177362 40724
rect 554774 40712 554780 40724
rect 177356 40684 554780 40712
rect 177356 40672 177362 40684
rect 554774 40672 554780 40684
rect 554832 40672 554838 40724
rect 144454 39992 144460 40044
rect 144512 40032 144518 40044
rect 145098 40032 145104 40044
rect 144512 40004 145104 40032
rect 144512 39992 144518 40004
rect 145098 39992 145104 40004
rect 145156 39992 145162 40044
rect 152734 39584 152740 39636
rect 152792 39624 152798 39636
rect 251174 39624 251180 39636
rect 152792 39596 251180 39624
rect 152792 39584 152798 39596
rect 251174 39584 251180 39596
rect 251232 39584 251238 39636
rect 160646 39516 160652 39568
rect 160704 39556 160710 39568
rect 357526 39556 357532 39568
rect 160704 39528 357532 39556
rect 160704 39516 160710 39528
rect 357526 39516 357532 39528
rect 357584 39516 357590 39568
rect 169478 39448 169484 39500
rect 169536 39488 169542 39500
rect 477494 39488 477500 39500
rect 169536 39460 477500 39488
rect 169536 39448 169542 39460
rect 477494 39448 477500 39460
rect 477552 39448 477558 39500
rect 170766 39380 170772 39432
rect 170824 39420 170830 39432
rect 484394 39420 484400 39432
rect 170824 39392 484400 39420
rect 170824 39380 170830 39392
rect 484394 39380 484400 39392
rect 484452 39380 484458 39432
rect 31754 39312 31760 39364
rect 31812 39352 31818 39364
rect 133874 39352 133880 39364
rect 31812 39324 133880 39352
rect 31812 39312 31818 39324
rect 133874 39312 133880 39324
rect 133932 39312 133938 39364
rect 145650 39312 145656 39364
rect 145708 39352 145714 39364
rect 168466 39352 168472 39364
rect 145708 39324 168472 39352
rect 145708 39312 145714 39324
rect 168466 39312 168472 39324
rect 168524 39312 168530 39364
rect 174722 39312 174728 39364
rect 174780 39352 174786 39364
rect 534074 39352 534080 39364
rect 174780 39324 534080 39352
rect 174780 39312 174786 39324
rect 534074 39312 534080 39324
rect 534132 39312 534138 39364
rect 154206 38156 154212 38208
rect 154264 38196 154270 38208
rect 267826 38196 267832 38208
rect 154264 38168 267832 38196
rect 154264 38156 154270 38168
rect 267826 38156 267832 38168
rect 267884 38156 267890 38208
rect 164970 38088 164976 38140
rect 165028 38128 165034 38140
rect 368474 38128 368480 38140
rect 165028 38100 368480 38128
rect 165028 38088 165034 38100
rect 368474 38088 368480 38100
rect 368532 38088 368538 38140
rect 170030 38020 170036 38072
rect 170088 38060 170094 38072
rect 488534 38060 488540 38072
rect 170088 38032 488540 38060
rect 170088 38020 170094 38032
rect 488534 38020 488540 38032
rect 488592 38020 488598 38072
rect 173526 37952 173532 38004
rect 173584 37992 173590 38004
rect 527818 37992 527824 38004
rect 173584 37964 527824 37992
rect 173584 37952 173590 37964
rect 527818 37952 527824 37964
rect 527876 37952 527882 38004
rect 38654 37884 38660 37936
rect 38712 37924 38718 37936
rect 135622 37924 135628 37936
rect 38712 37896 135628 37924
rect 38712 37884 38718 37896
rect 135622 37884 135628 37896
rect 135680 37884 135686 37936
rect 175366 37884 175372 37936
rect 175424 37924 175430 37936
rect 552014 37924 552020 37936
rect 175424 37896 552020 37924
rect 175424 37884 175430 37896
rect 552014 37884 552020 37896
rect 552072 37884 552078 37936
rect 135346 37272 135352 37324
rect 135404 37312 135410 37324
rect 142430 37312 142436 37324
rect 135404 37284 142436 37312
rect 135404 37272 135410 37284
rect 142430 37272 142436 37284
rect 142488 37272 142494 37324
rect 147490 36864 147496 36916
rect 147548 36904 147554 36916
rect 191834 36904 191840 36916
rect 147548 36876 191840 36904
rect 147548 36864 147554 36876
rect 191834 36864 191840 36876
rect 191892 36864 191898 36916
rect 148594 36796 148600 36848
rect 148652 36836 148658 36848
rect 205634 36836 205640 36848
rect 148652 36808 205640 36836
rect 148652 36796 148658 36808
rect 205634 36796 205640 36808
rect 205692 36796 205698 36848
rect 156782 36728 156788 36780
rect 156840 36768 156846 36780
rect 303614 36768 303620 36780
rect 156840 36740 303620 36768
rect 156840 36728 156846 36740
rect 303614 36728 303620 36740
rect 303672 36728 303678 36780
rect 170858 36660 170864 36712
rect 170916 36700 170922 36712
rect 490006 36700 490012 36712
rect 170916 36672 490012 36700
rect 170916 36660 170922 36672
rect 490006 36660 490012 36672
rect 490064 36660 490070 36712
rect 171410 36592 171416 36644
rect 171468 36632 171474 36644
rect 502334 36632 502340 36644
rect 171468 36604 502340 36632
rect 171468 36592 171474 36604
rect 502334 36592 502340 36604
rect 502392 36592 502398 36644
rect 145558 36524 145564 36576
rect 145616 36564 145622 36576
rect 170398 36564 170404 36576
rect 145616 36536 170404 36564
rect 145616 36524 145622 36536
rect 170398 36524 170404 36536
rect 170456 36524 170462 36576
rect 176194 36524 176200 36576
rect 176252 36564 176258 36576
rect 558914 36564 558920 36576
rect 176252 36536 558920 36564
rect 176252 36524 176258 36536
rect 558914 36524 558920 36536
rect 558972 36524 558978 36576
rect 151998 35368 152004 35420
rect 152056 35408 152062 35420
rect 266354 35408 266360 35420
rect 152056 35380 266360 35408
rect 152056 35368 152062 35380
rect 266354 35368 266360 35380
rect 266412 35368 266418 35420
rect 158346 35300 158352 35352
rect 158404 35340 158410 35352
rect 321554 35340 321560 35352
rect 158404 35312 321560 35340
rect 158404 35300 158410 35312
rect 321554 35300 321560 35312
rect 321612 35300 321618 35352
rect 169846 35232 169852 35284
rect 169904 35272 169910 35284
rect 491294 35272 491300 35284
rect 169904 35244 491300 35272
rect 169904 35232 169910 35244
rect 491294 35232 491300 35244
rect 491352 35232 491358 35284
rect 53834 35164 53840 35216
rect 53892 35204 53898 35216
rect 135438 35204 135444 35216
rect 53892 35176 135444 35204
rect 53892 35164 53898 35176
rect 135438 35164 135444 35176
rect 135496 35164 135502 35216
rect 177390 35164 177396 35216
rect 177448 35204 177454 35216
rect 576210 35204 576216 35216
rect 177448 35176 576216 35204
rect 177448 35164 177454 35176
rect 576210 35164 576216 35176
rect 576268 35164 576274 35216
rect 155678 34008 155684 34060
rect 155736 34048 155742 34060
rect 299566 34048 299572 34060
rect 155736 34020 299572 34048
rect 155736 34008 155742 34020
rect 299566 34008 299572 34020
rect 299624 34008 299630 34060
rect 163406 33940 163412 33992
rect 163464 33980 163470 33992
rect 340966 33980 340972 33992
rect 163464 33952 340972 33980
rect 163464 33940 163470 33952
rect 340966 33940 340972 33952
rect 341024 33940 341030 33992
rect 162210 33872 162216 33924
rect 162268 33912 162274 33924
rect 385034 33912 385040 33924
rect 162268 33884 385040 33912
rect 162268 33872 162274 33884
rect 385034 33872 385040 33884
rect 385092 33872 385098 33924
rect 167914 33804 167920 33856
rect 167972 33844 167978 33856
rect 460934 33844 460940 33856
rect 167972 33816 460940 33844
rect 167972 33804 167978 33816
rect 460934 33804 460940 33816
rect 460992 33804 460998 33856
rect 170490 33736 170496 33788
rect 170548 33776 170554 33788
rect 495434 33776 495440 33788
rect 170548 33748 495440 33776
rect 170548 33736 170554 33748
rect 495434 33736 495440 33748
rect 495492 33736 495498 33788
rect 147582 32648 147588 32700
rect 147640 32688 147646 32700
rect 194594 32688 194600 32700
rect 147640 32660 194600 32688
rect 147640 32648 147646 32660
rect 194594 32648 194600 32660
rect 194652 32648 194658 32700
rect 154114 32580 154120 32632
rect 154172 32620 154178 32632
rect 278774 32620 278780 32632
rect 154172 32592 278780 32620
rect 154172 32580 154178 32592
rect 278774 32580 278780 32592
rect 278832 32580 278838 32632
rect 160922 32512 160928 32564
rect 160980 32552 160986 32564
rect 356698 32552 356704 32564
rect 160980 32524 356704 32552
rect 160980 32512 160986 32524
rect 356698 32512 356704 32524
rect 356756 32512 356762 32564
rect 166442 32444 166448 32496
rect 166500 32484 166506 32496
rect 431954 32484 431960 32496
rect 166500 32456 431960 32484
rect 166500 32444 166506 32456
rect 431954 32444 431960 32456
rect 432012 32444 432018 32496
rect 172606 32376 172612 32428
rect 172664 32416 172670 32428
rect 531406 32416 531412 32428
rect 172664 32388 531412 32416
rect 172664 32376 172670 32388
rect 531406 32376 531412 32388
rect 531464 32376 531470 32428
rect 157150 31288 157156 31340
rect 157208 31328 157214 31340
rect 317414 31328 317420 31340
rect 157208 31300 317420 31328
rect 157208 31288 157214 31300
rect 317414 31288 317420 31300
rect 317472 31288 317478 31340
rect 159910 31220 159916 31272
rect 159968 31260 159974 31272
rect 350534 31260 350540 31272
rect 159968 31232 350540 31260
rect 159968 31220 159974 31232
rect 350534 31220 350540 31232
rect 350592 31220 350598 31272
rect 164234 31152 164240 31204
rect 164292 31192 164298 31204
rect 420914 31192 420920 31204
rect 164292 31164 420920 31192
rect 164292 31152 164298 31164
rect 420914 31152 420920 31164
rect 420972 31152 420978 31204
rect 169662 31084 169668 31136
rect 169720 31124 169726 31136
rect 474734 31124 474740 31136
rect 169720 31096 474740 31124
rect 169720 31084 169726 31096
rect 474734 31084 474740 31096
rect 474792 31084 474798 31136
rect 44266 31016 44272 31068
rect 44324 31056 44330 31068
rect 135530 31056 135536 31068
rect 44324 31028 135536 31056
rect 44324 31016 44330 31028
rect 135530 31016 135536 31028
rect 135588 31016 135594 31068
rect 177666 31016 177672 31068
rect 177724 31056 177730 31068
rect 571978 31056 571984 31068
rect 177724 31028 571984 31056
rect 177724 31016 177730 31028
rect 571978 31016 571984 31028
rect 572036 31016 572042 31068
rect 158438 29792 158444 29844
rect 158496 29832 158502 29844
rect 332686 29832 332692 29844
rect 158496 29804 332692 29832
rect 158496 29792 158502 29804
rect 332686 29792 332692 29804
rect 332744 29792 332750 29844
rect 162302 29724 162308 29776
rect 162360 29764 162366 29776
rect 378778 29764 378784 29776
rect 162360 29736 378784 29764
rect 162360 29724 162366 29736
rect 378778 29724 378784 29736
rect 378836 29724 378842 29776
rect 168006 29656 168012 29708
rect 168064 29696 168070 29708
rect 452654 29696 452660 29708
rect 168064 29668 452660 29696
rect 168064 29656 168070 29668
rect 452654 29656 452660 29668
rect 452712 29656 452718 29708
rect 171318 29588 171324 29640
rect 171376 29628 171382 29640
rect 506566 29628 506572 29640
rect 171376 29600 506572 29628
rect 171376 29588 171382 29600
rect 506566 29588 506572 29600
rect 506624 29588 506630 29640
rect 152642 28500 152648 28552
rect 152700 28540 152706 28552
rect 258074 28540 258080 28552
rect 152700 28512 258080 28540
rect 152700 28500 152706 28512
rect 258074 28500 258080 28512
rect 258132 28500 258138 28552
rect 159818 28432 159824 28484
rect 159876 28472 159882 28484
rect 339494 28472 339500 28484
rect 159876 28444 339500 28472
rect 159876 28432 159882 28444
rect 339494 28432 339500 28444
rect 339552 28432 339558 28484
rect 163866 28364 163872 28416
rect 163924 28404 163930 28416
rect 397454 28404 397460 28416
rect 163924 28376 397460 28404
rect 163924 28364 163930 28376
rect 397454 28364 397460 28376
rect 397512 28364 397518 28416
rect 169570 28296 169576 28348
rect 169628 28336 169634 28348
rect 470594 28336 470600 28348
rect 169628 28308 470600 28336
rect 169628 28296 169634 28308
rect 470594 28296 470600 28308
rect 470652 28296 470658 28348
rect 171226 28228 171232 28280
rect 171284 28268 171290 28280
rect 509234 28268 509240 28280
rect 171284 28240 509240 28268
rect 171284 28228 171290 28240
rect 509234 28228 509240 28240
rect 509292 28228 509298 28280
rect 165154 27072 165160 27124
rect 165212 27112 165218 27124
rect 409874 27112 409880 27124
rect 165212 27084 409880 27112
rect 165212 27072 165218 27084
rect 409874 27072 409880 27084
rect 409932 27072 409938 27124
rect 180702 27004 180708 27056
rect 180760 27044 180766 27056
rect 429194 27044 429200 27056
rect 180760 27016 429200 27044
rect 180760 27004 180766 27016
rect 429194 27004 429200 27016
rect 429252 27004 429258 27056
rect 171870 26936 171876 26988
rect 171928 26976 171934 26988
rect 513374 26976 513380 26988
rect 171928 26948 513380 26976
rect 171928 26936 171934 26948
rect 513374 26936 513380 26948
rect 513432 26936 513438 26988
rect 174906 26868 174912 26920
rect 174964 26908 174970 26920
rect 535454 26908 535460 26920
rect 174964 26880 535460 26908
rect 174964 26868 174970 26880
rect 535454 26868 535460 26880
rect 535512 26868 535518 26920
rect 156690 25780 156696 25832
rect 156748 25820 156754 25832
rect 310514 25820 310520 25832
rect 156748 25792 310520 25820
rect 156748 25780 156754 25792
rect 310514 25780 310520 25792
rect 310572 25780 310578 25832
rect 181622 25712 181628 25764
rect 181680 25752 181686 25764
rect 436094 25752 436100 25764
rect 181680 25724 436100 25752
rect 181680 25712 181686 25724
rect 436094 25712 436100 25724
rect 436152 25712 436158 25764
rect 173710 25644 173716 25696
rect 173768 25684 173774 25696
rect 520274 25684 520280 25696
rect 173768 25656 520280 25684
rect 173768 25644 173774 25656
rect 520274 25644 520280 25656
rect 520332 25644 520338 25696
rect 174998 25576 175004 25628
rect 175056 25616 175062 25628
rect 546494 25616 546500 25628
rect 175056 25588 546500 25616
rect 175056 25576 175062 25588
rect 546494 25576 546500 25588
rect 546552 25576 546558 25628
rect 145006 25508 145012 25560
rect 145064 25548 145070 25560
rect 171778 25548 171784 25560
rect 145064 25520 171784 25548
rect 145064 25508 145070 25520
rect 171778 25508 171784 25520
rect 171836 25508 171842 25560
rect 177758 25508 177764 25560
rect 177816 25548 177822 25560
rect 571334 25548 571340 25560
rect 177816 25520 571340 25548
rect 177816 25508 177822 25520
rect 571334 25508 571340 25520
rect 571392 25508 571398 25560
rect 154022 24352 154028 24404
rect 154080 24392 154086 24404
rect 284386 24392 284392 24404
rect 154080 24364 284392 24392
rect 154080 24352 154086 24364
rect 284386 24352 284392 24364
rect 284444 24352 284450 24404
rect 157334 24284 157340 24336
rect 157392 24324 157398 24336
rect 328454 24324 328460 24336
rect 157392 24296 328460 24324
rect 157392 24284 157398 24296
rect 328454 24284 328460 24296
rect 328512 24284 328518 24336
rect 168190 24216 168196 24268
rect 168248 24256 168254 24268
rect 449894 24256 449900 24268
rect 168248 24228 449900 24256
rect 168248 24216 168254 24228
rect 449894 24216 449900 24228
rect 449952 24216 449958 24268
rect 172514 24148 172520 24200
rect 172572 24188 172578 24200
rect 527174 24188 527180 24200
rect 172572 24160 527180 24188
rect 172572 24148 172578 24160
rect 527174 24148 527180 24160
rect 527232 24148 527238 24200
rect 176286 24080 176292 24132
rect 176344 24120 176350 24132
rect 564526 24120 564532 24132
rect 176344 24092 564532 24120
rect 176344 24080 176350 24092
rect 564526 24080 564532 24092
rect 564584 24080 564590 24132
rect 150066 22992 150072 23044
rect 150124 23032 150130 23044
rect 219434 23032 219440 23044
rect 150124 23004 219440 23032
rect 150124 22992 150130 23004
rect 219434 22992 219440 23004
rect 219492 22992 219498 23044
rect 161106 22924 161112 22976
rect 161164 22964 161170 22976
rect 365806 22964 365812 22976
rect 161164 22936 365812 22964
rect 161164 22924 161170 22936
rect 365806 22924 365812 22936
rect 365864 22924 365870 22976
rect 165246 22856 165252 22908
rect 165304 22896 165310 22908
rect 416774 22896 416780 22908
rect 165304 22868 416780 22896
rect 165304 22856 165310 22868
rect 416774 22856 416780 22868
rect 416832 22856 416838 22908
rect 173986 22788 173992 22840
rect 174044 22828 174050 22840
rect 538214 22828 538220 22840
rect 174044 22800 538220 22828
rect 174044 22788 174050 22800
rect 538214 22788 538220 22800
rect 538272 22788 538278 22840
rect 177850 22720 177856 22772
rect 177908 22760 177914 22772
rect 580258 22760 580264 22772
rect 177908 22732 580264 22760
rect 177908 22720 177914 22732
rect 580258 22720 580264 22732
rect 580316 22720 580322 22772
rect 158530 21632 158536 21684
rect 158588 21672 158594 21684
rect 329098 21672 329104 21684
rect 158588 21644 329104 21672
rect 158588 21632 158594 21644
rect 329098 21632 329104 21644
rect 329156 21632 329162 21684
rect 158162 21564 158168 21616
rect 158220 21604 158226 21616
rect 336734 21604 336740 21616
rect 158220 21576 336740 21604
rect 158220 21564 158226 21576
rect 336734 21564 336740 21576
rect 336792 21564 336798 21616
rect 337378 21564 337384 21616
rect 337436 21604 337442 21616
rect 471974 21604 471980 21616
rect 337436 21576 471980 21604
rect 337436 21564 337442 21576
rect 471974 21564 471980 21576
rect 472032 21564 472038 21616
rect 158806 21496 158812 21548
rect 158864 21536 158870 21548
rect 342898 21536 342904 21548
rect 158864 21508 342904 21536
rect 158864 21496 158870 21508
rect 342898 21496 342904 21508
rect 342956 21496 342962 21548
rect 178770 21428 178776 21480
rect 178828 21468 178834 21480
rect 415486 21468 415492 21480
rect 178828 21440 415492 21468
rect 178828 21428 178834 21440
rect 415486 21428 415492 21440
rect 415544 21428 415550 21480
rect 166626 21360 166632 21412
rect 166684 21400 166690 21412
rect 440326 21400 440332 21412
rect 166684 21372 440332 21400
rect 166684 21360 166690 21372
rect 440326 21360 440332 21372
rect 440384 21360 440390 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 187878 20652 187884 20664
rect 3476 20624 187884 20652
rect 3476 20612 3482 20624
rect 187878 20612 187884 20624
rect 187936 20612 187942 20664
rect 485038 20612 485044 20664
rect 485096 20652 485102 20664
rect 579982 20652 579988 20664
rect 485096 20624 579988 20652
rect 485096 20612 485102 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 154482 20204 154488 20256
rect 154540 20244 154546 20256
rect 280154 20244 280160 20256
rect 154540 20216 280160 20244
rect 154540 20204 154546 20216
rect 280154 20204 280160 20216
rect 280212 20204 280218 20256
rect 155770 20136 155776 20188
rect 155828 20176 155834 20188
rect 291194 20176 291200 20188
rect 155828 20148 291200 20176
rect 155828 20136 155834 20148
rect 291194 20136 291200 20148
rect 291252 20136 291258 20188
rect 155218 20068 155224 20120
rect 155276 20108 155282 20120
rect 287054 20108 287060 20120
rect 155276 20080 287060 20108
rect 155276 20068 155282 20080
rect 287054 20068 287060 20080
rect 287112 20068 287118 20120
rect 287698 20068 287704 20120
rect 287756 20108 287762 20120
rect 465166 20108 465172 20120
rect 287756 20080 465172 20108
rect 287756 20068 287762 20080
rect 465166 20068 465172 20080
rect 465224 20068 465230 20120
rect 161198 20000 161204 20052
rect 161256 20040 161262 20052
rect 372614 20040 372620 20052
rect 161256 20012 372620 20040
rect 161256 20000 161262 20012
rect 372614 20000 372620 20012
rect 372672 20000 372678 20052
rect 143626 19932 143632 19984
rect 143684 19972 143690 19984
rect 154574 19972 154580 19984
rect 143684 19944 154580 19972
rect 143684 19932 143690 19944
rect 154574 19932 154580 19944
rect 154632 19932 154638 19984
rect 182910 19932 182916 19984
rect 182968 19972 182974 19984
rect 442994 19972 443000 19984
rect 182968 19944 443000 19972
rect 182968 19932 182974 19944
rect 442994 19932 443000 19944
rect 443052 19932 443058 19984
rect 149054 18844 149060 18896
rect 149112 18884 149118 18896
rect 226334 18884 226340 18896
rect 149112 18856 226340 18884
rect 149112 18844 149118 18856
rect 226334 18844 226340 18856
rect 226392 18844 226398 18896
rect 155862 18776 155868 18828
rect 155920 18816 155926 18828
rect 300854 18816 300860 18828
rect 155920 18788 300860 18816
rect 155920 18776 155926 18788
rect 300854 18776 300860 18788
rect 300912 18776 300918 18828
rect 176378 18708 176384 18760
rect 176436 18748 176442 18760
rect 529198 18748 529204 18760
rect 176436 18720 529204 18748
rect 176436 18708 176442 18720
rect 529198 18708 529204 18720
rect 529256 18708 529262 18760
rect 175918 18640 175924 18692
rect 175976 18680 175982 18692
rect 567194 18680 567200 18692
rect 175976 18652 567200 18680
rect 175976 18640 175982 18652
rect 567194 18640 567200 18652
rect 567252 18640 567258 18692
rect 177942 18572 177948 18624
rect 178000 18612 178006 18624
rect 574094 18612 574100 18624
rect 178000 18584 574100 18612
rect 178000 18572 178006 18584
rect 574094 18572 574100 18584
rect 574152 18572 574158 18624
rect 151630 17484 151636 17536
rect 151688 17524 151694 17536
rect 241514 17524 241520 17536
rect 151688 17496 241520 17524
rect 151688 17484 151694 17496
rect 241514 17484 241520 17496
rect 241572 17484 241578 17536
rect 165338 17416 165344 17468
rect 165396 17456 165402 17468
rect 425054 17456 425060 17468
rect 165396 17428 425060 17456
rect 165396 17416 165402 17428
rect 425054 17416 425060 17428
rect 425112 17416 425118 17468
rect 166534 17348 166540 17400
rect 166592 17388 166598 17400
rect 441614 17388 441620 17400
rect 166592 17360 441620 17388
rect 166592 17348 166598 17360
rect 441614 17348 441620 17360
rect 441672 17348 441678 17400
rect 168098 17280 168104 17332
rect 168156 17320 168162 17332
rect 445754 17320 445760 17332
rect 168156 17292 445760 17320
rect 168156 17280 168162 17292
rect 445754 17280 445760 17292
rect 445812 17280 445818 17332
rect 146202 17212 146208 17264
rect 146260 17252 146266 17264
rect 165614 17252 165620 17264
rect 146260 17224 165620 17252
rect 146260 17212 146266 17224
rect 165614 17212 165620 17224
rect 165672 17212 165678 17264
rect 170950 17212 170956 17264
rect 171008 17252 171014 17264
rect 492674 17252 492680 17264
rect 171008 17224 492680 17252
rect 171008 17212 171014 17224
rect 492674 17212 492680 17224
rect 492732 17212 492738 17264
rect 152550 16056 152556 16108
rect 152608 16096 152614 16108
rect 252370 16096 252376 16108
rect 152608 16068 252376 16096
rect 152608 16056 152614 16068
rect 252370 16056 252376 16068
rect 252428 16056 252434 16108
rect 161290 15988 161296 16040
rect 161348 16028 161354 16040
rect 361114 16028 361120 16040
rect 161348 16000 361120 16028
rect 161348 15988 161354 16000
rect 361114 15988 361120 16000
rect 361172 15988 361178 16040
rect 161014 15920 161020 15972
rect 161072 15960 161078 15972
rect 364610 15960 364616 15972
rect 161072 15932 364616 15960
rect 161072 15920 161078 15932
rect 364610 15920 364616 15932
rect 364668 15920 364674 15972
rect 400858 15920 400864 15972
rect 400916 15960 400922 15972
rect 478874 15960 478880 15972
rect 400916 15932 478880 15960
rect 400916 15920 400922 15932
rect 478874 15920 478880 15932
rect 478932 15920 478938 15972
rect 166810 15852 166816 15904
rect 166868 15892 166874 15904
rect 432046 15892 432052 15904
rect 166868 15864 432052 15892
rect 166868 15852 166874 15864
rect 432046 15852 432052 15864
rect 432104 15852 432110 15904
rect 153930 14696 153936 14748
rect 153988 14736 153994 14748
rect 272426 14736 272432 14748
rect 153988 14708 272432 14736
rect 153988 14696 153994 14708
rect 272426 14696 272432 14708
rect 272484 14696 272490 14748
rect 155954 14628 155960 14680
rect 156012 14668 156018 14680
rect 314654 14668 314660 14680
rect 156012 14640 314660 14668
rect 156012 14628 156018 14640
rect 314654 14628 314660 14640
rect 314712 14628 314718 14680
rect 163958 14560 163964 14612
rect 164016 14600 164022 14612
rect 398926 14600 398932 14612
rect 164016 14572 398932 14600
rect 164016 14560 164022 14572
rect 398926 14560 398932 14572
rect 398984 14560 398990 14612
rect 164142 14492 164148 14544
rect 164200 14532 164206 14544
rect 404354 14532 404360 14544
rect 164200 14504 404360 14532
rect 164200 14492 164206 14504
rect 404354 14492 404360 14504
rect 404412 14492 404418 14544
rect 172238 14424 172244 14476
rect 172296 14464 172302 14476
rect 503714 14464 503720 14476
rect 172296 14436 503720 14464
rect 172296 14424 172302 14436
rect 503714 14424 503720 14436
rect 503772 14424 503778 14476
rect 157978 13200 157984 13252
rect 158036 13240 158042 13252
rect 324406 13240 324412 13252
rect 158036 13212 324412 13240
rect 158036 13200 158042 13212
rect 324406 13200 324412 13212
rect 324464 13200 324470 13252
rect 164050 13132 164056 13184
rect 164108 13172 164114 13184
rect 407206 13172 407212 13184
rect 164108 13144 407212 13172
rect 164108 13132 164114 13144
rect 407206 13132 407212 13144
rect 407264 13132 407270 13184
rect 172330 13064 172336 13116
rect 172388 13104 172394 13116
rect 511258 13104 511264 13116
rect 172388 13076 511264 13104
rect 172388 13064 172394 13076
rect 511258 13064 511264 13076
rect 511316 13064 511322 13116
rect 151446 11976 151452 12028
rect 151504 12016 151510 12028
rect 245194 12016 245200 12028
rect 151504 11988 245200 12016
rect 151504 11976 151510 11988
rect 245194 11976 245200 11988
rect 245252 11976 245258 12028
rect 160002 11908 160008 11960
rect 160060 11948 160066 11960
rect 342898 11948 342904 11960
rect 160060 11920 342904 11948
rect 160060 11908 160066 11920
rect 342898 11908 342904 11920
rect 342956 11908 342962 11960
rect 162486 11840 162492 11892
rect 162544 11880 162550 11892
rect 390646 11880 390652 11892
rect 162544 11852 390652 11880
rect 162544 11840 162550 11852
rect 390646 11840 390652 11852
rect 390704 11840 390710 11892
rect 166718 11772 166724 11824
rect 166776 11812 166782 11824
rect 435082 11812 435088 11824
rect 166776 11784 435088 11812
rect 166776 11772 166782 11784
rect 435082 11772 435088 11784
rect 435140 11772 435146 11824
rect 174538 11704 174544 11756
rect 174596 11744 174602 11756
rect 548610 11744 548616 11756
rect 174596 11716 548616 11744
rect 174596 11704 174602 11716
rect 548610 11704 548616 11716
rect 548668 11704 548674 11756
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 151078 10480 151084 10532
rect 151136 10520 151142 10532
rect 234614 10520 234620 10532
rect 151136 10492 234620 10520
rect 151136 10480 151142 10492
rect 234614 10480 234620 10492
rect 234672 10480 234678 10532
rect 159634 10412 159640 10464
rect 159692 10452 159698 10464
rect 349246 10452 349252 10464
rect 159692 10424 349252 10452
rect 159692 10412 159698 10424
rect 349246 10412 349252 10424
rect 349304 10412 349310 10464
rect 166902 10344 166908 10396
rect 166960 10384 166966 10396
rect 439130 10384 439136 10396
rect 166960 10356 439136 10384
rect 166960 10344 166966 10356
rect 439130 10344 439136 10356
rect 439188 10344 439194 10396
rect 105722 10276 105728 10328
rect 105780 10316 105786 10328
rect 139578 10316 139584 10328
rect 105780 10288 139584 10316
rect 105780 10276 105786 10288
rect 139578 10276 139584 10288
rect 139636 10276 139642 10328
rect 175274 10276 175280 10328
rect 175332 10316 175338 10328
rect 563054 10316 563060 10328
rect 175332 10288 563060 10316
rect 175332 10276 175338 10288
rect 563054 10276 563060 10288
rect 563112 10276 563118 10328
rect 142798 9596 142804 9648
rect 142856 9636 142862 9648
rect 143534 9636 143540 9648
rect 142856 9608 143540 9636
rect 142856 9596 142862 9608
rect 143534 9596 143540 9608
rect 143592 9596 143598 9648
rect 150342 9188 150348 9240
rect 150400 9228 150406 9240
rect 227530 9228 227536 9240
rect 150400 9200 227536 9228
rect 150400 9188 150406 9200
rect 227530 9188 227536 9200
rect 227588 9188 227594 9240
rect 161382 9120 161388 9172
rect 161440 9160 161446 9172
rect 371694 9160 371700 9172
rect 161440 9132 371700 9160
rect 161440 9120 161446 9132
rect 371694 9120 371700 9132
rect 371752 9120 371758 9172
rect 162578 9052 162584 9104
rect 162636 9092 162642 9104
rect 387150 9092 387156 9104
rect 162636 9064 387156 9092
rect 162636 9052 162642 9064
rect 387150 9052 387156 9064
rect 387208 9052 387214 9104
rect 168282 8984 168288 9036
rect 168340 9024 168346 9036
rect 456886 9024 456892 9036
rect 168340 8996 456892 9024
rect 168340 8984 168346 8996
rect 456886 8984 456892 8996
rect 456944 8984 456950 9036
rect 87966 8916 87972 8968
rect 88024 8956 88030 8968
rect 138198 8956 138204 8968
rect 88024 8928 138204 8956
rect 88024 8916 88030 8928
rect 138198 8916 138204 8928
rect 138256 8916 138262 8968
rect 176562 8916 176568 8968
rect 176620 8956 176626 8968
rect 556154 8956 556160 8968
rect 176620 8928 556160 8956
rect 176620 8916 176626 8928
rect 556154 8916 556160 8928
rect 556212 8916 556218 8968
rect 157242 7760 157248 7812
rect 157300 7800 157306 7812
rect 316218 7800 316224 7812
rect 157300 7772 316224 7800
rect 157300 7760 157306 7772
rect 316218 7760 316224 7772
rect 316276 7760 316282 7812
rect 162394 7692 162400 7744
rect 162452 7732 162458 7744
rect 378870 7732 378876 7744
rect 162452 7704 378876 7732
rect 162452 7692 162458 7704
rect 378870 7692 378876 7704
rect 378928 7692 378934 7744
rect 118694 7624 118700 7676
rect 118752 7664 118758 7676
rect 119890 7664 119896 7676
rect 118752 7636 119896 7664
rect 118752 7624 118758 7636
rect 119890 7624 119896 7636
rect 119948 7624 119954 7676
rect 169754 7624 169760 7676
rect 169812 7664 169818 7676
rect 482830 7664 482836 7676
rect 169812 7636 482836 7664
rect 169812 7624 169818 7636
rect 482830 7624 482836 7636
rect 482888 7624 482894 7676
rect 30098 7556 30104 7608
rect 30156 7596 30162 7608
rect 134150 7596 134156 7608
rect 30156 7568 134156 7596
rect 30156 7556 30162 7568
rect 134150 7556 134156 7568
rect 134208 7556 134214 7608
rect 175090 7556 175096 7608
rect 175148 7596 175154 7608
rect 545482 7596 545488 7608
rect 175148 7568 545488 7596
rect 175148 7556 175154 7568
rect 545482 7556 545488 7568
rect 545540 7556 545546 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 13078 6848 13084 6860
rect 3476 6820 13084 6848
rect 3476 6808 3482 6820
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 576118 6808 576124 6860
rect 576176 6848 576182 6860
rect 580166 6848 580172 6860
rect 576176 6820 580172 6848
rect 576176 6808 576182 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 153838 6332 153844 6384
rect 153896 6372 153902 6384
rect 276014 6372 276020 6384
rect 153896 6344 276020 6372
rect 153896 6332 153902 6344
rect 276014 6332 276020 6344
rect 276072 6332 276078 6384
rect 165522 6264 165528 6316
rect 165580 6304 165586 6316
rect 411898 6304 411904 6316
rect 165580 6276 411904 6304
rect 165580 6264 165586 6276
rect 411898 6264 411904 6276
rect 411956 6264 411962 6316
rect 165430 6196 165436 6248
rect 165488 6236 165494 6248
rect 414290 6236 414296 6248
rect 165488 6208 414296 6236
rect 165488 6196 165494 6208
rect 414290 6196 414296 6208
rect 414348 6196 414354 6248
rect 103330 6128 103336 6180
rect 103388 6168 103394 6180
rect 140314 6168 140320 6180
rect 103388 6140 140320 6168
rect 103388 6128 103394 6140
rect 140314 6128 140320 6140
rect 140372 6128 140378 6180
rect 173802 6128 173808 6180
rect 173860 6168 173866 6180
rect 525426 6168 525432 6180
rect 173860 6140 525432 6168
rect 173860 6128 173866 6140
rect 525426 6128 525432 6140
rect 525484 6128 525490 6180
rect 152366 5040 152372 5092
rect 152424 5080 152430 5092
rect 259546 5080 259552 5092
rect 152424 5052 259552 5080
rect 152424 5040 152430 5052
rect 259546 5040 259552 5052
rect 259604 5040 259610 5092
rect 162670 4972 162676 5024
rect 162728 5012 162734 5024
rect 382366 5012 382372 5024
rect 162728 4984 382372 5012
rect 162728 4972 162734 4984
rect 382366 4972 382372 4984
rect 382424 4972 382430 5024
rect 180150 4904 180156 4956
rect 180208 4944 180214 4956
rect 422570 4944 422576 4956
rect 180208 4916 422576 4944
rect 180208 4904 180214 4916
rect 422570 4904 422576 4916
rect 422628 4904 422634 4956
rect 171042 4836 171048 4888
rect 171100 4876 171106 4888
rect 486326 4876 486332 4888
rect 171100 4848 486332 4876
rect 171100 4836 171106 4848
rect 486326 4836 486332 4848
rect 486384 4836 486390 4888
rect 144822 4768 144828 4820
rect 144880 4808 144886 4820
rect 158898 4808 158904 4820
rect 144880 4780 158904 4808
rect 144880 4768 144886 4780
rect 158898 4768 158904 4780
rect 158956 4768 158962 4820
rect 175182 4768 175188 4820
rect 175240 4808 175246 4820
rect 541986 4808 541992 4820
rect 175240 4780 541992 4808
rect 175240 4768 175246 4780
rect 541986 4768 541992 4780
rect 542044 4768 542050 4820
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 118786 4088 118792 4140
rect 118844 4128 118850 4140
rect 121454 4128 121460 4140
rect 118844 4100 121460 4128
rect 118844 4088 118850 4100
rect 121454 4088 121460 4100
rect 121512 4088 121518 4140
rect 123478 4088 123484 4140
rect 123536 4128 123542 4140
rect 124950 4128 124956 4140
rect 123536 4100 124956 4128
rect 123536 4088 123542 4100
rect 124950 4088 124956 4100
rect 125008 4088 125014 4140
rect 131850 4128 131856 4140
rect 125060 4100 131856 4128
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 8938 4060 8944 4072
rect 1728 4032 8944 4060
rect 1728 4020 1734 4032
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 122282 4020 122288 4072
rect 122340 4060 122346 4072
rect 124858 4060 124864 4072
rect 122340 4032 124864 4060
rect 122340 4020 122346 4032
rect 124858 4020 124864 4032
rect 124916 4020 124922 4072
rect 125060 3992 125088 4100
rect 131850 4088 131856 4100
rect 131908 4088 131914 4140
rect 301590 4088 301596 4140
rect 301648 4128 301654 4140
rect 309042 4128 309048 4140
rect 301648 4100 309048 4128
rect 301648 4088 301654 4100
rect 309042 4088 309048 4100
rect 309100 4088 309106 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 317322 4128 317328 4140
rect 315356 4100 317328 4128
rect 315356 4088 315362 4100
rect 317322 4088 317328 4100
rect 317380 4088 317386 4140
rect 450538 4088 450544 4140
rect 450596 4128 450602 4140
rect 450998 4128 451004 4140
rect 450596 4100 451004 4128
rect 450596 4088 450602 4100
rect 450998 4088 451004 4100
rect 451056 4088 451062 4140
rect 527910 4088 527916 4140
rect 527968 4128 527974 4140
rect 529014 4128 529020 4140
rect 527968 4100 529020 4128
rect 527968 4088 527974 4100
rect 529014 4088 529020 4100
rect 529072 4088 529078 4140
rect 576210 4088 576216 4140
rect 576268 4128 576274 4140
rect 577406 4128 577412 4140
rect 576268 4100 577412 4128
rect 576268 4088 576274 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 125870 4020 125876 4072
rect 125928 4060 125934 4072
rect 129918 4060 129924 4072
rect 125928 4032 129924 4060
rect 125928 4020 125934 4032
rect 129918 4020 129924 4032
rect 129976 4020 129982 4072
rect 203610 4020 203616 4072
rect 203668 4060 203674 4072
rect 203668 4032 219434 4060
rect 203668 4020 203674 4032
rect 134518 3992 134524 4004
rect 118666 3964 125088 3992
rect 128326 3964 134524 3992
rect 45922 3884 45928 3936
rect 45980 3924 45986 3936
rect 46198 3924 46204 3936
rect 45980 3896 46204 3924
rect 45980 3884 45986 3896
rect 46198 3884 46204 3896
rect 46256 3884 46262 3936
rect 106918 3748 106924 3800
rect 106976 3788 106982 3800
rect 118666 3788 118694 3964
rect 128326 3924 128354 3964
rect 134518 3952 134524 3964
rect 134576 3952 134582 4004
rect 184198 3952 184204 4004
rect 184256 3992 184262 4004
rect 210970 3992 210976 4004
rect 184256 3964 210976 3992
rect 184256 3952 184262 3964
rect 210970 3952 210976 3964
rect 211028 3952 211034 4004
rect 106976 3760 118694 3788
rect 123496 3896 128354 3924
rect 106976 3748 106982 3760
rect 85666 3680 85672 3732
rect 85724 3720 85730 3732
rect 123496 3720 123524 3896
rect 131022 3884 131028 3936
rect 131080 3924 131086 3936
rect 144730 3924 144736 3936
rect 131080 3896 144736 3924
rect 131080 3884 131086 3896
rect 144730 3884 144736 3896
rect 144788 3884 144794 3936
rect 148502 3884 148508 3936
rect 148560 3924 148566 3936
rect 151814 3924 151820 3936
rect 148560 3896 151820 3924
rect 148560 3884 148566 3896
rect 151814 3884 151820 3896
rect 151872 3884 151878 3936
rect 181438 3884 181444 3936
rect 181496 3924 181502 3936
rect 190822 3924 190828 3936
rect 181496 3896 190828 3924
rect 181496 3884 181502 3896
rect 190822 3884 190828 3896
rect 190880 3884 190886 3936
rect 193858 3884 193864 3936
rect 193916 3924 193922 3936
rect 196802 3924 196808 3936
rect 193916 3896 196808 3924
rect 193916 3884 193922 3896
rect 196802 3884 196808 3896
rect 196860 3884 196866 3936
rect 196894 3884 196900 3936
rect 196952 3924 196958 3936
rect 203886 3924 203892 3936
rect 196952 3896 203892 3924
rect 196952 3884 196958 3896
rect 203886 3884 203892 3896
rect 203944 3884 203950 3936
rect 211798 3884 211804 3936
rect 211856 3924 211862 3936
rect 219406 3924 219434 4032
rect 247678 4020 247684 4072
rect 247736 4060 247742 4072
rect 248782 4060 248788 4072
rect 247736 4032 248788 4060
rect 247736 4020 247742 4032
rect 248782 4020 248788 4032
rect 248840 4020 248846 4072
rect 224218 3952 224224 4004
rect 224276 3992 224282 4004
rect 247586 3992 247592 4004
rect 224276 3964 247592 3992
rect 224276 3952 224282 3964
rect 247586 3952 247592 3964
rect 247644 3952 247650 4004
rect 231026 3924 231032 3936
rect 211856 3896 212304 3924
rect 219406 3896 231032 3924
rect 211856 3884 211862 3896
rect 124674 3816 124680 3868
rect 124732 3856 124738 3868
rect 140866 3856 140872 3868
rect 124732 3828 140872 3856
rect 124732 3816 124738 3828
rect 140866 3816 140872 3828
rect 140924 3816 140930 3868
rect 149698 3816 149704 3868
rect 149756 3856 149762 3868
rect 212166 3856 212172 3868
rect 149756 3828 212172 3856
rect 149756 3816 149762 3828
rect 212166 3816 212172 3828
rect 212224 3816 212230 3868
rect 212276 3856 212304 3896
rect 231026 3884 231032 3896
rect 231084 3884 231090 3936
rect 261478 3884 261484 3936
rect 261536 3924 261542 3936
rect 262950 3924 262956 3936
rect 261536 3896 262956 3924
rect 261536 3884 261542 3896
rect 262950 3884 262956 3896
rect 263008 3884 263014 3936
rect 240502 3856 240508 3868
rect 212276 3828 240508 3856
rect 240502 3816 240508 3828
rect 240560 3816 240566 3868
rect 242158 3816 242164 3868
rect 242216 3856 242222 3868
rect 298462 3856 298468 3868
rect 242216 3828 298468 3856
rect 242216 3816 242222 3828
rect 298462 3816 298468 3828
rect 298520 3816 298526 3868
rect 299566 3816 299572 3868
rect 299624 3856 299630 3868
rect 300762 3856 300768 3868
rect 299624 3828 300768 3856
rect 299624 3816 299630 3828
rect 300762 3816 300768 3828
rect 300820 3816 300826 3868
rect 311158 3816 311164 3868
rect 311216 3856 311222 3868
rect 312630 3856 312636 3868
rect 311216 3828 312636 3856
rect 311216 3816 311222 3828
rect 312630 3816 312636 3828
rect 312688 3816 312694 3868
rect 146938 3748 146944 3800
rect 146996 3788 147002 3800
rect 156598 3788 156604 3800
rect 146996 3760 156604 3788
rect 146996 3748 147002 3760
rect 156598 3748 156604 3760
rect 156656 3748 156662 3800
rect 156690 3748 156696 3800
rect 156748 3788 156754 3800
rect 170766 3788 170772 3800
rect 156748 3760 170772 3788
rect 156748 3748 156754 3760
rect 170766 3748 170772 3760
rect 170824 3748 170830 3800
rect 172422 3748 172428 3800
rect 172480 3788 172486 3800
rect 327994 3788 328000 3800
rect 172480 3760 328000 3788
rect 172480 3748 172486 3760
rect 327994 3748 328000 3760
rect 328052 3748 328058 3800
rect 357526 3748 357532 3800
rect 357584 3788 357590 3800
rect 358722 3788 358728 3800
rect 357584 3760 358728 3788
rect 357584 3748 357590 3760
rect 358722 3748 358728 3760
rect 358780 3748 358786 3800
rect 85724 3692 123524 3720
rect 85724 3680 85730 3692
rect 147122 3680 147128 3732
rect 147180 3680 147186 3732
rect 162762 3680 162768 3732
rect 162820 3720 162826 3732
rect 377674 3720 377680 3732
rect 162820 3692 377680 3720
rect 162820 3680 162826 3692
rect 377674 3680 377680 3692
rect 377732 3680 377738 3732
rect 66714 3612 66720 3664
rect 66772 3652 66778 3664
rect 72418 3652 72424 3664
rect 66772 3624 72424 3652
rect 66772 3612 66778 3624
rect 72418 3612 72424 3624
rect 72476 3612 72482 3664
rect 83274 3612 83280 3664
rect 83332 3652 83338 3664
rect 138106 3652 138112 3664
rect 83332 3624 138112 3652
rect 83332 3612 83338 3624
rect 138106 3612 138112 3624
rect 138164 3612 138170 3664
rect 147140 3652 147168 3680
rect 163682 3652 163688 3664
rect 147140 3624 163688 3652
rect 163682 3612 163688 3624
rect 163740 3612 163746 3664
rect 168374 3612 168380 3664
rect 168432 3652 168438 3664
rect 169570 3652 169576 3664
rect 168432 3624 169576 3652
rect 168432 3612 168438 3624
rect 169570 3612 169576 3624
rect 169628 3612 169634 3664
rect 178678 3612 178684 3664
rect 178736 3652 178742 3664
rect 408402 3652 408408 3664
rect 178736 3624 408408 3652
rect 178736 3612 178742 3624
rect 408402 3612 408408 3624
rect 408460 3612 408466 3664
rect 454678 3612 454684 3664
rect 454736 3652 454742 3664
rect 500586 3652 500592 3664
rect 454736 3624 500592 3652
rect 454736 3612 454742 3624
rect 500586 3612 500592 3624
rect 500644 3612 500650 3664
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 21358 3584 21364 3596
rect 19484 3556 21364 3584
rect 19484 3544 19490 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 44174 3544 44180 3596
rect 44232 3584 44238 3596
rect 45094 3584 45100 3596
rect 44232 3556 45100 3584
rect 44232 3544 44238 3556
rect 45094 3544 45100 3556
rect 45152 3544 45158 3596
rect 51350 3544 51356 3596
rect 51408 3584 51414 3596
rect 54478 3584 54484 3596
rect 51408 3556 54484 3584
rect 51408 3544 51414 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 64138 3584 64144 3596
rect 59688 3556 64144 3584
rect 59688 3544 59694 3556
rect 64138 3544 64144 3556
rect 64196 3544 64202 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 69164 3556 123616 3584
rect 69164 3544 69170 3556
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 120718 3516 120724 3528
rect 6512 3488 120724 3516
rect 6512 3476 6518 3488
rect 120718 3476 120724 3488
rect 120776 3476 120782 3528
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 10318 3448 10324 3460
rect 8812 3420 10324 3448
rect 8812 3408 8818 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 18598 3448 18604 3460
rect 17092 3420 18604 3448
rect 17092 3408 17098 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 27614 3408 27620 3460
rect 27672 3448 27678 3460
rect 28534 3448 28540 3460
rect 27672 3420 28540 3448
rect 27672 3408 27678 3420
rect 28534 3408 28540 3420
rect 28592 3408 28598 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 45922 3448 45928 3460
rect 33652 3420 45928 3448
rect 33652 3408 33658 3420
rect 45922 3408 45928 3420
rect 45980 3408 45986 3460
rect 52454 3408 52460 3460
rect 52512 3448 52518 3460
rect 53374 3448 53380 3460
rect 52512 3420 53380 3448
rect 52512 3408 52518 3420
rect 53374 3408 53380 3420
rect 53432 3408 53438 3460
rect 56042 3408 56048 3460
rect 56100 3448 56106 3460
rect 57238 3448 57244 3460
rect 56100 3420 57244 3448
rect 56100 3408 56106 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 60734 3408 60740 3460
rect 60792 3448 60798 3460
rect 61654 3448 61660 3460
rect 60792 3420 61660 3448
rect 60792 3408 60798 3420
rect 61654 3408 61660 3420
rect 61712 3408 61718 3460
rect 65518 3408 65524 3460
rect 65576 3448 65582 3460
rect 123588 3448 123616 3556
rect 128170 3544 128176 3596
rect 128228 3584 128234 3596
rect 130378 3584 130384 3596
rect 128228 3556 130384 3584
rect 128228 3544 128234 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 135254 3544 135260 3596
rect 135312 3584 135318 3596
rect 136450 3584 136456 3596
rect 135312 3556 136456 3584
rect 135312 3544 135318 3556
rect 136450 3544 136456 3556
rect 136508 3544 136514 3596
rect 137646 3544 137652 3596
rect 137704 3584 137710 3596
rect 138658 3584 138664 3596
rect 137704 3556 138664 3584
rect 137704 3544 137710 3556
rect 138658 3544 138664 3556
rect 138716 3544 138722 3596
rect 141418 3544 141424 3596
rect 141476 3584 141482 3596
rect 147122 3584 147128 3596
rect 141476 3556 147128 3584
rect 141476 3544 141482 3556
rect 147122 3544 147128 3556
rect 147180 3544 147186 3596
rect 152458 3544 152464 3596
rect 152516 3584 152522 3596
rect 175458 3584 175464 3596
rect 152516 3556 175464 3584
rect 152516 3544 152522 3556
rect 175458 3544 175464 3556
rect 175516 3544 175522 3596
rect 180058 3544 180064 3596
rect 180116 3544 180122 3596
rect 180334 3544 180340 3596
rect 180392 3584 180398 3596
rect 468294 3584 468300 3596
rect 180392 3556 468300 3584
rect 180392 3544 180398 3556
rect 468294 3544 468300 3556
rect 468352 3544 468358 3596
rect 468478 3544 468484 3596
rect 468536 3584 468542 3596
rect 469858 3584 469864 3596
rect 468536 3556 469864 3584
rect 468536 3544 468542 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 472618 3544 472624 3596
rect 472676 3584 472682 3596
rect 473446 3584 473452 3596
rect 472676 3556 473452 3584
rect 472676 3544 472682 3556
rect 473446 3544 473452 3556
rect 473504 3544 473510 3596
rect 475378 3544 475384 3596
rect 475436 3584 475442 3596
rect 518342 3584 518348 3596
rect 475436 3556 518348 3584
rect 475436 3544 475442 3556
rect 518342 3544 518348 3556
rect 518400 3544 518406 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 533706 3584 533712 3596
rect 525116 3556 533712 3584
rect 525116 3544 525122 3556
rect 533706 3544 533712 3556
rect 533764 3544 533770 3596
rect 538858 3544 538864 3596
rect 538916 3584 538922 3596
rect 539594 3584 539600 3596
rect 538916 3556 539600 3584
rect 538916 3544 538922 3556
rect 539594 3544 539600 3556
rect 539652 3544 539658 3596
rect 545758 3544 545764 3596
rect 545816 3584 545822 3596
rect 551462 3584 551468 3596
rect 545816 3556 551468 3584
rect 545816 3544 545822 3556
rect 551462 3544 551468 3556
rect 551520 3544 551526 3596
rect 572714 3584 572720 3596
rect 567166 3556 572720 3584
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128446 3516 128452 3528
rect 127032 3488 128452 3516
rect 127032 3476 127038 3488
rect 128446 3476 128452 3488
rect 128504 3476 128510 3528
rect 131206 3516 131212 3528
rect 128556 3488 131212 3516
rect 128556 3448 128584 3488
rect 131206 3476 131212 3488
rect 131264 3476 131270 3528
rect 134150 3476 134156 3528
rect 134208 3516 134214 3528
rect 136910 3516 136916 3528
rect 134208 3488 136916 3516
rect 134208 3476 134214 3488
rect 136910 3476 136916 3488
rect 136968 3476 136974 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148376 3488 171640 3516
rect 148376 3476 148382 3488
rect 65576 3420 115934 3448
rect 123588 3420 128584 3448
rect 65576 3408 65582 3420
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 17218 3380 17224 3392
rect 15988 3352 17224 3380
rect 15988 3340 15994 3352
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 77294 3340 77300 3392
rect 77352 3380 77358 3392
rect 78214 3380 78220 3392
rect 77352 3352 78220 3380
rect 77352 3340 77358 3352
rect 78214 3340 78220 3352
rect 78272 3340 78278 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 102778 3380 102784 3392
rect 101088 3352 102784 3380
rect 101088 3340 101094 3352
rect 102778 3340 102784 3352
rect 102836 3340 102842 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 115906 3380 115934 3420
rect 130930 3408 130936 3460
rect 130988 3448 130994 3460
rect 162486 3448 162492 3460
rect 130988 3420 162492 3448
rect 130988 3408 130994 3420
rect 162486 3408 162492 3420
rect 162544 3408 162550 3460
rect 129918 3380 129924 3392
rect 115906 3352 129924 3380
rect 129918 3340 129924 3352
rect 129976 3340 129982 3392
rect 132954 3340 132960 3392
rect 133012 3380 133018 3392
rect 141510 3380 141516 3392
rect 133012 3352 141516 3380
rect 133012 3340 133018 3352
rect 141510 3340 141516 3352
rect 141568 3340 141574 3392
rect 162118 3340 162124 3392
rect 162176 3380 162182 3392
rect 164878 3380 164884 3392
rect 162176 3352 164884 3380
rect 162176 3340 162182 3352
rect 164878 3340 164884 3352
rect 164936 3340 164942 3392
rect 171612 3380 171640 3488
rect 171778 3476 171784 3528
rect 171836 3516 171842 3528
rect 173158 3516 173164 3528
rect 171836 3488 173164 3516
rect 171836 3476 171842 3488
rect 173158 3476 173164 3488
rect 173216 3476 173222 3528
rect 180076 3516 180104 3544
rect 180076 3488 180794 3516
rect 176654 3380 176660 3392
rect 171612 3352 176660 3380
rect 176654 3340 176660 3352
rect 176712 3340 176718 3392
rect 120718 3272 120724 3324
rect 120776 3312 120782 3324
rect 131758 3312 131764 3324
rect 120776 3284 131764 3312
rect 120776 3272 120782 3284
rect 131758 3272 131764 3284
rect 131816 3272 131822 3324
rect 147030 3272 147036 3324
rect 147088 3312 147094 3324
rect 150618 3312 150624 3324
rect 147088 3284 150624 3312
rect 147088 3272 147094 3284
rect 150618 3272 150624 3284
rect 150676 3272 150682 3324
rect 170398 3272 170404 3324
rect 170456 3312 170462 3324
rect 174262 3312 174268 3324
rect 170456 3284 174268 3312
rect 170456 3272 170462 3284
rect 174262 3272 174268 3284
rect 174320 3272 174326 3324
rect 180766 3312 180794 3488
rect 181530 3476 181536 3528
rect 181588 3516 181594 3528
rect 186130 3516 186136 3528
rect 181588 3488 186136 3516
rect 181588 3476 181594 3488
rect 186130 3476 186136 3488
rect 186188 3476 186194 3528
rect 186332 3488 504128 3516
rect 182082 3340 182088 3392
rect 182140 3380 182146 3392
rect 186332 3380 186360 3488
rect 182140 3352 186360 3380
rect 190426 3420 489914 3448
rect 182140 3340 182146 3352
rect 190426 3312 190454 3420
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260650 3380 260656 3392
rect 259512 3352 260656 3380
rect 259512 3340 259518 3352
rect 260650 3340 260656 3352
rect 260708 3340 260714 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 329098 3340 329104 3392
rect 329156 3380 329162 3392
rect 330386 3380 330392 3392
rect 329156 3352 330392 3380
rect 329156 3340 329162 3352
rect 330386 3340 330392 3352
rect 330444 3340 330450 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 342990 3340 342996 3392
rect 343048 3380 343054 3392
rect 344554 3380 344560 3392
rect 343048 3352 344560 3380
rect 343048 3340 343054 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 356698 3340 356704 3392
rect 356756 3380 356762 3392
rect 357526 3380 357532 3392
rect 356756 3352 357532 3380
rect 356756 3340 356762 3352
rect 357526 3340 357532 3352
rect 357584 3340 357590 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 378778 3340 378784 3392
rect 378836 3380 378842 3392
rect 379974 3380 379980 3392
rect 378836 3352 379980 3380
rect 378836 3340 378842 3352
rect 379974 3340 379980 3352
rect 380032 3340 380038 3392
rect 382918 3340 382924 3392
rect 382976 3380 382982 3392
rect 384758 3380 384764 3392
rect 382976 3352 384764 3380
rect 382976 3340 382982 3352
rect 384758 3340 384764 3352
rect 384816 3340 384822 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 416682 3380 416688 3392
rect 414716 3352 416688 3380
rect 414716 3340 414722 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 418798 3340 418804 3392
rect 418856 3380 418862 3392
rect 420178 3380 420184 3392
rect 418856 3352 420184 3380
rect 418856 3340 418862 3352
rect 420178 3340 420184 3352
rect 420236 3340 420242 3392
rect 431954 3340 431960 3392
rect 432012 3380 432018 3392
rect 433242 3380 433248 3392
rect 432012 3352 433248 3380
rect 432012 3340 432018 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 446398 3340 446404 3392
rect 446456 3380 446462 3392
rect 447410 3380 447416 3392
rect 446456 3352 447416 3380
rect 446456 3340 446462 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 453390 3340 453396 3392
rect 453448 3380 453454 3392
rect 454494 3380 454500 3392
rect 453448 3352 454500 3380
rect 453448 3340 453454 3352
rect 454494 3340 454500 3352
rect 454552 3340 454558 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 486418 3340 486424 3392
rect 486476 3380 486482 3392
rect 487614 3380 487620 3392
rect 486476 3352 487620 3380
rect 486476 3340 486482 3352
rect 487614 3340 487620 3352
rect 487672 3340 487678 3392
rect 180766 3284 190454 3312
rect 324958 3272 324964 3324
rect 325016 3312 325022 3324
rect 326798 3312 326804 3324
rect 325016 3284 326804 3312
rect 325016 3272 325022 3284
rect 326798 3272 326804 3284
rect 326856 3272 326862 3324
rect 382274 3272 382280 3324
rect 382332 3312 382338 3324
rect 383562 3312 383568 3324
rect 382332 3284 383568 3312
rect 382332 3272 382338 3284
rect 383562 3272 383568 3284
rect 383620 3272 383626 3324
rect 450998 3272 451004 3324
rect 451056 3312 451062 3324
rect 452102 3312 452108 3324
rect 451056 3284 452108 3312
rect 451056 3272 451062 3284
rect 452102 3272 452108 3284
rect 452160 3272 452166 3324
rect 489886 3312 489914 3420
rect 496078 3408 496084 3460
rect 496136 3448 496142 3460
rect 497090 3448 497096 3460
rect 496136 3420 497096 3448
rect 496136 3408 496142 3420
rect 497090 3408 497096 3420
rect 497148 3408 497154 3460
rect 504100 3380 504128 3488
rect 504358 3476 504364 3528
rect 504416 3516 504422 3528
rect 507670 3516 507676 3528
rect 504416 3488 507676 3516
rect 504416 3476 504422 3488
rect 507670 3476 507676 3488
rect 507728 3476 507734 3528
rect 529198 3476 529204 3528
rect 529256 3516 529262 3528
rect 560846 3516 560852 3528
rect 529256 3488 560852 3516
rect 529256 3476 529262 3488
rect 560846 3476 560852 3488
rect 560904 3476 560910 3528
rect 560938 3476 560944 3528
rect 560996 3516 561002 3528
rect 567166 3516 567194 3556
rect 572714 3544 572720 3556
rect 572772 3544 572778 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 576302 3584 576308 3596
rect 574796 3556 576308 3584
rect 574796 3544 574802 3556
rect 576302 3544 576308 3556
rect 576360 3544 576366 3596
rect 560996 3488 567194 3516
rect 560996 3476 561002 3488
rect 567838 3476 567844 3528
rect 567896 3516 567902 3528
rect 569126 3516 569132 3528
rect 567896 3488 569132 3516
rect 567896 3476 567902 3488
rect 569126 3476 569132 3488
rect 569184 3476 569190 3528
rect 580258 3476 580264 3528
rect 580316 3516 580322 3528
rect 580994 3516 581000 3528
rect 580316 3488 581000 3516
rect 580316 3476 580322 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 583386 3448 583392 3460
rect 509206 3420 583392 3448
rect 505370 3380 505376 3392
rect 504100 3352 505376 3380
rect 505370 3340 505376 3352
rect 505428 3340 505434 3392
rect 509206 3312 509234 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 489886 3284 509234 3312
rect 192478 3204 192484 3256
rect 192536 3244 192542 3256
rect 193214 3244 193220 3256
rect 192536 3216 193220 3244
rect 192536 3204 192542 3216
rect 193214 3204 193220 3216
rect 193272 3204 193278 3256
rect 400950 3204 400956 3256
rect 401008 3244 401014 3256
rect 402514 3244 402520 3256
rect 401008 3216 402520 3244
rect 401008 3204 401014 3216
rect 402514 3204 402520 3216
rect 402572 3204 402578 3256
rect 520918 3204 520924 3256
rect 520976 3244 520982 3256
rect 524230 3244 524236 3256
rect 520976 3216 524236 3244
rect 520976 3204 520982 3216
rect 524230 3204 524236 3216
rect 524288 3204 524294 3256
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 39298 3176 39304 3188
rect 38436 3148 39304 3176
rect 38436 3136 38442 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 511350 3136 511356 3188
rect 511408 3176 511414 3188
rect 514754 3176 514760 3188
rect 511408 3148 514760 3176
rect 511408 3136 511414 3148
rect 514754 3136 514760 3148
rect 514812 3136 514818 3188
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22738 3040 22744 3052
rect 20680 3012 22744 3040
rect 20680 3000 20686 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 23014 3000 23020 3052
rect 23072 3040 23078 3052
rect 25498 3040 25504 3052
rect 23072 3012 25504 3040
rect 23072 3000 23078 3012
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 147214 3000 147220 3052
rect 147272 3040 147278 3052
rect 148318 3040 148324 3052
rect 147272 3012 148324 3040
rect 147272 3000 147278 3012
rect 148318 3000 148324 3012
rect 148376 3000 148382 3052
rect 148410 3000 148416 3052
rect 148468 3040 148474 3052
rect 154206 3040 154212 3052
rect 148468 3012 154212 3040
rect 148468 3000 148474 3012
rect 154206 3000 154212 3012
rect 154264 3000 154270 3052
rect 175918 3000 175924 3052
rect 175976 3040 175982 3052
rect 177850 3040 177856 3052
rect 175976 3012 177856 3040
rect 175976 3000 175982 3012
rect 177850 3000 177856 3012
rect 177908 3000 177914 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 565630 3040 565636 3052
rect 563756 3012 565636 3040
rect 563756 3000 563762 3012
rect 565630 3000 565636 3012
rect 565688 3000 565694 3052
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 14458 2972 14464 2984
rect 12400 2944 14464 2972
rect 12400 2932 12406 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 182818 2932 182824 2984
rect 182876 2972 182882 2984
rect 189718 2972 189724 2984
rect 182876 2944 189724 2972
rect 182876 2932 182882 2944
rect 189718 2932 189724 2944
rect 189776 2932 189782 2984
rect 423674 2864 423680 2916
rect 423732 2904 423738 2916
rect 424962 2904 424968 2916
rect 423732 2876 424968 2904
rect 423732 2864 423738 2876
rect 424962 2864 424968 2876
rect 425020 2864 425026 2916
rect 440234 2592 440240 2644
rect 440292 2632 440298 2644
rect 441522 2632 441528 2644
rect 440292 2604 441528 2632
rect 440292 2592 440298 2604
rect 441522 2592 441528 2604
rect 441580 2592 441586 2644
rect 390554 2456 390560 2508
rect 390612 2496 390618 2508
rect 391842 2496 391848 2508
rect 390612 2468 391848 2496
rect 390612 2456 390618 2468
rect 391842 2456 391848 2468
rect 391900 2456 391906 2508
rect 340874 1776 340880 1828
rect 340932 1816 340938 1828
rect 342162 1816 342168 1828
rect 340932 1788 342168 1816
rect 340932 1776 340938 1788
rect 342162 1776 342168 1788
rect 342220 1776 342226 1828
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 137836 700816 137888 700868
rect 157340 700816 157392 700868
rect 155960 700748 156012 700800
rect 202788 700748 202840 700800
rect 89168 700680 89220 700732
rect 160744 700680 160796 700732
rect 154580 700612 154632 700664
rect 267648 700612 267700 700664
rect 24308 700544 24360 700596
rect 162216 700544 162268 700596
rect 8116 700476 8168 700528
rect 162124 700476 162176 700528
rect 153292 700408 153344 700460
rect 332508 700408 332560 700460
rect 152464 700340 152516 700392
rect 413652 700340 413704 700392
rect 489184 700340 489236 700392
rect 527180 700340 527232 700392
rect 527824 700340 527876 700392
rect 559656 700340 559708 700392
rect 148324 700272 148376 700324
rect 543464 700272 543516 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 146300 696940 146352 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 161480 683204 161532 683256
rect 146944 683136 146996 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 163504 670692 163556 670744
rect 498844 670692 498896 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 163596 656888 163648 656940
rect 182824 643084 182876 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 164240 632068 164292 632120
rect 188344 630640 188396 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 164884 618264 164936 618316
rect 143632 616836 143684 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 164976 605820 165028 605872
rect 142344 590656 142396 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 165620 579640 165672 579692
rect 144184 576852 144236 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 167644 565836 167696 565888
rect 142804 563048 142856 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 166264 553392 166316 553444
rect 181444 536800 181496 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 167000 527144 167052 527196
rect 142896 524424 142948 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 7564 514768 7616 514820
rect 180064 510620 180116 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 167736 500964 167788 501016
rect 139400 484372 139452 484424
rect 580172 484372 580224 484424
rect 140044 470568 140096 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 170404 462340 170456 462392
rect 178684 456764 178736 456816
rect 580172 456764 580224 456816
rect 157432 450508 157484 450560
rect 169760 450508 169812 450560
rect 3148 448536 3200 448588
rect 170496 448536 170548 448588
rect 138664 430584 138716 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 169760 422288 169812 422340
rect 138756 418140 138808 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 171784 409844 171836 409896
rect 185584 404336 185636 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 171876 397468 171928 397520
rect 196624 378156 196676 378208
rect 580172 378156 580224 378208
rect 2780 371288 2832 371340
rect 4804 371288 4856 371340
rect 3516 358368 3568 358420
rect 8944 358368 8996 358420
rect 135260 351908 135312 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 149704 345040 149756 345092
rect 134524 324300 134576 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 173900 318792 173952 318844
rect 135904 311856 135956 311908
rect 579988 311856 580040 311908
rect 3516 304988 3568 305040
rect 175924 304988 175976 305040
rect 134616 298120 134668 298172
rect 580172 298120 580224 298172
rect 3516 292544 3568 292596
rect 174544 292544 174596 292596
rect 145564 289076 145616 289128
rect 188344 289076 188396 289128
rect 149060 287648 149112 287700
rect 462320 287648 462372 287700
rect 137284 286288 137336 286340
rect 196624 286288 196676 286340
rect 147680 283568 147732 283620
rect 489184 283568 489236 283620
rect 144920 282140 144972 282192
rect 182824 282140 182876 282192
rect 140780 280780 140832 280832
rect 181444 280780 181496 280832
rect 40040 279420 40092 279472
rect 160100 279420 160152 279472
rect 151084 275272 151136 275324
rect 428464 275272 428516 275324
rect 8944 273912 8996 273964
rect 173164 273912 173216 273964
rect 186688 273912 186740 273964
rect 364340 273912 364392 273964
rect 151912 273232 151964 273284
rect 186688 273232 186740 273284
rect 187148 273232 187200 273284
rect 133144 271872 133196 271924
rect 580172 271872 580224 271924
rect 7564 271192 7616 271244
rect 169024 271192 169076 271244
rect 149152 271124 149204 271176
rect 494060 271124 494112 271176
rect 71780 269764 71832 269816
rect 119988 269764 120040 269816
rect 147772 269764 147824 269816
rect 527824 269764 527876 269816
rect 119988 269084 120040 269136
rect 158720 269084 158772 269136
rect 4804 268404 4856 268456
rect 172704 268404 172756 268456
rect 146208 268336 146260 268388
rect 498844 268336 498896 268388
rect 137836 266976 137888 267028
rect 185584 266976 185636 267028
rect 3056 266364 3108 266416
rect 175924 266364 175976 266416
rect 140964 265684 141016 265736
rect 180064 265684 180116 265736
rect 3424 265616 3476 265668
rect 169208 265616 169260 265668
rect 174544 265548 174596 265600
rect 193588 265480 193640 265532
rect 173440 265412 173492 265464
rect 193772 265412 193824 265464
rect 170220 265344 170272 265396
rect 170496 265344 170548 265396
rect 192024 265344 192076 265396
rect 175832 265276 175884 265328
rect 197820 265276 197872 265328
rect 171692 265208 171744 265260
rect 171876 265208 171928 265260
rect 194968 265208 195020 265260
rect 171784 265140 171836 265192
rect 195152 265140 195204 265192
rect 170404 265072 170456 265124
rect 170680 265072 170732 265124
rect 196256 265072 196308 265124
rect 169116 265004 169168 265056
rect 197912 265004 197964 265056
rect 163504 264936 163556 264988
rect 195060 264936 195112 264988
rect 149704 264324 149756 264376
rect 173256 264324 173308 264376
rect 139400 264256 139452 264308
rect 178684 264256 178736 264308
rect 106924 264188 106976 264240
rect 158720 264188 158772 264240
rect 116952 264052 117004 264104
rect 133144 264052 133196 264104
rect 133328 264052 133380 264104
rect 118332 263984 118384 264036
rect 134248 263984 134300 264036
rect 134616 263984 134668 264036
rect 119712 263916 119764 263968
rect 137836 263916 137888 263968
rect 120908 263848 120960 263900
rect 139400 263848 139452 263900
rect 121736 263780 121788 263832
rect 142620 263780 142672 263832
rect 121000 263712 121052 263764
rect 140964 263712 141016 263764
rect 172704 263712 172756 263764
rect 190828 263712 190880 263764
rect 114192 263644 114244 263696
rect 137192 263644 137244 263696
rect 173256 263644 173308 263696
rect 190920 263644 190972 263696
rect 121092 263576 121144 263628
rect 151084 263576 151136 263628
rect 158720 263576 158772 263628
rect 159364 263576 159416 263628
rect 187884 263576 187936 263628
rect 137468 263508 137520 263560
rect 580264 263508 580316 263560
rect 150440 263440 150492 263492
rect 151360 263440 151412 263492
rect 188528 263440 188580 263492
rect 347780 263440 347832 263492
rect 193128 263372 193180 263424
rect 218060 263372 218112 263424
rect 3516 263032 3568 263084
rect 177396 263032 177448 263084
rect 132040 262964 132092 263016
rect 580356 262964 580408 263016
rect 118424 262896 118476 262948
rect 125968 262896 126020 262948
rect 131120 262896 131172 262948
rect 131764 262896 131816 262948
rect 580448 262896 580500 262948
rect 3424 262828 3476 262880
rect 179052 262828 179104 262880
rect 179236 262828 179288 262880
rect 189632 262828 189684 262880
rect 116860 262760 116912 262812
rect 131120 262760 131172 262812
rect 167828 262760 167880 262812
rect 192392 262760 192444 262812
rect 116768 262692 116820 262744
rect 134524 262692 134576 262744
rect 134800 262692 134852 262744
rect 153200 262692 153252 262744
rect 158720 262692 158772 262744
rect 166264 262692 166316 262744
rect 192208 262692 192260 262744
rect 114008 262624 114060 262676
rect 128728 262624 128780 262676
rect 153844 262624 153896 262676
rect 187976 262624 188028 262676
rect 188528 262624 188580 262676
rect 119804 262556 119856 262608
rect 131120 262556 131172 262608
rect 155868 262556 155920 262608
rect 191012 262556 191064 262608
rect 282920 262828 282972 262880
rect 122380 262488 122432 262540
rect 152188 262488 152240 262540
rect 152464 262488 152516 262540
rect 157156 262488 157208 262540
rect 192300 262488 192352 262540
rect 193128 262488 193180 262540
rect 118056 262420 118108 262472
rect 129280 262420 129332 262472
rect 181444 262420 181496 262472
rect 192116 262420 192168 262472
rect 119620 262352 119672 262404
rect 127716 262352 127768 262404
rect 184756 262352 184808 262404
rect 193680 262352 193732 262404
rect 113916 262284 113968 262336
rect 127072 262284 127124 262336
rect 182916 262284 182968 262336
rect 190460 262284 190512 262336
rect 181168 262216 181220 262268
rect 187700 262216 187752 262268
rect 129832 261400 129884 261452
rect 188344 261400 188396 261452
rect 179052 261332 179104 261384
rect 198096 261332 198148 261384
rect 131120 261264 131172 261316
rect 471244 261264 471296 261316
rect 177948 261196 178000 261248
rect 191288 261196 191340 261248
rect 180708 261128 180760 261180
rect 196716 261128 196768 261180
rect 120816 261060 120868 261112
rect 133236 261060 133288 261112
rect 177396 261060 177448 261112
rect 196532 261060 196584 261112
rect 115296 260992 115348 261044
rect 130384 260992 130436 261044
rect 181996 260992 182048 261044
rect 196440 260992 196492 261044
rect 14464 260924 14516 260976
rect 176200 260924 176252 260976
rect 189724 260924 189776 260976
rect 115572 260856 115624 260908
rect 132040 260856 132092 260908
rect 184020 260856 184072 260908
rect 198004 260856 198056 260908
rect 118240 260788 118292 260840
rect 124312 260788 124364 260840
rect 181260 260516 181312 260568
rect 188068 260516 188120 260568
rect 179696 260448 179748 260500
rect 192300 260448 192352 260500
rect 4804 260380 4856 260432
rect 177948 260380 178000 260432
rect 178684 260380 178736 260432
rect 191104 260380 191156 260432
rect 133236 260312 133288 260364
rect 169208 260244 169260 260296
rect 178684 260244 178736 260296
rect 472624 260312 472676 260364
rect 122196 260108 122248 260160
rect 135260 260176 135312 260228
rect 136226 260176 136278 260228
rect 157340 260176 157392 260228
rect 158306 260176 158358 260228
rect 167000 260176 167052 260228
rect 167690 260176 167742 260228
rect 169760 260176 169812 260228
rect 171002 260176 171054 260228
rect 189356 260176 189408 260228
rect 175924 260108 175976 260160
rect 189540 260108 189592 260160
rect 115480 260040 115532 260092
rect 126842 260040 126894 260092
rect 167690 260040 167742 260092
rect 118148 259972 118200 260024
rect 139676 259972 139728 260024
rect 189448 260040 189500 260092
rect 178500 259972 178552 260024
rect 181628 259972 181680 260024
rect 181720 259972 181772 260024
rect 184664 259972 184716 260024
rect 119528 259904 119580 259956
rect 140780 259904 140832 259956
rect 141424 259904 141476 259956
rect 164700 259904 164752 259956
rect 187976 259972 188028 260024
rect 121920 259836 121972 259888
rect 146300 259836 146352 259888
rect 166172 259836 166224 259888
rect 191196 259836 191248 259888
rect 121184 259768 121236 259820
rect 147680 259768 147732 259820
rect 158076 259768 158128 259820
rect 181260 259768 181312 259820
rect 181628 259768 181680 259820
rect 188252 259768 188304 259820
rect 119436 259700 119488 259752
rect 153200 259700 153252 259752
rect 158628 259700 158680 259752
rect 179696 259700 179748 259752
rect 180156 259700 180208 259752
rect 134340 259632 134392 259684
rect 120632 259564 120684 259616
rect 178040 259564 178092 259616
rect 120724 259496 120776 259548
rect 125600 259496 125652 259548
rect 174452 259496 174504 259548
rect 181720 259564 181772 259616
rect 116676 259428 116728 259480
rect 128360 259428 128412 259480
rect 184572 259700 184624 259752
rect 190552 259700 190604 259752
rect 184664 259632 184716 259684
rect 187332 259632 187384 259684
rect 187240 259564 187292 259616
rect 183468 259496 183520 259548
rect 195244 259496 195296 259548
rect 580172 259360 580224 259412
rect 472624 245556 472676 245608
rect 580172 245556 580224 245608
rect 3516 241408 3568 241460
rect 14464 241408 14516 241460
rect 2780 215228 2832 215280
rect 4804 215228 4856 215280
rect 471244 206932 471296 206984
rect 579804 206932 579856 206984
rect 111708 200608 111760 200660
rect 131948 200608 132000 200660
rect 115848 200540 115900 200592
rect 122748 200472 122800 200524
rect 112996 200404 113048 200456
rect 132040 200404 132092 200456
rect 107200 200336 107252 200388
rect 113088 200268 113140 200320
rect 130936 200268 130988 200320
rect 122564 200132 122616 200184
rect 125600 200064 125652 200116
rect 125232 199928 125284 199980
rect 127532 199860 127584 199912
rect 132914 199860 132966 199912
rect 133098 199860 133150 199912
rect 133190 199860 133242 199912
rect 133466 199860 133518 199912
rect 133742 199860 133794 199912
rect 134018 199860 134070 199912
rect 134110 199860 134162 199912
rect 134478 199860 134530 199912
rect 134570 199860 134622 199912
rect 134662 199860 134714 199912
rect 135214 199860 135266 199912
rect 135490 199860 135542 199912
rect 135674 199860 135726 199912
rect 136042 199860 136094 199912
rect 136318 199860 136370 199912
rect 136502 199860 136554 199912
rect 136686 199860 136738 199912
rect 136870 199860 136922 199912
rect 132868 199724 132920 199776
rect 111248 199656 111300 199708
rect 128820 199656 128872 199708
rect 133282 199792 133334 199844
rect 133328 199656 133380 199708
rect 133420 199656 133472 199708
rect 111524 199588 111576 199640
rect 131580 199588 131632 199640
rect 133144 199588 133196 199640
rect 134064 199588 134116 199640
rect 134524 199724 134576 199776
rect 134616 199724 134668 199776
rect 135536 199724 135588 199776
rect 135628 199656 135680 199708
rect 134708 199588 134760 199640
rect 135352 199588 135404 199640
rect 136180 199588 136232 199640
rect 136732 199724 136784 199776
rect 136824 199724 136876 199776
rect 137054 199860 137106 199912
rect 137422 199860 137474 199912
rect 137790 199860 137842 199912
rect 138250 199860 138302 199912
rect 138342 199860 138394 199912
rect 138526 199860 138578 199912
rect 138802 199860 138854 199912
rect 137238 199792 137290 199844
rect 137100 199656 137152 199708
rect 137192 199656 137244 199708
rect 136456 199588 136508 199640
rect 136548 199588 136600 199640
rect 137836 199724 137888 199776
rect 138204 199724 138256 199776
rect 138204 199588 138256 199640
rect 138480 199588 138532 199640
rect 138664 199588 138716 199640
rect 139078 199860 139130 199912
rect 139170 199860 139222 199912
rect 139262 199860 139314 199912
rect 139354 199860 139406 199912
rect 139906 199860 139958 199912
rect 140090 199860 140142 199912
rect 140274 199860 140326 199912
rect 140458 199860 140510 199912
rect 140826 199860 140878 199912
rect 140918 199860 140970 199912
rect 141010 199860 141062 199912
rect 141102 199860 141154 199912
rect 141194 199860 141246 199912
rect 141286 199860 141338 199912
rect 141378 199860 141430 199912
rect 141562 199860 141614 199912
rect 141654 199860 141706 199912
rect 141746 199860 141798 199912
rect 141838 199860 141890 199912
rect 138940 199588 138992 199640
rect 139124 199724 139176 199776
rect 139216 199656 139268 199708
rect 139308 199588 139360 199640
rect 139952 199588 140004 199640
rect 140366 199792 140418 199844
rect 140642 199792 140694 199844
rect 140734 199792 140786 199844
rect 140320 199656 140372 199708
rect 140412 199656 140464 199708
rect 140918 199724 140970 199776
rect 141102 199656 141154 199708
rect 141240 199656 141292 199708
rect 140228 199588 140280 199640
rect 140596 199588 140648 199640
rect 140688 199588 140740 199640
rect 140780 199588 140832 199640
rect 141010 199588 141062 199640
rect 141424 199588 141476 199640
rect 141608 199724 141660 199776
rect 141700 199724 141752 199776
rect 141792 199656 141844 199708
rect 142390 199860 142442 199912
rect 142574 199860 142626 199912
rect 142666 199860 142718 199912
rect 142758 199860 142810 199912
rect 142942 199860 142994 199912
rect 143310 199860 143362 199912
rect 143402 199860 143454 199912
rect 143862 199860 143914 199912
rect 143954 199860 144006 199912
rect 144598 199860 144650 199912
rect 144690 199860 144742 199912
rect 144966 199860 145018 199912
rect 145242 199860 145294 199912
rect 145334 199860 145386 199912
rect 145426 199860 145478 199912
rect 145610 199860 145662 199912
rect 146070 199860 146122 199912
rect 146162 199860 146214 199912
rect 142436 199724 142488 199776
rect 142712 199724 142764 199776
rect 142528 199656 142580 199708
rect 142620 199656 142672 199708
rect 143356 199656 143408 199708
rect 143448 199656 143500 199708
rect 141976 199588 142028 199640
rect 142252 199588 142304 199640
rect 142896 199588 142948 199640
rect 144092 199656 144144 199708
rect 143908 199588 143960 199640
rect 144000 199588 144052 199640
rect 115664 199520 115716 199572
rect 143632 199520 143684 199572
rect 144092 199520 144144 199572
rect 144644 199724 144696 199776
rect 144920 199656 144972 199708
rect 145380 199724 145432 199776
rect 145288 199656 145340 199708
rect 144368 199588 144420 199640
rect 145564 199724 145616 199776
rect 146116 199724 146168 199776
rect 146024 199588 146076 199640
rect 146438 199860 146490 199912
rect 146622 199860 146674 199912
rect 146898 199860 146950 199912
rect 147082 199860 147134 199912
rect 147174 199860 147226 199912
rect 147358 199860 147410 199912
rect 147634 199860 147686 199912
rect 147818 199860 147870 199912
rect 148094 199860 148146 199912
rect 148278 199860 148330 199912
rect 148462 199860 148514 199912
rect 148738 199860 148790 199912
rect 148830 199860 148882 199912
rect 148922 199860 148974 199912
rect 149106 199860 149158 199912
rect 149382 199860 149434 199912
rect 144828 199520 144880 199572
rect 145104 199520 145156 199572
rect 146576 199588 146628 199640
rect 146944 199588 146996 199640
rect 147036 199588 147088 199640
rect 147312 199588 147364 199640
rect 112812 199452 112864 199504
rect 148048 199724 148100 199776
rect 148692 199724 148744 199776
rect 148784 199724 148836 199776
rect 149566 199860 149618 199912
rect 149612 199724 149664 199776
rect 147772 199588 147824 199640
rect 148232 199588 148284 199640
rect 148416 199588 148468 199640
rect 148876 199588 148928 199640
rect 147588 199520 147640 199572
rect 149842 199860 149894 199912
rect 149934 199860 149986 199912
rect 150118 199860 150170 199912
rect 150302 199860 150354 199912
rect 150394 199860 150446 199912
rect 149888 199724 149940 199776
rect 150072 199724 150124 199776
rect 150348 199656 150400 199708
rect 150256 199588 150308 199640
rect 150072 199520 150124 199572
rect 150670 199860 150722 199912
rect 150762 199860 150814 199912
rect 150854 199860 150906 199912
rect 150946 199860 150998 199912
rect 151222 199860 151274 199912
rect 151314 199860 151366 199912
rect 151406 199860 151458 199912
rect 149244 199452 149296 199504
rect 150716 199724 150768 199776
rect 151176 199656 151228 199708
rect 151084 199588 151136 199640
rect 151544 199588 151596 199640
rect 151360 199520 151412 199572
rect 151268 199452 151320 199504
rect 177856 200608 177908 200660
rect 180064 200608 180116 200660
rect 183836 200540 183888 200592
rect 186872 200540 186924 200592
rect 151774 199860 151826 199912
rect 151866 199860 151918 199912
rect 151958 199860 152010 199912
rect 152142 199860 152194 199912
rect 153062 199860 153114 199912
rect 153246 199860 153298 199912
rect 153338 199860 153390 199912
rect 153522 199860 153574 199912
rect 153706 199860 153758 199912
rect 153798 199860 153850 199912
rect 154074 199860 154126 199912
rect 154258 199860 154310 199912
rect 154534 199860 154586 199912
rect 154718 199860 154770 199912
rect 154994 199860 155046 199912
rect 155086 199860 155138 199912
rect 155178 199860 155230 199912
rect 155362 199860 155414 199912
rect 155454 199860 155506 199912
rect 155822 199860 155874 199912
rect 156098 199860 156150 199912
rect 156466 199860 156518 199912
rect 156650 199860 156702 199912
rect 156742 199860 156794 199912
rect 156926 199860 156978 199912
rect 157110 199860 157162 199912
rect 157294 199860 157346 199912
rect 157386 199860 157438 199912
rect 157662 199860 157714 199912
rect 157938 199860 157990 199912
rect 158214 199860 158266 199912
rect 158490 199860 158542 199912
rect 158766 199860 158818 199912
rect 158950 199860 159002 199912
rect 159226 199860 159278 199912
rect 159318 199860 159370 199912
rect 159502 199860 159554 199912
rect 159870 199860 159922 199912
rect 151820 199724 151872 199776
rect 151912 199656 151964 199708
rect 152004 199588 152056 199640
rect 152694 199792 152746 199844
rect 152786 199792 152838 199844
rect 152970 199792 153022 199844
rect 152464 199520 152516 199572
rect 152648 199520 152700 199572
rect 152924 199588 152976 199640
rect 119896 199384 119948 199436
rect 145656 199384 145708 199436
rect 146852 199384 146904 199436
rect 121184 199316 121236 199368
rect 148140 199316 148192 199368
rect 117228 199248 117280 199300
rect 145196 199248 145248 199300
rect 108856 199180 108908 199232
rect 131488 199180 131540 199232
rect 131580 199180 131632 199232
rect 136824 199180 136876 199232
rect 138848 199180 138900 199232
rect 139032 199180 139084 199232
rect 114376 199112 114428 199164
rect 145932 199180 145984 199232
rect 151452 199384 151504 199436
rect 151820 199384 151872 199436
rect 152280 199452 152332 199504
rect 153200 199520 153252 199572
rect 153752 199656 153804 199708
rect 153476 199588 153528 199640
rect 153660 199588 153712 199640
rect 153936 199588 153988 199640
rect 153844 199520 153896 199572
rect 153936 199452 153988 199504
rect 154028 199452 154080 199504
rect 154304 199724 154356 199776
rect 154764 199656 154816 199708
rect 154672 199520 154724 199572
rect 155224 199724 155276 199776
rect 155408 199724 155460 199776
rect 156282 199792 156334 199844
rect 155776 199588 155828 199640
rect 155960 199588 156012 199640
rect 156144 199588 156196 199640
rect 156236 199588 156288 199640
rect 155316 199520 155368 199572
rect 155868 199520 155920 199572
rect 156420 199656 156472 199708
rect 156604 199588 156656 199640
rect 156880 199724 156932 199776
rect 157340 199656 157392 199708
rect 157248 199588 157300 199640
rect 156696 199520 156748 199572
rect 157064 199520 157116 199572
rect 155040 199452 155092 199504
rect 155592 199452 155644 199504
rect 158260 199588 158312 199640
rect 158444 199588 158496 199640
rect 158628 199520 158680 199572
rect 158996 199724 159048 199776
rect 159272 199724 159324 199776
rect 159180 199588 159232 199640
rect 159548 199588 159600 199640
rect 153016 199384 153068 199436
rect 153292 199384 153344 199436
rect 158812 199452 158864 199504
rect 159824 199588 159876 199640
rect 160146 199860 160198 199912
rect 160330 199860 160382 199912
rect 160514 199860 160566 199912
rect 160698 199860 160750 199912
rect 160790 199860 160842 199912
rect 161158 199860 161210 199912
rect 161434 199860 161486 199912
rect 160192 199588 160244 199640
rect 160376 199588 160428 199640
rect 160468 199588 160520 199640
rect 160744 199656 160796 199708
rect 160928 199588 160980 199640
rect 161710 199860 161762 199912
rect 161894 199860 161946 199912
rect 162170 199860 162222 199912
rect 162262 199860 162314 199912
rect 162354 199860 162406 199912
rect 162446 199860 162498 199912
rect 161572 199588 161624 199640
rect 160652 199520 160704 199572
rect 161664 199520 161716 199572
rect 159916 199452 159968 199504
rect 156144 199384 156196 199436
rect 161204 199384 161256 199436
rect 150808 199316 150860 199368
rect 155960 199316 156012 199368
rect 159364 199316 159416 199368
rect 162078 199724 162130 199776
rect 162032 199520 162084 199572
rect 162308 199724 162360 199776
rect 162630 199860 162682 199912
rect 162584 199588 162636 199640
rect 163044 199588 163096 199640
rect 197360 200472 197412 200524
rect 198832 200404 198884 200456
rect 178868 200336 178920 200388
rect 193312 200268 193364 200320
rect 178040 200200 178092 200252
rect 193496 200200 193548 200252
rect 163918 199860 163970 199912
rect 164562 199860 164614 199912
rect 164654 199860 164706 199912
rect 164746 199860 164798 199912
rect 163780 199588 163832 199640
rect 164516 199588 164568 199640
rect 164930 199860 164982 199912
rect 165022 199860 165074 199912
rect 165114 199860 165166 199912
rect 165298 199860 165350 199912
rect 165390 199860 165442 199912
rect 165482 199860 165534 199912
rect 165574 199860 165626 199912
rect 165666 199860 165718 199912
rect 165758 199860 165810 199912
rect 164792 199656 164844 199708
rect 164700 199588 164752 199640
rect 165436 199724 165488 199776
rect 166034 199792 166086 199844
rect 164976 199656 165028 199708
rect 165068 199656 165120 199708
rect 165344 199656 165396 199708
rect 165528 199656 165580 199708
rect 165712 199656 165764 199708
rect 165160 199588 165212 199640
rect 165988 199588 166040 199640
rect 162492 199520 162544 199572
rect 166218 199860 166270 199912
rect 166770 199860 166822 199912
rect 166862 199860 166914 199912
rect 167046 199860 167098 199912
rect 167138 199860 167190 199912
rect 167230 199860 167282 199912
rect 167414 199860 167466 199912
rect 166310 199792 166362 199844
rect 166724 199724 166776 199776
rect 166908 199724 166960 199776
rect 166816 199656 166868 199708
rect 166816 199520 166868 199572
rect 162216 199452 162268 199504
rect 162768 199452 162820 199504
rect 164240 199452 164292 199504
rect 166172 199452 166224 199504
rect 167184 199656 167236 199708
rect 167368 199588 167420 199640
rect 167000 199520 167052 199572
rect 165252 199384 165304 199436
rect 165620 199384 165672 199436
rect 162768 199316 162820 199368
rect 167874 199860 167926 199912
rect 167966 199860 168018 199912
rect 168058 199860 168110 199912
rect 168426 199860 168478 199912
rect 168794 199860 168846 199912
rect 168886 199860 168938 199912
rect 168978 199860 169030 199912
rect 169254 199860 169306 199912
rect 167920 199724 167972 199776
rect 168012 199656 168064 199708
rect 168472 199588 168524 199640
rect 168840 199656 168892 199708
rect 168932 199656 168984 199708
rect 169392 199588 169444 199640
rect 169208 199520 169260 199572
rect 169622 199860 169674 199912
rect 169714 199860 169766 199912
rect 169806 199860 169858 199912
rect 169898 199860 169950 199912
rect 170082 199860 170134 199912
rect 170174 199860 170226 199912
rect 170542 199860 170594 199912
rect 170634 199860 170686 199912
rect 170726 199860 170778 199912
rect 170818 199860 170870 199912
rect 169576 199656 169628 199708
rect 169668 199656 169720 199708
rect 169576 199520 169628 199572
rect 168656 199452 168708 199504
rect 167736 199316 167788 199368
rect 170036 199724 170088 199776
rect 169852 199656 169904 199708
rect 170496 199724 170548 199776
rect 170588 199656 170640 199708
rect 170128 199588 170180 199640
rect 186780 200132 186832 200184
rect 186872 200132 186924 200184
rect 190552 200132 190604 200184
rect 181904 200064 181956 200116
rect 171094 199860 171146 199912
rect 171048 199724 171100 199776
rect 170864 199520 170916 199572
rect 171278 199860 171330 199912
rect 171830 199860 171882 199912
rect 171922 199860 171974 199912
rect 172198 199860 172250 199912
rect 172566 199860 172618 199912
rect 172750 199860 172802 199912
rect 173118 199860 173170 199912
rect 171876 199656 171928 199708
rect 171324 199588 171376 199640
rect 172060 199588 172112 199640
rect 172244 199588 172296 199640
rect 172152 199520 172204 199572
rect 172336 199520 172388 199572
rect 172428 199520 172480 199572
rect 172796 199520 172848 199572
rect 169760 199452 169812 199504
rect 170772 199452 170824 199504
rect 171600 199452 171652 199504
rect 171968 199452 172020 199504
rect 151084 199248 151136 199300
rect 157156 199248 157208 199300
rect 160560 199248 160612 199300
rect 161848 199248 161900 199300
rect 164884 199248 164936 199300
rect 169760 199316 169812 199368
rect 171968 199316 172020 199368
rect 173578 199860 173630 199912
rect 173532 199520 173584 199572
rect 174038 199860 174090 199912
rect 174130 199860 174182 199912
rect 174222 199860 174274 199912
rect 174406 199860 174458 199912
rect 174498 199860 174550 199912
rect 174084 199724 174136 199776
rect 174268 199520 174320 199572
rect 173348 199452 173400 199504
rect 174176 199452 174228 199504
rect 174452 199656 174504 199708
rect 174682 199860 174734 199912
rect 174774 199860 174826 199912
rect 174958 199860 175010 199912
rect 174820 199588 174872 199640
rect 175004 199588 175056 199640
rect 174728 199520 174780 199572
rect 187516 199996 187568 200048
rect 175510 199860 175562 199912
rect 175602 199860 175654 199912
rect 175970 199860 176022 199912
rect 176062 199860 176114 199912
rect 176154 199860 176206 199912
rect 176246 199860 176298 199912
rect 176706 199860 176758 199912
rect 176798 199860 176850 199912
rect 176982 199860 177034 199912
rect 177258 199860 177310 199912
rect 177672 199860 177724 199912
rect 175924 199724 175976 199776
rect 176108 199724 176160 199776
rect 175556 199656 175608 199708
rect 195520 199792 195572 199844
rect 176844 199724 176896 199776
rect 176936 199724 176988 199776
rect 177166 199724 177218 199776
rect 199568 199724 199620 199776
rect 176016 199588 176068 199640
rect 176200 199588 176252 199640
rect 177396 199520 177448 199572
rect 177672 199520 177724 199572
rect 177948 199520 178000 199572
rect 178224 199520 178276 199572
rect 186596 199520 186648 199572
rect 175188 199452 175240 199504
rect 175924 199452 175976 199504
rect 176384 199452 176436 199504
rect 177580 199452 177632 199504
rect 178132 199452 178184 199504
rect 173808 199384 173860 199436
rect 180340 199384 180392 199436
rect 182824 199384 182876 199436
rect 190460 199384 190512 199436
rect 156144 199180 156196 199232
rect 159732 199180 159784 199232
rect 143632 199112 143684 199164
rect 148416 199112 148468 199164
rect 152832 199112 152884 199164
rect 115756 199044 115808 199096
rect 147588 199044 147640 199096
rect 159456 199044 159508 199096
rect 160008 199044 160060 199096
rect 162400 199112 162452 199164
rect 165712 199112 165764 199164
rect 164884 199044 164936 199096
rect 178040 199248 178092 199300
rect 169392 199180 169444 199232
rect 171140 199112 171192 199164
rect 172336 199180 172388 199232
rect 173716 199180 173768 199232
rect 203064 199316 203116 199368
rect 175188 199112 175240 199164
rect 201040 199112 201092 199164
rect 169392 199044 169444 199096
rect 169944 199044 169996 199096
rect 170772 199044 170824 199096
rect 175740 199044 175792 199096
rect 186412 199044 186464 199096
rect 187516 199044 187568 199096
rect 198740 199044 198792 199096
rect 133144 198976 133196 199028
rect 159824 198976 159876 199028
rect 166356 198976 166408 199028
rect 200212 198976 200264 199028
rect 114468 198908 114520 198960
rect 147036 198908 147088 198960
rect 159640 198908 159692 198960
rect 160008 198908 160060 198960
rect 169392 198908 169444 198960
rect 170772 198908 170824 198960
rect 174268 198908 174320 198960
rect 178776 198908 178828 198960
rect 181076 198908 181128 198960
rect 187700 198908 187752 198960
rect 121368 198840 121420 198892
rect 140320 198840 140372 198892
rect 159180 198840 159232 198892
rect 162768 198840 162820 198892
rect 167460 198840 167512 198892
rect 201868 198840 201920 198892
rect 126336 198772 126388 198824
rect 147680 198772 147732 198824
rect 150256 198772 150308 198824
rect 157432 198772 157484 198824
rect 158996 198772 159048 198824
rect 167736 198772 167788 198824
rect 167828 198772 167880 198824
rect 170128 198772 170180 198824
rect 171140 198772 171192 198824
rect 174268 198772 174320 198824
rect 118608 198704 118660 198756
rect 144368 198704 144420 198756
rect 170772 198704 170824 198756
rect 180156 198772 180208 198824
rect 186412 198772 186464 198824
rect 200948 198772 201000 198824
rect 174820 198704 174872 198756
rect 200580 198704 200632 198756
rect 130936 198636 130988 198688
rect 144828 198636 144880 198688
rect 173072 198636 173124 198688
rect 195980 198636 196032 198688
rect 126704 198568 126756 198620
rect 146668 198568 146720 198620
rect 167092 198568 167144 198620
rect 178684 198568 178736 198620
rect 181904 198568 181956 198620
rect 194048 198568 194100 198620
rect 108672 198500 108724 198552
rect 133328 198500 133380 198552
rect 157892 198500 157944 198552
rect 171784 198500 171836 198552
rect 123300 198432 123352 198484
rect 143724 198432 143776 198484
rect 156696 198432 156748 198484
rect 171508 198432 171560 198484
rect 173256 198432 173308 198484
rect 199108 198432 199160 198484
rect 108396 198364 108448 198416
rect 132500 198364 132552 198416
rect 159824 198364 159876 198416
rect 171324 198364 171376 198416
rect 177396 198364 177448 198416
rect 197728 198364 197780 198416
rect 122472 198296 122524 198348
rect 148232 198296 148284 198348
rect 169944 198296 169996 198348
rect 196624 198296 196676 198348
rect 106924 198228 106976 198280
rect 127532 198228 127584 198280
rect 136548 198228 136600 198280
rect 138020 198228 138072 198280
rect 172520 198228 172572 198280
rect 198188 198228 198240 198280
rect 122288 198160 122340 198212
rect 149152 198160 149204 198212
rect 156420 198160 156472 198212
rect 171324 198160 171376 198212
rect 172152 198160 172204 198212
rect 181444 198160 181496 198212
rect 199568 198160 199620 198212
rect 204720 198160 204772 198212
rect 103336 198092 103388 198144
rect 134892 198092 134944 198144
rect 153384 198092 153436 198144
rect 171140 198092 171192 198144
rect 173900 198092 173952 198144
rect 200396 198092 200448 198144
rect 103428 198024 103480 198076
rect 133604 198024 133656 198076
rect 173348 198024 173400 198076
rect 200672 198024 200724 198076
rect 102876 197956 102928 198008
rect 125600 197956 125652 198008
rect 157616 197956 157668 198008
rect 169760 197956 169812 198008
rect 172244 197956 172296 198008
rect 199384 197956 199436 198008
rect 132224 197820 132276 197872
rect 151176 197888 151228 197940
rect 163320 197888 163372 197940
rect 163504 197888 163556 197940
rect 138296 197820 138348 197872
rect 149428 197820 149480 197872
rect 155040 197820 155092 197872
rect 171876 197888 171928 197940
rect 173532 197888 173584 197940
rect 193864 197888 193916 197940
rect 170496 197820 170548 197872
rect 187700 197820 187752 197872
rect 126152 197752 126204 197804
rect 144828 197752 144880 197804
rect 170220 197752 170272 197804
rect 186688 197752 186740 197804
rect 163780 197684 163832 197736
rect 189080 197684 189132 197736
rect 131028 197616 131080 197668
rect 138296 197616 138348 197668
rect 171784 197616 171836 197668
rect 180432 197616 180484 197668
rect 165620 197548 165672 197600
rect 181628 197548 181680 197600
rect 145472 197480 145524 197532
rect 147680 197480 147732 197532
rect 171324 197480 171376 197532
rect 172428 197480 172480 197532
rect 120448 197412 120500 197464
rect 144184 197412 144236 197464
rect 171508 197412 171560 197464
rect 172152 197412 172204 197464
rect 117320 197344 117372 197396
rect 138940 197344 138992 197396
rect 174084 197344 174136 197396
rect 174452 197344 174504 197396
rect 130568 197276 130620 197328
rect 150532 197276 150584 197328
rect 164792 197276 164844 197328
rect 199016 197276 199068 197328
rect 112904 197208 112956 197260
rect 117136 197140 117188 197192
rect 120448 197140 120500 197192
rect 132960 197140 133012 197192
rect 140044 197140 140096 197192
rect 164148 197208 164200 197260
rect 193220 197208 193272 197260
rect 142896 197140 142948 197192
rect 164424 197140 164476 197192
rect 199660 197140 199712 197192
rect 111616 197072 111668 197124
rect 143264 197072 143316 197124
rect 147588 197072 147640 197124
rect 154856 197072 154908 197124
rect 163504 197072 163556 197124
rect 197452 197072 197504 197124
rect 117044 197004 117096 197056
rect 148600 197004 148652 197056
rect 160836 197004 160888 197056
rect 194692 197004 194744 197056
rect 112720 196936 112772 196988
rect 132776 196936 132828 196988
rect 133144 196936 133196 196988
rect 142528 196936 142580 196988
rect 163688 196936 163740 196988
rect 197544 196936 197596 196988
rect 110328 196868 110380 196920
rect 142804 196868 142856 196920
rect 160376 196868 160428 196920
rect 194876 196868 194928 196920
rect 111340 196800 111392 196852
rect 132960 196800 133012 196852
rect 106832 196732 106884 196784
rect 140136 196800 140188 196852
rect 177856 196800 177908 196852
rect 196348 196800 196400 196852
rect 140044 196732 140096 196784
rect 143724 196732 143776 196784
rect 158996 196732 159048 196784
rect 187792 196732 187844 196784
rect 109776 196664 109828 196716
rect 133144 196664 133196 196716
rect 171784 196664 171836 196716
rect 197636 196664 197688 196716
rect 106096 196596 106148 196648
rect 139584 196596 139636 196648
rect 159548 196596 159600 196648
rect 193404 196596 193456 196648
rect 123392 196460 123444 196512
rect 133328 196460 133380 196512
rect 144092 196460 144144 196512
rect 162308 196460 162360 196512
rect 180248 196528 180300 196580
rect 143448 196392 143500 196444
rect 132776 196256 132828 196308
rect 133328 196256 133380 196308
rect 147956 196188 148008 196240
rect 157892 196188 157944 196240
rect 165620 196188 165672 196240
rect 166172 196188 166224 196240
rect 134156 196052 134208 196104
rect 134708 196052 134760 196104
rect 133696 195984 133748 196036
rect 135996 195984 136048 196036
rect 122656 195916 122708 195968
rect 154304 195916 154356 195968
rect 172152 195916 172204 195968
rect 190644 195916 190696 195968
rect 111432 195848 111484 195900
rect 133696 195848 133748 195900
rect 114100 195780 114152 195832
rect 152004 195848 152056 195900
rect 152648 195848 152700 195900
rect 172428 195848 172480 195900
rect 190736 195848 190788 195900
rect 145012 195780 145064 195832
rect 156972 195780 157024 195832
rect 166264 195780 166316 195832
rect 169760 195780 169812 195832
rect 192576 195780 192628 195832
rect 103060 195712 103112 195764
rect 134340 195712 134392 195764
rect 135996 195712 136048 195764
rect 142436 195712 142488 195764
rect 158076 195712 158128 195764
rect 191840 195712 191892 195764
rect 107016 195644 107068 195696
rect 137928 195644 137980 195696
rect 165712 195644 165764 195696
rect 196072 195644 196124 195696
rect 110236 195576 110288 195628
rect 143080 195576 143132 195628
rect 161572 195576 161624 195628
rect 194600 195576 194652 195628
rect 114284 195508 114336 195560
rect 147128 195508 147180 195560
rect 166264 195508 166316 195560
rect 190460 195508 190512 195560
rect 118884 195440 118936 195492
rect 153108 195440 153160 195492
rect 162216 195440 162268 195492
rect 196164 195440 196216 195492
rect 105636 195372 105688 195424
rect 117320 195372 117372 195424
rect 138664 195372 138716 195424
rect 140780 195372 140832 195424
rect 157340 195372 157392 195424
rect 190552 195372 190604 195424
rect 105820 195304 105872 195356
rect 139860 195304 139912 195356
rect 158720 195304 158772 195356
rect 191932 195304 191984 195356
rect 112628 195236 112680 195288
rect 145104 195236 145156 195288
rect 157248 195236 157300 195288
rect 157800 195236 157852 195288
rect 161848 195236 161900 195288
rect 194784 195236 194836 195288
rect 118516 195168 118568 195220
rect 148968 195168 149020 195220
rect 164976 195168 165028 195220
rect 165160 195168 165212 195220
rect 169024 195168 169076 195220
rect 169576 195168 169628 195220
rect 148232 195100 148284 195152
rect 148784 195100 148836 195152
rect 168748 195100 168800 195152
rect 169208 195100 169260 195152
rect 171876 194896 171928 194948
rect 189172 195168 189224 195220
rect 171140 194828 171192 194880
rect 188160 195100 188212 195152
rect 124864 194760 124916 194812
rect 137652 194760 137704 194812
rect 167000 194624 167052 194676
rect 184204 194624 184256 194676
rect 122104 194488 122156 194540
rect 149428 194488 149480 194540
rect 167000 194488 167052 194540
rect 168656 194488 168708 194540
rect 104164 194420 104216 194472
rect 132592 194420 132644 194472
rect 111064 194352 111116 194404
rect 141792 194352 141844 194404
rect 166080 194352 166132 194404
rect 182916 194352 182968 194404
rect 108764 194284 108816 194336
rect 136916 194284 136968 194336
rect 138756 194284 138808 194336
rect 138940 194284 138992 194336
rect 104716 194216 104768 194268
rect 136364 194216 136416 194268
rect 161480 194216 161532 194268
rect 161756 194216 161808 194268
rect 168012 194216 168064 194268
rect 201592 194216 201644 194268
rect 104348 194148 104400 194200
rect 135720 194148 135772 194200
rect 168564 194148 168616 194200
rect 203340 194148 203392 194200
rect 104532 194080 104584 194132
rect 136088 194080 136140 194132
rect 169116 194080 169168 194132
rect 203248 194080 203300 194132
rect 100576 194012 100628 194064
rect 125232 194012 125284 194064
rect 167184 194012 167236 194064
rect 202052 194012 202104 194064
rect 101680 193944 101732 193996
rect 134064 193944 134116 193996
rect 153936 193944 153988 193996
rect 205824 193944 205876 193996
rect 103152 193876 103204 193928
rect 135536 193876 135588 193928
rect 161848 193876 161900 193928
rect 205732 193876 205784 193928
rect 105912 193808 105964 193860
rect 140504 193808 140556 193860
rect 151268 193808 151320 193860
rect 206100 193808 206152 193860
rect 112536 193740 112588 193792
rect 117688 193740 117740 193792
rect 122012 193672 122064 193724
rect 147956 193672 148008 193724
rect 123208 193604 123260 193656
rect 146024 193604 146076 193656
rect 176016 193536 176068 193588
rect 188712 193536 188764 193588
rect 105728 193128 105780 193180
rect 137008 193128 137060 193180
rect 156328 193128 156380 193180
rect 183100 193128 183152 193180
rect 188344 193128 188396 193180
rect 580172 193128 580224 193180
rect 108304 193060 108356 193112
rect 140688 193060 140740 193112
rect 176844 193060 176896 193112
rect 204352 193060 204404 193112
rect 110144 192992 110196 193044
rect 144736 192992 144788 193044
rect 165528 192992 165580 193044
rect 192484 192992 192536 193044
rect 111156 192924 111208 192976
rect 144368 192924 144420 192976
rect 153384 192924 153436 192976
rect 154028 192924 154080 192976
rect 170128 192924 170180 192976
rect 201776 192924 201828 192976
rect 110052 192856 110104 192908
rect 144000 192856 144052 192908
rect 167276 192856 167328 192908
rect 168288 192856 168340 192908
rect 174452 192856 174504 192908
rect 205916 192856 205968 192908
rect 106004 192788 106056 192840
rect 131580 192788 131632 192840
rect 163044 192788 163096 192840
rect 163412 192788 163464 192840
rect 172704 192788 172756 192840
rect 206008 192788 206060 192840
rect 115388 192720 115440 192772
rect 149796 192720 149848 192772
rect 164240 192720 164292 192772
rect 195980 192720 196032 192772
rect 104256 192652 104308 192704
rect 136548 192652 136600 192704
rect 169484 192652 169536 192704
rect 202880 192652 202932 192704
rect 109868 192584 109920 192636
rect 144552 192584 144604 192636
rect 168196 192584 168248 192636
rect 201684 192584 201736 192636
rect 102784 192516 102836 192568
rect 136824 192516 136876 192568
rect 178684 192516 178736 192568
rect 200304 192516 200356 192568
rect 108580 192448 108632 192500
rect 141976 192448 142028 192500
rect 166816 192448 166868 192500
rect 200764 192448 200816 192500
rect 107476 192380 107528 192432
rect 137744 192380 137796 192432
rect 156236 192380 156288 192432
rect 181536 192380 181588 192432
rect 157524 192312 157576 192364
rect 181444 192312 181496 192364
rect 157432 192244 157484 192296
rect 158260 192244 158312 192296
rect 165804 192244 165856 192296
rect 166724 192244 166776 192296
rect 158996 191224 159048 191276
rect 159916 191224 159968 191276
rect 164332 191224 164384 191276
rect 164608 191224 164660 191276
rect 167092 191224 167144 191276
rect 168104 191224 168156 191276
rect 150532 191156 150584 191208
rect 151820 191156 151872 191208
rect 173992 191156 174044 191208
rect 175004 191156 175056 191208
rect 146760 191088 146812 191140
rect 147312 191088 147364 191140
rect 151728 191088 151780 191140
rect 152188 191088 152240 191140
rect 157616 191088 157668 191140
rect 158444 191088 158496 191140
rect 160376 191088 160428 191140
rect 161296 191088 161348 191140
rect 161664 191088 161716 191140
rect 162584 191088 162636 191140
rect 170680 191088 170732 191140
rect 171508 191088 171560 191140
rect 174268 191088 174320 191140
rect 174728 191088 174780 191140
rect 160192 191020 160244 191072
rect 160928 191020 160980 191072
rect 171968 191020 172020 191072
rect 172704 191020 172756 191072
rect 160100 190952 160152 191004
rect 161020 190952 161072 191004
rect 145656 190816 145708 190868
rect 151912 190816 151964 190868
rect 151912 190680 151964 190732
rect 152648 190680 152700 190732
rect 141424 190544 141476 190596
rect 143816 190544 143868 190596
rect 173900 190544 173952 190596
rect 174176 190544 174228 190596
rect 113824 190408 113876 190460
rect 141884 190408 141936 190460
rect 174176 190408 174228 190460
rect 174544 190408 174596 190460
rect 110972 190340 111024 190392
rect 138664 190340 138716 190392
rect 109960 190272 110012 190324
rect 139952 190272 140004 190324
rect 112352 190204 112404 190256
rect 141240 190204 141292 190256
rect 157248 190204 157300 190256
rect 158812 190204 158864 190256
rect 107568 190136 107620 190188
rect 140228 190136 140280 190188
rect 101772 190068 101824 190120
rect 134064 190068 134116 190120
rect 101864 190000 101916 190052
rect 134800 190000 134852 190052
rect 102968 189932 103020 189984
rect 136180 189932 136232 189984
rect 101588 189864 101640 189916
rect 134984 189864 135036 189916
rect 150992 189864 151044 189916
rect 151636 189864 151688 189916
rect 102048 189796 102100 189848
rect 135904 189796 135956 189848
rect 101956 189728 102008 189780
rect 135260 189728 135312 189780
rect 134156 189660 134208 189712
rect 134432 189660 134484 189712
rect 162860 189660 162912 189712
rect 163228 189660 163280 189712
rect 126428 189456 126480 189508
rect 149704 189456 149756 189508
rect 149704 189320 149756 189372
rect 153200 189320 153252 189372
rect 162860 189320 162912 189372
rect 163964 189320 164016 189372
rect 3424 188980 3476 189032
rect 120632 188980 120684 189032
rect 169760 188980 169812 189032
rect 170956 188980 171008 189032
rect 132868 188912 132920 188964
rect 133420 188912 133472 188964
rect 171416 188912 171468 188964
rect 171600 188912 171652 188964
rect 154764 188776 154816 188828
rect 155500 188776 155552 188828
rect 169944 188640 169996 188692
rect 170588 188640 170640 188692
rect 131764 188436 131816 188488
rect 139400 188436 139452 188488
rect 125508 188368 125560 188420
rect 143540 188368 143592 188420
rect 176844 188368 176896 188420
rect 177948 188368 178000 188420
rect 130384 188300 130436 188352
rect 139308 188300 139360 188352
rect 176752 188300 176804 188352
rect 177764 188300 177816 188352
rect 135628 188232 135680 188284
rect 136272 188232 136324 188284
rect 176660 187892 176712 187944
rect 178132 187892 178184 187944
rect 132684 187484 132736 187536
rect 133880 187484 133932 187536
rect 126244 187416 126296 187468
rect 150072 187416 150124 187468
rect 149520 186328 149572 186380
rect 150164 186328 150216 186380
rect 148692 185784 148744 185836
rect 154580 185784 154632 185836
rect 141148 185444 141200 185496
rect 142068 185444 142120 185496
rect 161480 185104 161532 185156
rect 162124 185104 162176 185156
rect 145748 184968 145800 185020
rect 156512 184968 156564 185020
rect 175280 184968 175332 185020
rect 176108 184968 176160 185020
rect 153476 184696 153528 184748
rect 154304 184696 154356 184748
rect 175556 184696 175608 184748
rect 175924 184696 175976 184748
rect 159272 184016 159324 184068
rect 160008 184016 160060 184068
rect 172612 183472 172664 183524
rect 172888 183472 172940 183524
rect 164332 183336 164384 183388
rect 165344 183336 165396 183388
rect 129096 183064 129148 183116
rect 137376 183064 137428 183116
rect 127624 181976 127676 182028
rect 141608 181976 141660 182028
rect 171140 181432 171192 181484
rect 171324 181432 171376 181484
rect 129280 180276 129332 180328
rect 149888 180276 149940 180328
rect 145840 179120 145892 179172
rect 146576 179120 146628 179172
rect 188620 178032 188672 178084
rect 580172 178032 580224 178084
rect 189816 165588 189868 165640
rect 580172 165588 580224 165640
rect 168656 155320 168708 155372
rect 203432 155320 203484 155372
rect 169576 155252 169628 155304
rect 203524 155252 203576 155304
rect 167276 155184 167328 155236
rect 202328 155184 202380 155236
rect 163136 153144 163188 153196
rect 185952 153144 186004 153196
rect 161756 153076 161808 153128
rect 185584 153076 185636 153128
rect 160284 153008 160336 153060
rect 184296 153008 184348 153060
rect 161848 152940 161900 152992
rect 186044 152940 186096 152992
rect 160468 152872 160520 152924
rect 185676 152872 185728 152924
rect 158996 152804 159048 152856
rect 184388 152804 184440 152856
rect 160376 152736 160428 152788
rect 186136 152736 186188 152788
rect 160008 152668 160060 152720
rect 184756 152668 184808 152720
rect 167092 152600 167144 152652
rect 199200 152600 199252 152652
rect 164608 152532 164660 152584
rect 199292 152532 199344 152584
rect 165712 152464 165764 152516
rect 200856 152464 200908 152516
rect 163228 152396 163280 152448
rect 185860 152396 185912 152448
rect 165804 152328 165856 152380
rect 184572 152328 184624 152380
rect 168380 152260 168432 152312
rect 183192 152260 183244 152312
rect 100208 151172 100260 151224
rect 132684 151172 132736 151224
rect 100300 151104 100352 151156
rect 134248 151104 134300 151156
rect 100392 151036 100444 151088
rect 134432 151036 134484 151088
rect 176936 150356 176988 150408
rect 202788 150356 202840 150408
rect 176844 150288 176896 150340
rect 201408 150288 201460 150340
rect 184204 150220 184256 150272
rect 202236 150220 202288 150272
rect 175556 150152 175608 150204
rect 204536 150152 204588 150204
rect 175464 150084 175516 150136
rect 204628 150084 204680 150136
rect 174360 150016 174412 150068
rect 203708 150016 203760 150068
rect 174176 149948 174228 150000
rect 203616 149948 203668 150000
rect 175648 149880 175700 149932
rect 206192 149880 206244 149932
rect 175280 149812 175332 149864
rect 206284 149812 206336 149864
rect 175372 149744 175424 149796
rect 206376 149744 206428 149796
rect 148968 149676 149020 149728
rect 184664 149676 184716 149728
rect 3424 149064 3476 149116
rect 9588 149064 9640 149116
rect 126612 148996 126664 149048
rect 154856 148996 154908 149048
rect 113364 148928 113416 148980
rect 142620 148928 142672 148980
rect 125048 148860 125100 148912
rect 153476 148860 153528 148912
rect 123116 148792 123168 148844
rect 152096 148792 152148 148844
rect 102692 148724 102744 148776
rect 131856 148724 131908 148776
rect 178684 148724 178736 148776
rect 195520 148724 195572 148776
rect 124496 148656 124548 148708
rect 156144 148656 156196 148708
rect 164424 148656 164476 148708
rect 186964 148656 187016 148708
rect 104072 148588 104124 148640
rect 135628 148588 135680 148640
rect 160192 148588 160244 148640
rect 184112 148588 184164 148640
rect 120448 148520 120500 148572
rect 153292 148520 153344 148572
rect 167000 148520 167052 148572
rect 198280 148520 198332 148572
rect 117596 148452 117648 148504
rect 152188 148452 152240 148504
rect 163044 148452 163096 148504
rect 196992 148452 197044 148504
rect 116216 148384 116268 148436
rect 151728 148384 151780 148436
rect 164516 148384 164568 148436
rect 199476 148384 199528 148436
rect 9588 148316 9640 148368
rect 180892 148316 180944 148368
rect 196716 148316 196768 148368
rect 113548 148248 113600 148300
rect 142988 148248 143040 148300
rect 116124 148180 116176 148232
rect 142528 148180 142580 148232
rect 126520 148112 126572 148164
rect 148324 148112 148376 148164
rect 178224 147568 178276 147620
rect 196532 147568 196584 147620
rect 178040 147500 178092 147552
rect 198096 147500 198148 147552
rect 171232 147432 171284 147484
rect 194324 147432 194376 147484
rect 172796 147364 172848 147416
rect 195336 147364 195388 147416
rect 172888 147296 172940 147348
rect 196532 147296 196584 147348
rect 113916 147228 113968 147280
rect 126980 147228 127032 147280
rect 170036 147228 170088 147280
rect 193956 147228 194008 147280
rect 115020 147160 115072 147212
rect 137284 147160 137336 147212
rect 171324 147160 171376 147212
rect 195428 147160 195480 147212
rect 114928 147092 114980 147144
rect 140964 147092 141016 147144
rect 172704 147092 172756 147144
rect 198372 147092 198424 147144
rect 112260 147024 112312 147076
rect 138480 147024 138532 147076
rect 171416 147024 171468 147076
rect 196716 147024 196768 147076
rect 117504 146956 117556 147008
rect 145656 146956 145708 147008
rect 171508 146956 171560 147008
rect 198096 146956 198148 147008
rect 110880 146888 110932 146940
rect 139768 146888 139820 146940
rect 173992 146888 174044 146940
rect 206468 146888 206520 146940
rect 179604 146820 179656 146872
rect 197912 146820 197964 146872
rect 178408 146752 178460 146804
rect 195152 146752 195204 146804
rect 179696 146684 179748 146736
rect 193772 146684 193824 146736
rect 116860 146208 116912 146260
rect 131304 146208 131356 146260
rect 178316 146208 178368 146260
rect 188252 146208 188304 146260
rect 116768 146140 116820 146192
rect 131212 146140 131264 146192
rect 178132 146140 178184 146192
rect 191288 146140 191340 146192
rect 121920 146072 121972 146124
rect 146668 146072 146720 146124
rect 175556 146072 175608 146124
rect 197820 146072 197872 146124
rect 121828 146004 121880 146056
rect 149520 146004 149572 146056
rect 161572 146004 161624 146056
rect 188344 146004 188396 146056
rect 118792 145936 118844 145988
rect 146576 145936 146628 145988
rect 165620 145936 165672 145988
rect 194140 145936 194192 145988
rect 118976 145868 119028 145920
rect 146484 145868 146536 145920
rect 161480 145868 161532 145920
rect 190092 145868 190144 145920
rect 119068 145800 119120 145852
rect 147680 145800 147732 145852
rect 162952 145800 163004 145852
rect 194232 145800 194284 145852
rect 120356 145732 120408 145784
rect 153108 145732 153160 145784
rect 160100 145732 160152 145784
rect 195152 145732 195204 145784
rect 116400 145664 116452 145716
rect 150624 145664 150676 145716
rect 159916 145664 159968 145716
rect 191380 145664 191432 145716
rect 119988 145596 120040 145648
rect 160100 145596 160152 145648
rect 161664 145596 161716 145648
rect 192944 145596 192996 145648
rect 3516 145528 3568 145580
rect 179788 145528 179840 145580
rect 189632 145528 189684 145580
rect 116768 145460 116820 145512
rect 130568 145460 130620 145512
rect 180432 145460 180484 145512
rect 190184 145460 190236 145512
rect 116952 145392 117004 145444
rect 129740 145392 129792 145444
rect 180340 145392 180392 145444
rect 190000 145392 190052 145444
rect 179420 145324 179472 145376
rect 189724 145324 189776 145376
rect 183008 144848 183060 144900
rect 192760 144848 192812 144900
rect 179512 144780 179564 144832
rect 193588 144780 193640 144832
rect 118056 144712 118108 144764
rect 130016 144712 130068 144764
rect 173808 144712 173860 144764
rect 190920 144712 190972 144764
rect 119712 144644 119764 144696
rect 138112 144644 138164 144696
rect 170772 144644 170824 144696
rect 192024 144644 192076 144696
rect 116492 144576 116544 144628
rect 143816 144576 143868 144628
rect 172428 144576 172480 144628
rect 194968 144576 195020 144628
rect 122380 144508 122432 144560
rect 152648 144508 152700 144560
rect 169116 144508 169168 144560
rect 192392 144508 192444 144560
rect 122564 144440 122616 144492
rect 153844 144440 153896 144492
rect 158168 144440 158220 144492
rect 192852 144440 192904 144492
rect 119712 144372 119764 144424
rect 150532 144372 150584 144424
rect 152556 144372 152608 144424
rect 186412 144372 186464 144424
rect 116860 144304 116912 144356
rect 148600 144304 148652 144356
rect 156420 144304 156472 144356
rect 191012 144304 191064 144356
rect 115296 144236 115348 144288
rect 131396 144236 131448 144288
rect 188620 144236 188672 144288
rect 116676 144168 116728 144220
rect 129372 144168 129424 144220
rect 130016 144168 130068 144220
rect 189816 144168 189868 144220
rect 188160 143896 188212 143948
rect 188160 143624 188212 143676
rect 119988 143556 120040 143608
rect 145288 143556 145340 143608
rect 187884 143556 187936 143608
rect 188068 143556 188120 143608
rect 113732 143488 113784 143540
rect 123852 143488 123904 143540
rect 124036 143488 124088 143540
rect 124588 143488 124640 143540
rect 119804 143420 119856 143472
rect 131488 143488 131540 143540
rect 131580 143488 131632 143540
rect 580356 143488 580408 143540
rect 131120 143420 131172 143472
rect 137560 143420 137612 143472
rect 146300 143420 146352 143472
rect 149152 143420 149204 143472
rect 175464 143420 175516 143472
rect 179512 143420 179564 143472
rect 181536 143420 181588 143472
rect 187056 143420 187108 143472
rect 187424 143420 187476 143472
rect 187884 143420 187936 143472
rect 120816 143352 120868 143404
rect 133144 143352 133196 143404
rect 174636 143352 174688 143404
rect 179696 143352 179748 143404
rect 185676 143352 185728 143404
rect 193680 143420 193732 143472
rect 115112 143284 115164 143336
rect 123760 143284 123812 143336
rect 123852 143284 123904 143336
rect 124864 143284 124916 143336
rect 131212 143284 131264 143336
rect 135444 143284 135496 143336
rect 172980 143284 173032 143336
rect 178408 143284 178460 143336
rect 122196 143216 122248 143268
rect 136640 143216 136692 143268
rect 176568 143216 176620 143268
rect 185952 143284 186004 143336
rect 195060 143352 195112 143404
rect 189540 143284 189592 143336
rect 114008 143148 114060 143200
rect 129556 143148 129608 143200
rect 129832 143148 129884 143200
rect 135904 143148 135956 143200
rect 169668 143148 169720 143200
rect 179604 143148 179656 143200
rect 118332 143080 118384 143132
rect 134800 143080 134852 143132
rect 177396 143080 177448 143132
rect 179420 143080 179472 143132
rect 115572 143012 115624 143064
rect 132592 143012 132644 143064
rect 170220 143012 170272 143064
rect 188436 143216 188488 143268
rect 195244 143284 195296 143336
rect 182456 143148 182508 143200
rect 196440 143148 196492 143200
rect 184480 143080 184532 143132
rect 198004 143080 198056 143132
rect 191104 143012 191156 143064
rect 120908 142944 120960 142996
rect 139768 142944 139820 142996
rect 168288 142944 168340 142996
rect 182088 142944 182140 142996
rect 121000 142876 121052 142928
rect 141516 142876 141568 142928
rect 166908 142876 166960 142928
rect 191196 142876 191248 142928
rect 121092 142808 121144 142860
rect 151360 142808 151412 142860
rect 158628 142808 158680 142860
rect 188252 142808 188304 142860
rect 119620 142740 119672 142792
rect 128452 142740 128504 142792
rect 129372 142740 129424 142792
rect 131580 142740 131632 142792
rect 183100 142740 183152 142792
rect 190920 142740 190972 142792
rect 123760 142672 123812 142724
rect 129096 142672 129148 142724
rect 131212 142672 131264 142724
rect 131396 142672 131448 142724
rect 177948 142672 178000 142724
rect 178224 142672 178276 142724
rect 182088 142672 182140 142724
rect 189448 142672 189500 142724
rect 183744 142604 183796 142656
rect 188436 142604 188488 142656
rect 129924 142264 129976 142316
rect 134248 142264 134300 142316
rect 129740 142196 129792 142248
rect 133880 142196 133932 142248
rect 155684 142196 155736 142248
rect 157340 142196 157392 142248
rect 159180 142196 159232 142248
rect 161480 142196 161532 142248
rect 3424 142128 3476 142180
rect 183744 142128 183796 142180
rect 185952 142128 186004 142180
rect 187884 142128 187936 142180
rect 161480 142060 161532 142112
rect 192300 142060 192352 142112
rect 118424 141992 118476 142044
rect 126888 141992 126940 142044
rect 115480 141924 115532 141976
rect 127348 141924 127400 141976
rect 180340 141924 180392 141976
rect 187240 141924 187292 141976
rect 115296 141856 115348 141908
rect 130384 141856 130436 141908
rect 182088 141856 182140 141908
rect 192116 141856 192168 141908
rect 116584 141788 116636 141840
rect 131764 141788 131816 141840
rect 183192 141788 183244 141840
rect 196440 141788 196492 141840
rect 113640 141720 113692 141772
rect 132868 141720 132920 141772
rect 175188 141720 175240 141772
rect 187332 141720 187384 141772
rect 118148 141652 118200 141704
rect 140320 141652 140372 141704
rect 173532 141652 173584 141704
rect 190828 141652 190880 141704
rect 114192 141584 114244 141636
rect 137008 141584 137060 141636
rect 171876 141584 171928 141636
rect 189356 141584 189408 141636
rect 119988 141516 120040 141568
rect 151912 141516 151964 141568
rect 167460 141516 167512 141568
rect 192208 141516 192260 141568
rect 119528 141448 119580 141500
rect 142252 141448 142304 141500
rect 164332 141448 164384 141500
rect 189540 141448 189592 141500
rect 119436 141380 119488 141432
rect 153568 141380 153620 141432
rect 162860 141380 162912 141432
rect 198004 141380 198056 141432
rect 121000 141312 121052 141364
rect 126520 141312 126572 141364
rect 118240 141244 118292 141296
rect 125416 141244 125468 141296
rect 129556 141040 129608 141092
rect 187976 141040 188028 141092
rect 117780 140972 117832 141024
rect 182088 140972 182140 141024
rect 8944 140904 8996 140956
rect 182824 140904 182876 140956
rect 184572 140904 184624 140956
rect 188436 140904 188488 140956
rect 126888 140836 126940 140888
rect 464344 140836 464396 140888
rect 124588 140768 124640 140820
rect 124956 140768 125008 140820
rect 485044 140768 485096 140820
rect 125968 140700 126020 140752
rect 126612 140700 126664 140752
rect 126980 140700 127032 140752
rect 127716 140700 127768 140752
rect 131304 140700 131356 140752
rect 132316 140700 132368 140752
rect 178040 140700 178092 140752
rect 178960 140700 179012 140752
rect 184756 140700 184808 140752
rect 192024 140700 192076 140752
rect 120632 140632 120684 140684
rect 126336 140632 126388 140684
rect 172520 140632 172572 140684
rect 180156 140632 180208 140684
rect 118148 140564 118200 140616
rect 126244 140564 126296 140616
rect 171692 140564 171744 140616
rect 179052 140564 179104 140616
rect 180248 140564 180300 140616
rect 188252 140564 188304 140616
rect 117872 140496 117924 140548
rect 126428 140496 126480 140548
rect 184112 140496 184164 140548
rect 188620 140496 188672 140548
rect 120724 140428 120776 140480
rect 147036 140428 147088 140480
rect 182916 140428 182968 140480
rect 190828 140428 190880 140480
rect 119252 140360 119304 140412
rect 146944 140360 146996 140412
rect 185768 140360 185820 140412
rect 193864 140360 193916 140412
rect 120540 140292 120592 140344
rect 148232 140292 148284 140344
rect 181444 140292 181496 140344
rect 189908 140292 189960 140344
rect 117964 140224 118016 140276
rect 145564 140224 145616 140276
rect 180064 140224 180116 140276
rect 189356 140224 189408 140276
rect 118056 140156 118108 140208
rect 147956 140156 148008 140208
rect 184296 140156 184348 140208
rect 189816 140156 189868 140208
rect 121920 140088 121972 140140
rect 152464 140088 152516 140140
rect 169852 140088 169904 140140
rect 119344 140020 119396 140072
rect 129280 140020 129332 140072
rect 129740 140020 129792 140072
rect 184664 140088 184716 140140
rect 187240 140088 187292 140140
rect 130016 139952 130068 140004
rect 130476 139952 130528 140004
rect 187332 140020 187384 140072
rect 188068 139952 188120 140004
rect 184388 139884 184440 139936
rect 194048 139952 194100 140004
rect 188620 139884 188672 139936
rect 192300 139884 192352 139936
rect 171140 139816 171192 139868
rect 128820 139748 128872 139800
rect 183468 139748 183520 139800
rect 125876 139680 125928 139732
rect 184664 139680 184716 139732
rect 196256 139816 196308 139868
rect 118700 139612 118752 139664
rect 180064 139612 180116 139664
rect 122840 139544 122892 139596
rect 123852 139544 123904 139596
rect 184572 139544 184624 139596
rect 31024 139476 31076 139528
rect 181168 139476 181220 139528
rect 185584 139476 185636 139528
rect 187424 139476 187476 139528
rect 13084 139408 13136 139460
rect 185032 139408 185084 139460
rect 186136 139408 186188 139460
rect 187148 139408 187200 139460
rect 186044 139340 186096 139392
rect 186872 139340 186924 139392
rect 188252 139408 188304 139460
rect 187976 139340 188028 139392
rect 580172 139340 580224 139392
rect 187976 139204 188028 139256
rect 3516 137912 3568 137964
rect 118700 137912 118752 137964
rect 3148 111732 3200 111784
rect 31024 111732 31076 111784
rect 464344 86912 464396 86964
rect 580172 86912 580224 86964
rect 3516 85484 3568 85536
rect 117780 85484 117832 85536
rect 123024 81064 123076 81116
rect 119068 80928 119120 80980
rect 122288 80860 122340 80912
rect 123024 80860 123076 80912
rect 108212 80792 108264 80844
rect 85580 80724 85632 80776
rect 105636 80724 105688 80776
rect 71780 80656 71832 80708
rect 108212 80656 108264 80708
rect 119988 80656 120040 80708
rect 104256 80384 104308 80436
rect 131948 80656 132000 80708
rect 132132 80656 132184 80708
rect 132224 80588 132276 80640
rect 132224 80384 132276 80436
rect 131856 80316 131908 80368
rect 104164 80180 104216 80232
rect 110972 80044 111024 80096
rect 131028 80248 131080 80300
rect 127532 80180 127584 80232
rect 131948 80044 132000 80096
rect 132730 79908 132782 79960
rect 133098 79908 133150 79960
rect 126980 79840 127032 79892
rect 132914 79840 132966 79892
rect 119252 79636 119304 79688
rect 132408 79636 132460 79688
rect 106832 79568 106884 79620
rect 113824 79500 113876 79552
rect 125692 79500 125744 79552
rect 127440 79500 127492 79552
rect 111064 79432 111116 79484
rect 125600 79432 125652 79484
rect 127532 79432 127584 79484
rect 133052 79568 133104 79620
rect 133374 79908 133426 79960
rect 133650 79908 133702 79960
rect 133466 79840 133518 79892
rect 133420 79704 133472 79756
rect 133328 79568 133380 79620
rect 132868 79500 132920 79552
rect 133834 79908 133886 79960
rect 134018 79908 134070 79960
rect 134110 79908 134162 79960
rect 134662 79908 134714 79960
rect 134846 79908 134898 79960
rect 133696 79636 133748 79688
rect 133604 79568 133656 79620
rect 133880 79772 133932 79824
rect 133972 79772 134024 79824
rect 134478 79840 134530 79892
rect 134202 79772 134254 79824
rect 134064 79704 134116 79756
rect 134156 79568 134208 79620
rect 134340 79568 134392 79620
rect 134938 79840 134990 79892
rect 134662 79772 134714 79824
rect 134754 79704 134806 79756
rect 111248 79364 111300 79416
rect 128360 79364 128412 79416
rect 131028 79364 131080 79416
rect 100116 79296 100168 79348
rect 100300 79296 100352 79348
rect 112444 79296 112496 79348
rect 130384 79296 130436 79348
rect 132684 79364 132736 79416
rect 134340 79432 134392 79484
rect 134616 79500 134668 79552
rect 134892 79636 134944 79688
rect 135306 79908 135358 79960
rect 136226 79908 136278 79960
rect 136318 79908 136370 79960
rect 136594 79908 136646 79960
rect 136962 79908 137014 79960
rect 137054 79908 137106 79960
rect 137238 79908 137290 79960
rect 137514 79908 137566 79960
rect 138250 79908 138302 79960
rect 138894 79908 138946 79960
rect 139078 79908 139130 79960
rect 139446 79908 139498 79960
rect 139630 79908 139682 79960
rect 139722 79908 139774 79960
rect 140642 79908 140694 79960
rect 140826 79908 140878 79960
rect 141010 79908 141062 79960
rect 141194 79908 141246 79960
rect 141562 79908 141614 79960
rect 135076 79432 135128 79484
rect 135766 79840 135818 79892
rect 135950 79840 136002 79892
rect 136042 79840 136094 79892
rect 135582 79772 135634 79824
rect 135260 79568 135312 79620
rect 135628 79568 135680 79620
rect 135996 79636 136048 79688
rect 136410 79772 136462 79824
rect 136456 79636 136508 79688
rect 136824 79704 136876 79756
rect 136180 79568 136232 79620
rect 136364 79568 136416 79620
rect 136548 79568 136600 79620
rect 136088 79500 136140 79552
rect 136916 79636 136968 79688
rect 137100 79636 137152 79688
rect 137422 79840 137474 79892
rect 137790 79840 137842 79892
rect 137468 79704 137520 79756
rect 137836 79636 137888 79688
rect 138112 79636 138164 79688
rect 138986 79840 139038 79892
rect 138388 79636 138440 79688
rect 138480 79636 138532 79688
rect 137008 79568 137060 79620
rect 137284 79568 137336 79620
rect 139814 79840 139866 79892
rect 139492 79636 139544 79688
rect 139584 79568 139636 79620
rect 140182 79840 140234 79892
rect 140458 79840 140510 79892
rect 139768 79500 139820 79552
rect 140044 79500 140096 79552
rect 135536 79432 135588 79484
rect 135720 79432 135772 79484
rect 137008 79432 137060 79484
rect 137928 79432 137980 79484
rect 140320 79636 140372 79688
rect 140596 79772 140648 79824
rect 141056 79704 141108 79756
rect 141286 79840 141338 79892
rect 141470 79840 141522 79892
rect 141654 79840 141706 79892
rect 140780 79568 140832 79620
rect 141148 79636 141200 79688
rect 141056 79568 141108 79620
rect 141240 79500 141292 79552
rect 141332 79500 141384 79552
rect 141516 79432 141568 79484
rect 141838 79908 141890 79960
rect 142390 79908 142442 79960
rect 142482 79840 142534 79892
rect 143402 79908 143454 79960
rect 143586 79908 143638 79960
rect 142206 79772 142258 79824
rect 141976 79636 142028 79688
rect 142068 79500 142120 79552
rect 142942 79840 142994 79892
rect 143218 79840 143270 79892
rect 143494 79840 143546 79892
rect 142758 79772 142810 79824
rect 142620 79568 142672 79620
rect 142804 79568 142856 79620
rect 142896 79500 142948 79552
rect 142528 79432 142580 79484
rect 143678 79840 143730 79892
rect 143540 79704 143592 79756
rect 143172 79432 143224 79484
rect 143448 79432 143500 79484
rect 141148 79364 141200 79416
rect 141608 79364 141660 79416
rect 144138 79840 144190 79892
rect 143954 79772 144006 79824
rect 143816 79636 143868 79688
rect 144000 79636 144052 79688
rect 144368 79500 144420 79552
rect 144782 79908 144834 79960
rect 144874 79908 144926 79960
rect 144598 79840 144650 79892
rect 145702 79908 145754 79960
rect 145794 79908 145846 79960
rect 145978 79908 146030 79960
rect 146070 79908 146122 79960
rect 146254 79908 146306 79960
rect 144828 79772 144880 79824
rect 144644 79636 144696 79688
rect 144552 79500 144604 79552
rect 145518 79840 145570 79892
rect 145564 79704 145616 79756
rect 145196 79500 145248 79552
rect 145656 79636 145708 79688
rect 145656 79500 145708 79552
rect 123300 79228 123352 79280
rect 144460 79296 144512 79348
rect 145012 79432 145064 79484
rect 146346 79840 146398 79892
rect 146530 79840 146582 79892
rect 146024 79772 146076 79824
rect 146116 79772 146168 79824
rect 146300 79704 146352 79756
rect 146714 79908 146766 79960
rect 146668 79704 146720 79756
rect 146576 79568 146628 79620
rect 146990 79908 147042 79960
rect 147082 79908 147134 79960
rect 147174 79908 147226 79960
rect 147450 79908 147502 79960
rect 147542 79908 147594 79960
rect 147910 79908 147962 79960
rect 148094 79908 148146 79960
rect 146944 79704 146996 79756
rect 147220 79704 147272 79756
rect 147496 79704 147548 79756
rect 147036 79636 147088 79688
rect 147128 79636 147180 79688
rect 147220 79568 147272 79620
rect 147404 79500 147456 79552
rect 147588 79500 147640 79552
rect 147818 79840 147870 79892
rect 147772 79704 147824 79756
rect 147864 79636 147916 79688
rect 148278 79840 148330 79892
rect 148370 79840 148422 79892
rect 148232 79704 148284 79756
rect 148324 79636 148376 79688
rect 147772 79568 147824 79620
rect 147956 79568 148008 79620
rect 148830 79908 148882 79960
rect 148922 79908 148974 79960
rect 149106 79908 149158 79960
rect 149198 79908 149250 79960
rect 148692 79636 148744 79688
rect 146760 79432 146812 79484
rect 148600 79432 148652 79484
rect 147404 79364 147456 79416
rect 148876 79772 148928 79824
rect 149152 79772 149204 79824
rect 149060 79636 149112 79688
rect 149244 79568 149296 79620
rect 149658 79908 149710 79960
rect 149750 79908 149802 79960
rect 149842 79908 149894 79960
rect 149474 79840 149526 79892
rect 149704 79772 149756 79824
rect 149796 79704 149848 79756
rect 150118 79840 150170 79892
rect 149888 79636 149940 79688
rect 187424 80860 187476 80912
rect 188620 80860 188672 80912
rect 206100 80860 206152 80912
rect 234620 80860 234672 80912
rect 177948 80656 178000 80708
rect 178040 80656 178092 80708
rect 178592 80656 178644 80708
rect 186780 80792 186832 80844
rect 252560 80792 252612 80844
rect 188160 80724 188212 80776
rect 270500 80724 270552 80776
rect 188620 80656 188672 80708
rect 189264 80656 189316 80708
rect 288440 80656 288492 80708
rect 187424 80452 187476 80504
rect 150670 79908 150722 79960
rect 150946 79840 150998 79892
rect 151222 79908 151274 79960
rect 151406 79908 151458 79960
rect 152050 79908 152102 79960
rect 152418 79908 152470 79960
rect 152878 79908 152930 79960
rect 152970 79908 153022 79960
rect 153430 79908 153482 79960
rect 154166 79908 154218 79960
rect 154258 79908 154310 79960
rect 154350 79908 154402 79960
rect 154442 79908 154494 79960
rect 154810 79908 154862 79960
rect 154994 79908 155046 79960
rect 155178 79908 155230 79960
rect 151176 79772 151228 79824
rect 150348 79704 150400 79756
rect 151866 79840 151918 79892
rect 150440 79636 150492 79688
rect 151360 79636 151412 79688
rect 152234 79772 152286 79824
rect 152188 79636 152240 79688
rect 150992 79568 151044 79620
rect 151820 79568 151872 79620
rect 152694 79840 152746 79892
rect 152648 79636 152700 79688
rect 152556 79568 152608 79620
rect 153154 79840 153206 79892
rect 153706 79840 153758 79892
rect 152970 79772 153022 79824
rect 153016 79636 153068 79688
rect 153890 79772 153942 79824
rect 153292 79568 153344 79620
rect 153752 79568 153804 79620
rect 150164 79500 150216 79552
rect 153476 79500 153528 79552
rect 154212 79772 154264 79824
rect 154396 79772 154448 79824
rect 154304 79636 154356 79688
rect 154626 79840 154678 79892
rect 154764 79704 154816 79756
rect 154672 79636 154724 79688
rect 153936 79568 153988 79620
rect 154948 79568 155000 79620
rect 178776 80316 178828 80368
rect 185216 80248 185268 80300
rect 156282 79908 156334 79960
rect 156374 79908 156426 79960
rect 156558 79908 156610 79960
rect 155362 79840 155414 79892
rect 155914 79840 155966 79892
rect 156190 79840 156242 79892
rect 155132 79500 155184 79552
rect 155454 79772 155506 79824
rect 155500 79636 155552 79688
rect 156144 79500 156196 79552
rect 156236 79432 156288 79484
rect 156742 79908 156794 79960
rect 156926 79908 156978 79960
rect 157294 79908 157346 79960
rect 156834 79840 156886 79892
rect 156788 79704 156840 79756
rect 156604 79636 156656 79688
rect 156696 79568 156748 79620
rect 156880 79636 156932 79688
rect 157248 79568 157300 79620
rect 157064 79432 157116 79484
rect 152648 79296 152700 79348
rect 156972 79296 157024 79348
rect 157478 79908 157530 79960
rect 157570 79908 157622 79960
rect 157662 79908 157714 79960
rect 157754 79908 157806 79960
rect 157524 79636 157576 79688
rect 157524 79500 157576 79552
rect 158214 79908 158266 79960
rect 158490 79908 158542 79960
rect 158030 79840 158082 79892
rect 157938 79772 157990 79824
rect 158398 79840 158450 79892
rect 158766 79908 158818 79960
rect 158858 79908 158910 79960
rect 159042 79908 159094 79960
rect 158812 79772 158864 79824
rect 159134 79840 159186 79892
rect 159088 79704 159140 79756
rect 159594 79908 159646 79960
rect 159686 79908 159738 79960
rect 159502 79772 159554 79824
rect 158260 79636 158312 79688
rect 158352 79636 158404 79688
rect 158536 79636 158588 79688
rect 158628 79636 158680 79688
rect 158904 79636 158956 79688
rect 159640 79636 159692 79688
rect 158444 79568 158496 79620
rect 159548 79568 159600 79620
rect 160054 79908 160106 79960
rect 160238 79908 160290 79960
rect 160422 79908 160474 79960
rect 160606 79908 160658 79960
rect 160146 79840 160198 79892
rect 160330 79840 160382 79892
rect 160008 79636 160060 79688
rect 160284 79704 160336 79756
rect 160560 79636 160612 79688
rect 160100 79568 160152 79620
rect 160376 79568 160428 79620
rect 160882 79908 160934 79960
rect 160974 79908 161026 79960
rect 161158 79908 161210 79960
rect 161710 79908 161762 79960
rect 160744 79568 160796 79620
rect 161342 79840 161394 79892
rect 161204 79772 161256 79824
rect 161664 79772 161716 79824
rect 161296 79704 161348 79756
rect 161020 79636 161072 79688
rect 161986 79908 162038 79960
rect 162078 79908 162130 79960
rect 162262 79908 162314 79960
rect 161894 79840 161946 79892
rect 161940 79636 161992 79688
rect 162032 79568 162084 79620
rect 157892 79500 157944 79552
rect 159824 79500 159876 79552
rect 160836 79500 160888 79552
rect 162124 79500 162176 79552
rect 162538 79840 162590 79892
rect 163274 79908 163326 79960
rect 163458 79908 163510 79960
rect 163826 79908 163878 79960
rect 162814 79840 162866 79892
rect 162998 79840 163050 79892
rect 163182 79840 163234 79892
rect 162584 79636 162636 79688
rect 162860 79636 162912 79688
rect 162492 79500 162544 79552
rect 163136 79636 163188 79688
rect 163136 79500 163188 79552
rect 163366 79840 163418 79892
rect 157800 79432 157852 79484
rect 158168 79432 158220 79484
rect 162952 79432 163004 79484
rect 157984 79364 158036 79416
rect 158076 79364 158128 79416
rect 162400 79364 162452 79416
rect 162768 79364 162820 79416
rect 163734 79840 163786 79892
rect 163642 79772 163694 79824
rect 163780 79704 163832 79756
rect 163596 79568 163648 79620
rect 163688 79500 163740 79552
rect 163504 79432 163556 79484
rect 164102 79840 164154 79892
rect 164470 79840 164522 79892
rect 164378 79772 164430 79824
rect 164148 79704 164200 79756
rect 164654 79772 164706 79824
rect 164424 79636 164476 79688
rect 164608 79636 164660 79688
rect 165022 79908 165074 79960
rect 165114 79908 165166 79960
rect 164056 79500 164108 79552
rect 164792 79500 164844 79552
rect 165298 79840 165350 79892
rect 165206 79772 165258 79824
rect 165160 79636 165212 79688
rect 165252 79568 165304 79620
rect 165942 79908 165994 79960
rect 166126 79908 166178 79960
rect 166034 79840 166086 79892
rect 166402 79908 166454 79960
rect 166494 79908 166546 79960
rect 166770 79908 166822 79960
rect 165758 79772 165810 79824
rect 165896 79772 165948 79824
rect 165804 79568 165856 79620
rect 165436 79500 165488 79552
rect 165620 79500 165672 79552
rect 166448 79636 166500 79688
rect 166356 79568 166408 79620
rect 166862 79840 166914 79892
rect 166816 79568 166868 79620
rect 167230 79908 167282 79960
rect 167506 79908 167558 79960
rect 167874 79908 167926 79960
rect 167966 79908 168018 79960
rect 167138 79840 167190 79892
rect 167414 79840 167466 79892
rect 167092 79568 167144 79620
rect 167184 79500 167236 79552
rect 166540 79432 166592 79484
rect 167460 79704 167512 79756
rect 167782 79840 167834 79892
rect 167920 79772 167972 79824
rect 167828 79704 167880 79756
rect 168518 79908 168570 79960
rect 168794 79908 168846 79960
rect 169070 79908 169122 79960
rect 167644 79636 167696 79688
rect 168288 79636 168340 79688
rect 169024 79568 169076 79620
rect 169346 79908 169398 79960
rect 169530 79908 169582 79960
rect 169714 79908 169766 79960
rect 170266 79908 170318 79960
rect 170358 79908 170410 79960
rect 169622 79840 169674 79892
rect 169392 79636 169444 79688
rect 169484 79636 169536 79688
rect 169576 79568 169628 79620
rect 169898 79840 169950 79892
rect 170174 79840 170226 79892
rect 169852 79568 169904 79620
rect 169392 79500 169444 79552
rect 168748 79432 168800 79484
rect 169760 79432 169812 79484
rect 170128 79704 170180 79756
rect 177764 80180 177816 80232
rect 177856 80180 177908 80232
rect 178408 80180 178460 80232
rect 178592 80180 178644 80232
rect 182548 80180 182600 80232
rect 238760 80180 238812 80232
rect 170726 79908 170778 79960
rect 170818 79908 170870 79960
rect 170910 79908 170962 79960
rect 171830 79908 171882 79960
rect 172198 79908 172250 79960
rect 172474 79908 172526 79960
rect 173026 79908 173078 79960
rect 170404 79772 170456 79824
rect 170634 79772 170686 79824
rect 170128 79500 170180 79552
rect 170496 79500 170548 79552
rect 170588 79500 170640 79552
rect 171278 79840 171330 79892
rect 171094 79772 171146 79824
rect 171646 79840 171698 79892
rect 171140 79568 171192 79620
rect 170956 79500 171008 79552
rect 171048 79432 171100 79484
rect 157708 79296 157760 79348
rect 158444 79296 158496 79348
rect 164976 79296 165028 79348
rect 171508 79636 171560 79688
rect 172290 79840 172342 79892
rect 172842 79840 172894 79892
rect 172934 79840 172986 79892
rect 172428 79772 172480 79824
rect 172658 79772 172710 79824
rect 173118 79840 173170 79892
rect 173210 79840 173262 79892
rect 172980 79704 173032 79756
rect 173072 79704 173124 79756
rect 173164 79704 173216 79756
rect 172060 79636 172112 79688
rect 172336 79636 172388 79688
rect 172704 79636 172756 79688
rect 172888 79636 172940 79688
rect 173394 79772 173446 79824
rect 171784 79568 171836 79620
rect 173164 79568 173216 79620
rect 173256 79568 173308 79620
rect 173348 79568 173400 79620
rect 171876 79500 171928 79552
rect 178316 80112 178368 80164
rect 185216 80112 185268 80164
rect 302240 80112 302292 80164
rect 380900 80044 380952 80096
rect 173578 79908 173630 79960
rect 172796 79432 172848 79484
rect 173440 79432 173492 79484
rect 173670 79840 173722 79892
rect 173716 79704 173768 79756
rect 178592 79976 178644 80028
rect 174038 79908 174090 79960
rect 174314 79908 174366 79960
rect 174406 79908 174458 79960
rect 174774 79908 174826 79960
rect 175050 79908 175102 79960
rect 175234 79908 175286 79960
rect 175418 79908 175470 79960
rect 175510 79908 175562 79960
rect 175786 79908 175838 79960
rect 175970 79908 176022 79960
rect 176062 79908 176114 79960
rect 177672 79908 177724 79960
rect 177856 79908 177908 79960
rect 173946 79772 173998 79824
rect 173992 79636 174044 79688
rect 174084 79568 174136 79620
rect 174590 79840 174642 79892
rect 174728 79772 174780 79824
rect 174360 79704 174412 79756
rect 174452 79704 174504 79756
rect 174544 79704 174596 79756
rect 174820 79636 174872 79688
rect 175004 79568 175056 79620
rect 174820 79500 174872 79552
rect 175188 79568 175240 79620
rect 175464 79704 175516 79756
rect 175280 79500 175332 79552
rect 175694 79840 175746 79892
rect 175740 79704 175792 79756
rect 176246 79840 176298 79892
rect 176016 79772 176068 79824
rect 176016 79636 176068 79688
rect 176522 79840 176574 79892
rect 176798 79840 176850 79892
rect 176890 79840 176942 79892
rect 177074 79840 177126 79892
rect 175648 79568 175700 79620
rect 176384 79568 176436 79620
rect 175924 79500 175976 79552
rect 176614 79772 176666 79824
rect 176568 79568 176620 79620
rect 176936 79636 176988 79688
rect 177028 79636 177080 79688
rect 177120 79568 177172 79620
rect 176108 79432 176160 79484
rect 176292 79432 176344 79484
rect 182180 79432 182232 79484
rect 171784 79364 171836 79416
rect 174176 79364 174228 79416
rect 174360 79364 174412 79416
rect 174820 79364 174872 79416
rect 175280 79364 175332 79416
rect 178132 79364 178184 79416
rect 178316 79364 178368 79416
rect 194324 79364 194376 79416
rect 172152 79296 172204 79348
rect 175096 79296 175148 79348
rect 177488 79296 177540 79348
rect 177764 79296 177816 79348
rect 196808 79296 196860 79348
rect 132408 79228 132460 79280
rect 147128 79228 147180 79280
rect 147956 79228 148008 79280
rect 122472 79160 122524 79212
rect 147680 79160 147732 79212
rect 148232 79160 148284 79212
rect 151912 79160 151964 79212
rect 152280 79160 152332 79212
rect 159548 79228 159600 79280
rect 170312 79228 170364 79280
rect 171416 79228 171468 79280
rect 171876 79228 171928 79280
rect 173164 79228 173216 79280
rect 199108 79228 199160 79280
rect 525800 79296 525852 79348
rect 170772 79160 170824 79212
rect 171600 79160 171652 79212
rect 172244 79160 172296 79212
rect 172336 79160 172388 79212
rect 198096 79160 198148 79212
rect 118792 79092 118844 79144
rect 145012 79092 145064 79144
rect 146668 79092 146720 79144
rect 118976 79024 119028 79076
rect 146300 79024 146352 79076
rect 147036 79024 147088 79076
rect 147220 79024 147272 79076
rect 150992 79092 151044 79144
rect 159548 79092 159600 79144
rect 162216 79092 162268 79144
rect 162584 79092 162636 79144
rect 164884 79092 164936 79144
rect 165620 79092 165672 79144
rect 158444 79024 158496 79076
rect 159088 79024 159140 79076
rect 159824 79024 159876 79076
rect 164976 79024 165028 79076
rect 173624 79024 173676 79076
rect 191196 79092 191248 79144
rect 174268 79024 174320 79076
rect 203708 79024 203760 79076
rect 120632 78956 120684 79008
rect 141700 78956 141752 79008
rect 119344 78888 119396 78940
rect 146300 78888 146352 78940
rect 147036 78888 147088 78940
rect 148692 78956 148744 79008
rect 161756 78956 161808 79008
rect 167460 78956 167512 79008
rect 172520 78956 172572 79008
rect 174084 78956 174136 79008
rect 174728 78956 174780 79008
rect 175096 78956 175148 79008
rect 175372 78956 175424 79008
rect 206376 78956 206428 79008
rect 149060 78888 149112 78940
rect 149980 78888 150032 78940
rect 164240 78888 164292 78940
rect 165620 78888 165672 78940
rect 171232 78888 171284 78940
rect 195428 78888 195480 78940
rect 196256 78888 196308 78940
rect 196624 78888 196676 78940
rect 483020 78888 483072 78940
rect 117872 78820 117924 78872
rect 149244 78820 149296 78872
rect 159640 78820 159692 78872
rect 191380 78820 191432 78872
rect 198740 78820 198792 78872
rect 199384 78820 199436 78872
rect 500960 78820 501012 78872
rect 132408 78752 132460 78804
rect 137744 78752 137796 78804
rect 139676 78752 139728 78804
rect 139860 78752 139912 78804
rect 141700 78752 141752 78804
rect 147772 78752 147824 78804
rect 171968 78752 172020 78804
rect 196716 78752 196768 78804
rect 196808 78752 196860 78804
rect 523132 78752 523184 78804
rect 127440 78684 127492 78736
rect 132500 78684 132552 78736
rect 133604 78684 133656 78736
rect 133880 78684 133932 78736
rect 134524 78684 134576 78736
rect 138480 78684 138532 78736
rect 144368 78684 144420 78736
rect 150624 78684 150676 78736
rect 151176 78684 151228 78736
rect 162032 78684 162084 78736
rect 102140 78616 102192 78668
rect 102876 78616 102928 78668
rect 133972 78616 134024 78668
rect 138756 78616 138808 78668
rect 139032 78616 139084 78668
rect 151268 78616 151320 78668
rect 151636 78616 151688 78668
rect 152004 78616 152056 78668
rect 153108 78616 153160 78668
rect 153936 78616 153988 78668
rect 154488 78616 154540 78668
rect 163136 78616 163188 78668
rect 163780 78616 163832 78668
rect 164332 78616 164384 78668
rect 164516 78616 164568 78668
rect 173348 78684 173400 78736
rect 196532 78684 196584 78736
rect 199108 78684 199160 78736
rect 199568 78684 199620 78736
rect 536840 78684 536892 78736
rect 104256 78548 104308 78600
rect 132592 78548 132644 78600
rect 132684 78548 132736 78600
rect 142344 78548 142396 78600
rect 170772 78548 170824 78600
rect 176292 78548 176344 78600
rect 176752 78616 176804 78668
rect 177212 78616 177264 78668
rect 177672 78548 177724 78600
rect 178776 78548 178828 78600
rect 123024 78480 123076 78532
rect 131304 78480 131356 78532
rect 132408 78480 132460 78532
rect 132500 78480 132552 78532
rect 46940 78344 46992 78396
rect 107292 78412 107344 78464
rect 136180 78412 136232 78464
rect 139768 78480 139820 78532
rect 140136 78480 140188 78532
rect 170220 78480 170272 78532
rect 196256 78480 196308 78532
rect 141884 78412 141936 78464
rect 159548 78412 159600 78464
rect 161940 78412 161992 78464
rect 162400 78412 162452 78464
rect 167184 78412 167236 78464
rect 182916 78412 182968 78464
rect 122104 78344 122156 78396
rect 149152 78344 149204 78396
rect 173256 78344 173308 78396
rect 173808 78344 173860 78396
rect 173900 78344 173952 78396
rect 174544 78344 174596 78396
rect 174728 78344 174780 78396
rect 175280 78344 175332 78396
rect 175648 78344 175700 78396
rect 176108 78344 176160 78396
rect 178500 78344 178552 78396
rect 57980 78276 58032 78328
rect 107292 78276 107344 78328
rect 122012 78276 122064 78328
rect 148324 78276 148376 78328
rect 169024 78276 169076 78328
rect 203340 78344 203392 78396
rect 287704 78344 287756 78396
rect 20720 78140 20772 78192
rect 102140 78140 102192 78192
rect 6920 78072 6972 78124
rect 106924 78208 106976 78260
rect 126980 78208 127032 78260
rect 132316 78208 132368 78260
rect 146576 78208 146628 78260
rect 179420 78208 179472 78260
rect 2872 78004 2924 78056
rect 104256 78004 104308 78056
rect 2780 77936 2832 77988
rect 108396 77936 108448 77988
rect 127164 78140 127216 78192
rect 141056 78140 141108 78192
rect 141700 78140 141752 78192
rect 142896 78140 142948 78192
rect 171876 78140 171928 78192
rect 172336 78140 172388 78192
rect 175280 78140 175332 78192
rect 176200 78140 176252 78192
rect 255964 78276 256016 78328
rect 192576 78208 192628 78260
rect 324320 78208 324372 78260
rect 337384 78140 337436 78192
rect 123208 78072 123260 78124
rect 146116 78072 146168 78124
rect 162952 78072 163004 78124
rect 393320 78072 393372 78124
rect 113640 78004 113692 78056
rect 130660 78004 130712 78056
rect 113732 77936 113784 77988
rect 123024 77936 123076 77988
rect 115112 77800 115164 77852
rect 129832 77936 129884 77988
rect 137284 78004 137336 78056
rect 139124 78004 139176 78056
rect 139400 78004 139452 78056
rect 164792 78004 164844 78056
rect 165528 78004 165580 78056
rect 169576 78004 169628 78056
rect 400864 78004 400916 78056
rect 131580 77936 131632 77988
rect 142436 77936 142488 77988
rect 163412 77936 163464 77988
rect 400220 77936 400272 77988
rect 123392 77868 123444 77920
rect 142620 77868 142672 77920
rect 142988 77868 143040 77920
rect 166632 77868 166684 77920
rect 181628 77868 181680 77920
rect 130660 77800 130712 77852
rect 132868 77800 132920 77852
rect 134156 77800 134208 77852
rect 134432 77800 134484 77852
rect 135996 77800 136048 77852
rect 136456 77800 136508 77852
rect 136824 77800 136876 77852
rect 137192 77800 137244 77852
rect 142436 77800 142488 77852
rect 143448 77800 143500 77852
rect 165804 77800 165856 77852
rect 180708 77800 180760 77852
rect 107292 77732 107344 77784
rect 136088 77732 136140 77784
rect 137836 77732 137888 77784
rect 143724 77732 143776 77784
rect 144368 77732 144420 77784
rect 153476 77732 153528 77784
rect 154396 77732 154448 77784
rect 164608 77732 164660 77784
rect 178776 77732 178828 77784
rect 132960 77664 133012 77716
rect 141700 77664 141752 77716
rect 157616 77664 157668 77716
rect 192576 77664 192628 77716
rect 131028 77596 131080 77648
rect 144920 77596 144972 77648
rect 148324 77596 148376 77648
rect 148508 77596 148560 77648
rect 164608 77596 164660 77648
rect 164884 77596 164936 77648
rect 165160 77596 165212 77648
rect 180156 77596 180208 77648
rect 176016 77528 176068 77580
rect 176384 77528 176436 77580
rect 176844 77528 176896 77580
rect 177120 77528 177172 77580
rect 140964 77460 141016 77512
rect 141332 77460 141384 77512
rect 146116 77460 146168 77512
rect 148324 77460 148376 77512
rect 162952 77460 163004 77512
rect 163320 77460 163372 77512
rect 170312 77460 170364 77512
rect 178868 77460 178920 77512
rect 173624 77392 173676 77444
rect 178040 77392 178092 77444
rect 160652 77324 160704 77376
rect 163320 77324 163372 77376
rect 151544 77256 151596 77308
rect 112628 77188 112680 77240
rect 146300 77188 146352 77240
rect 151452 77188 151504 77240
rect 163228 77256 163280 77308
rect 166264 77256 166316 77308
rect 171324 77256 171376 77308
rect 171692 77256 171744 77308
rect 172520 77256 172572 77308
rect 173348 77256 173400 77308
rect 161572 77188 161624 77240
rect 196716 77188 196768 77240
rect 72424 76780 72476 76832
rect 102784 77120 102836 77172
rect 137468 77120 137520 77172
rect 163044 77120 163096 77172
rect 197820 77120 197872 77172
rect 198188 77120 198240 77172
rect 114560 77052 114612 77104
rect 115204 77052 115256 77104
rect 115664 77052 115716 77104
rect 100760 76984 100812 77036
rect 101588 76984 101640 77036
rect 134984 76984 135036 77036
rect 135352 76984 135404 77036
rect 135628 76984 135680 77036
rect 159732 77052 159784 77104
rect 193588 77052 193640 77104
rect 148416 76984 148468 77036
rect 155500 76984 155552 77036
rect 117044 76916 117096 76968
rect 148876 76916 148928 76968
rect 155960 76916 156012 76968
rect 156880 76916 156932 76968
rect 162124 76984 162176 77036
rect 162768 76984 162820 77036
rect 191104 76984 191156 77036
rect 177764 76916 177816 76968
rect 177948 76916 178000 76968
rect 180064 76916 180116 76968
rect 188988 76916 189040 76968
rect 189172 76916 189224 76968
rect 64144 76712 64196 76764
rect 105728 76848 105780 76900
rect 136916 76848 136968 76900
rect 145288 76848 145340 76900
rect 146208 76848 146260 76900
rect 151084 76848 151136 76900
rect 211804 76848 211856 76900
rect 119712 76780 119764 76832
rect 151452 76780 151504 76832
rect 224224 76780 224276 76832
rect 111340 76712 111392 76764
rect 141056 76712 141108 76764
rect 141424 76712 141476 76764
rect 143172 76712 143224 76764
rect 143448 76712 143500 76764
rect 149152 76712 149204 76764
rect 149796 76712 149848 76764
rect 152648 76712 152700 76764
rect 260840 76712 260892 76764
rect 34520 76644 34572 76696
rect 100760 76644 100812 76696
rect 115204 76644 115256 76696
rect 127164 76644 127216 76696
rect 153200 76644 153252 76696
rect 153476 76644 153528 76696
rect 155224 76644 155276 76696
rect 171784 76644 171836 76696
rect 52460 76576 52512 76628
rect 135352 76576 135404 76628
rect 149520 76576 149572 76628
rect 149980 76576 150032 76628
rect 168472 76576 168524 76628
rect 169300 76576 169352 76628
rect 35900 76508 35952 76560
rect 134248 76508 134300 76560
rect 147128 76508 147180 76560
rect 181444 76644 181496 76696
rect 193588 76644 193640 76696
rect 194048 76644 194100 76696
rect 353300 76644 353352 76696
rect 112536 76440 112588 76492
rect 138296 76440 138348 76492
rect 170864 76440 170916 76492
rect 187700 76576 187752 76628
rect 196716 76576 196768 76628
rect 374000 76576 374052 76628
rect 174544 76508 174596 76560
rect 174728 76508 174780 76560
rect 170680 76372 170732 76424
rect 186688 76508 186740 76560
rect 197820 76508 197872 76560
rect 391940 76508 391992 76560
rect 131856 76304 131908 76356
rect 140596 76304 140648 76356
rect 145472 76304 145524 76356
rect 145932 76304 145984 76356
rect 170772 76304 170824 76356
rect 187332 76372 187384 76424
rect 180708 76304 180760 76356
rect 200764 76304 200816 76356
rect 177028 76168 177080 76220
rect 177948 76168 178000 76220
rect 170128 76100 170180 76152
rect 170680 76100 170732 76152
rect 124864 76032 124916 76084
rect 125600 76032 125652 76084
rect 171232 76032 171284 76084
rect 171600 76032 171652 76084
rect 172796 76032 172848 76084
rect 177212 76032 177264 76084
rect 171784 75964 171836 76016
rect 179880 75964 179932 76016
rect 289820 75964 289872 76016
rect 167920 75896 167972 75948
rect 168288 75896 168340 75948
rect 168932 75896 168984 75948
rect 169576 75896 169628 75948
rect 169852 75896 169904 75948
rect 170588 75896 170640 75948
rect 177764 75896 177816 75948
rect 181352 75896 181404 75948
rect 296720 75896 296772 75948
rect 111524 75828 111576 75880
rect 145472 75828 145524 75880
rect 167552 75828 167604 75880
rect 202328 75828 202380 75880
rect 115388 75760 115440 75812
rect 96620 75692 96672 75744
rect 105820 75692 105872 75744
rect 139676 75692 139728 75744
rect 130752 75624 130804 75676
rect 131028 75624 131080 75676
rect 134248 75624 134300 75676
rect 134708 75624 134760 75676
rect 135444 75624 135496 75676
rect 136456 75624 136508 75676
rect 107016 75556 107068 75608
rect 139124 75556 139176 75608
rect 156420 75760 156472 75812
rect 156880 75760 156932 75812
rect 161664 75760 161716 75812
rect 162768 75760 162820 75812
rect 196348 75760 196400 75812
rect 146300 75692 146352 75744
rect 180800 75692 180852 75744
rect 146760 75624 146812 75676
rect 185032 75624 185084 75676
rect 117228 75488 117280 75540
rect 145380 75488 145432 75540
rect 147864 75556 147916 75608
rect 198740 75556 198792 75608
rect 121184 75420 121236 75472
rect 148140 75420 148192 75472
rect 150164 75488 150216 75540
rect 216680 75488 216732 75540
rect 149612 75420 149664 75472
rect 223580 75420 223632 75472
rect 122748 75352 122800 75404
rect 149888 75352 149940 75404
rect 165712 75352 165764 75404
rect 165988 75352 166040 75404
rect 167552 75352 167604 75404
rect 168012 75352 168064 75404
rect 171508 75352 171560 75404
rect 118608 75284 118660 75336
rect 145564 75284 145616 75336
rect 156052 75284 156104 75336
rect 156788 75284 156840 75336
rect 160468 75284 160520 75336
rect 162032 75284 162084 75336
rect 166080 75284 166132 75336
rect 171968 75284 172020 75336
rect 174176 75352 174228 75404
rect 504364 75352 504416 75404
rect 454684 75284 454736 75336
rect 81440 75216 81492 75268
rect 138664 75216 138716 75268
rect 145380 75216 145432 75268
rect 145748 75216 145800 75268
rect 167000 75216 167052 75268
rect 168104 75216 168156 75268
rect 172888 75216 172940 75268
rect 173716 75216 173768 75268
rect 174360 75216 174412 75268
rect 511264 75216 511316 75268
rect 67640 75148 67692 75200
rect 132592 75148 132644 75200
rect 132684 75148 132736 75200
rect 133788 75148 133840 75200
rect 135812 75148 135864 75200
rect 136548 75148 136600 75200
rect 136640 75148 136692 75200
rect 137192 75148 137244 75200
rect 168656 75148 168708 75200
rect 169116 75148 169168 75200
rect 172980 75148 173032 75200
rect 521660 75148 521712 75200
rect 115940 75080 115992 75132
rect 116492 75080 116544 75132
rect 141332 75080 141384 75132
rect 157524 75080 157576 75132
rect 189908 75080 189960 75132
rect 114468 75012 114520 75064
rect 147220 75012 147272 75064
rect 159824 75012 159876 75064
rect 160008 75012 160060 75064
rect 164792 75012 164844 75064
rect 192484 75012 192536 75064
rect 134340 74944 134392 74996
rect 135168 74944 135220 74996
rect 135444 74944 135496 74996
rect 136272 74944 136324 74996
rect 173716 74944 173768 74996
rect 198372 74944 198424 74996
rect 132592 74876 132644 74928
rect 137652 74876 137704 74928
rect 158812 74876 158864 74928
rect 159824 74876 159876 74928
rect 176844 74876 176896 74928
rect 177764 74876 177816 74928
rect 129924 74672 129976 74724
rect 142160 74672 142212 74724
rect 158904 74604 158956 74656
rect 159456 74604 159508 74656
rect 168564 74604 168616 74656
rect 169208 74604 169260 74656
rect 111156 74468 111208 74520
rect 143540 74468 143592 74520
rect 143724 74468 143776 74520
rect 144092 74468 144144 74520
rect 145012 74468 145064 74520
rect 145380 74468 145432 74520
rect 161020 74468 161072 74520
rect 161480 74468 161532 74520
rect 165896 74468 165948 74520
rect 166816 74468 166868 74520
rect 200856 74468 200908 74520
rect 111708 74400 111760 74452
rect 144276 74400 144328 74452
rect 168748 74400 168800 74452
rect 202052 74400 202104 74452
rect 120356 74332 120408 74384
rect 152096 74332 152148 74384
rect 160560 74332 160612 74384
rect 161296 74332 161348 74384
rect 193864 74332 193916 74384
rect 108304 74264 108356 74316
rect 140688 74264 140740 74316
rect 150256 74264 150308 74316
rect 203616 74264 203668 74316
rect 114100 74196 114152 74248
rect 145012 74196 145064 74248
rect 150900 74196 150952 74248
rect 237380 74196 237432 74248
rect 112720 74128 112772 74180
rect 143724 74128 143776 74180
rect 151728 74128 151780 74180
rect 247684 74128 247736 74180
rect 117964 74060 118016 74112
rect 148048 74060 148100 74112
rect 154212 74060 154264 74112
rect 284300 74060 284352 74112
rect 112996 73992 113048 74044
rect 142436 73992 142488 74044
rect 157524 73992 157576 74044
rect 158260 73992 158312 74044
rect 159364 73992 159416 74044
rect 347780 73992 347832 74044
rect 113456 73924 113508 73976
rect 138572 73924 138624 73976
rect 141608 73924 141660 73976
rect 141976 73924 142028 73976
rect 152188 73924 152240 73976
rect 255320 73924 255372 73976
rect 255964 73924 256016 73976
rect 456800 73924 456852 73976
rect 95240 73856 95292 73908
rect 140044 73856 140096 73908
rect 157340 73856 157392 73908
rect 158352 73856 158404 73908
rect 172428 73856 172480 73908
rect 190184 73856 190236 73908
rect 202052 73856 202104 73908
rect 446404 73856 446456 73908
rect 54484 73788 54536 73840
rect 107384 73788 107436 73840
rect 115204 73788 115256 73840
rect 138388 73788 138440 73840
rect 143540 73788 143592 73840
rect 144184 73788 144236 73840
rect 152188 73788 152240 73840
rect 152924 73788 152976 73840
rect 261484 73788 261536 73840
rect 264244 73788 264296 73840
rect 518900 73788 518952 73840
rect 117688 73720 117740 73772
rect 129740 73720 129792 73772
rect 132960 73720 133012 73772
rect 176200 73720 176252 73772
rect 204628 73720 204680 73772
rect 169392 73652 169444 73704
rect 180248 73652 180300 73704
rect 107384 73584 107436 73636
rect 136364 73584 136416 73636
rect 158996 73244 159048 73296
rect 159180 73244 159232 73296
rect 107660 73176 107712 73228
rect 108304 73176 108356 73228
rect 124956 73176 125008 73228
rect 125692 73176 125744 73228
rect 105912 73108 105964 73160
rect 139584 73108 139636 73160
rect 140504 73108 140556 73160
rect 114284 73040 114336 73092
rect 146668 73108 146720 73160
rect 164700 73108 164752 73160
rect 165252 73108 165304 73160
rect 199476 73108 199528 73160
rect 327724 73108 327776 73160
rect 579988 73108 580040 73160
rect 142252 73040 142304 73092
rect 143448 73040 143500 73092
rect 157064 73040 157116 73092
rect 191012 73040 191064 73092
rect 121276 72972 121328 73024
rect 100208 72904 100260 72956
rect 133604 72904 133656 72956
rect 153752 72972 153804 73024
rect 156512 72972 156564 73024
rect 187056 72972 187108 73024
rect 187608 72972 187660 73024
rect 154856 72904 154908 72956
rect 242164 72904 242216 72956
rect 122656 72836 122708 72888
rect 154028 72836 154080 72888
rect 160100 72836 160152 72888
rect 160744 72836 160796 72888
rect 189816 72836 189868 72888
rect 191012 72836 191064 72888
rect 301504 72836 301556 72888
rect 104348 72768 104400 72820
rect 135260 72768 135312 72820
rect 187608 72768 187660 72820
rect 305000 72768 305052 72820
rect 111432 72700 111484 72752
rect 142896 72700 142948 72752
rect 156972 72700 157024 72752
rect 311164 72700 311216 72752
rect 111616 72632 111668 72684
rect 142252 72632 142304 72684
rect 157432 72632 157484 72684
rect 318800 72632 318852 72684
rect 70400 72564 70452 72616
rect 137928 72564 137980 72616
rect 153292 72564 153344 72616
rect 153660 72564 153712 72616
rect 157708 72564 157760 72616
rect 324964 72564 325016 72616
rect 21364 72496 21416 72548
rect 100208 72496 100260 72548
rect 112904 72496 112956 72548
rect 142528 72496 142580 72548
rect 157800 72496 157852 72548
rect 332600 72496 332652 72548
rect 45560 72428 45612 72480
rect 135536 72428 135588 72480
rect 145656 72428 145708 72480
rect 156328 72428 156380 72480
rect 167460 72428 167512 72480
rect 375380 72428 375432 72480
rect 119804 72360 119856 72412
rect 141516 72360 141568 72412
rect 146668 72360 146720 72412
rect 147404 72360 147456 72412
rect 162216 72360 162268 72412
rect 190092 72360 190144 72412
rect 121368 72292 121420 72344
rect 129924 72292 129976 72344
rect 135260 72292 135312 72344
rect 135536 72292 135588 72344
rect 160008 72292 160060 72344
rect 187240 72292 187292 72344
rect 174912 72224 174964 72276
rect 205916 72224 205968 72276
rect 164240 72156 164292 72208
rect 165528 72156 165580 72208
rect 195520 72156 195572 72208
rect 148048 72088 148100 72140
rect 148784 72088 148836 72140
rect 152096 72088 152148 72140
rect 152832 72088 152884 72140
rect 164240 72020 164292 72072
rect 164608 72020 164660 72072
rect 161848 71952 161900 72004
rect 162400 71952 162452 72004
rect 166356 71816 166408 71868
rect 166908 71816 166960 71868
rect 118700 71748 118752 71800
rect 119804 71748 119856 71800
rect 163964 71748 164016 71800
rect 117596 71680 117648 71732
rect 151820 71680 151872 71732
rect 164332 71680 164384 71732
rect 165436 71680 165488 71732
rect 165988 71680 166040 71732
rect 166356 71680 166408 71732
rect 3516 71612 3568 71664
rect 8944 71612 8996 71664
rect 120816 71612 120868 71664
rect 154580 71612 154632 71664
rect 155224 71612 155276 71664
rect 182180 71680 182232 71732
rect 192116 71680 192168 71732
rect 198004 71612 198056 71664
rect 100116 71544 100168 71596
rect 134616 71544 134668 71596
rect 138572 71544 138624 71596
rect 139308 71544 139360 71596
rect 141516 71544 141568 71596
rect 142896 71544 142948 71596
rect 165160 71544 165212 71596
rect 165620 71544 165672 71596
rect 199292 71544 199344 71596
rect 118148 71476 118200 71528
rect 150808 71476 150860 71528
rect 120448 71408 120500 71460
rect 104440 71340 104492 71392
rect 134156 71340 134208 71392
rect 134800 71340 134852 71392
rect 142344 71408 142396 71460
rect 143172 71408 143224 71460
rect 151820 71408 151872 71460
rect 152740 71408 152792 71460
rect 163688 71408 163740 71460
rect 163964 71408 164016 71460
rect 196992 71476 197044 71528
rect 153568 71340 153620 71392
rect 161020 71340 161072 71392
rect 192300 71408 192352 71460
rect 169484 71340 169536 71392
rect 196440 71340 196492 71392
rect 108580 71272 108632 71324
rect 121460 71272 121512 71324
rect 123116 71272 123168 71324
rect 152556 71272 152608 71324
rect 161388 71272 161440 71324
rect 187148 71272 187200 71324
rect 108856 71204 108908 71256
rect 138388 71204 138440 71256
rect 139032 71204 139084 71256
rect 162400 71204 162452 71256
rect 188344 71204 188396 71256
rect 113364 71136 113416 71188
rect 142344 71136 142396 71188
rect 153568 71136 153620 71188
rect 153936 71136 153988 71188
rect 165436 71136 165488 71188
rect 186964 71136 187016 71188
rect 115296 71068 115348 71120
rect 138572 71068 138624 71120
rect 148876 71068 148928 71120
rect 27620 71000 27672 71052
rect 100116 71000 100168 71052
rect 102784 71000 102836 71052
rect 106832 71000 106884 71052
rect 116124 71000 116176 71052
rect 136916 71000 136968 71052
rect 142804 71000 142856 71052
rect 153568 71000 153620 71052
rect 154120 71000 154172 71052
rect 184204 71000 184256 71052
rect 192116 71000 192168 71052
rect 192852 71000 192904 71052
rect 200120 71000 200172 71052
rect 121460 70932 121512 70984
rect 142068 70932 142120 70984
rect 142436 70864 142488 70916
rect 142804 70864 142856 70916
rect 150808 70864 150860 70916
rect 151268 70864 151320 70916
rect 166356 70864 166408 70916
rect 200028 70864 200080 70916
rect 187608 70456 187660 70508
rect 480260 70456 480312 70508
rect 190368 70388 190420 70440
rect 531320 70388 531372 70440
rect 116768 70320 116820 70372
rect 151084 70320 151136 70372
rect 168104 70320 168156 70372
rect 202236 70320 202288 70372
rect 121000 70252 121052 70304
rect 154672 70252 154724 70304
rect 155408 70252 155460 70304
rect 166540 70252 166592 70304
rect 166724 70252 166776 70304
rect 169576 70252 169628 70304
rect 203524 70252 203576 70304
rect 117504 70184 117556 70236
rect 152280 70184 152332 70236
rect 152556 70184 152608 70236
rect 168288 70184 168340 70236
rect 198280 70184 198332 70236
rect 106004 70116 106056 70168
rect 140228 70116 140280 70168
rect 165896 70116 165948 70168
rect 166724 70116 166776 70168
rect 194140 70116 194192 70168
rect 122196 70048 122248 70100
rect 154948 70048 155000 70100
rect 155316 70048 155368 70100
rect 166908 70048 166960 70100
rect 192576 70048 192628 70100
rect 102140 69980 102192 70032
rect 102968 69980 103020 70032
rect 136548 69980 136600 70032
rect 171968 69980 172020 70032
rect 192760 69980 192812 70032
rect 103520 69912 103572 69964
rect 106004 69912 106056 69964
rect 110236 69912 110288 69964
rect 142620 69912 142672 69964
rect 175832 69912 175884 69964
rect 199568 69912 199620 69964
rect 89720 69844 89772 69896
rect 107016 69844 107068 69896
rect 110328 69844 110380 69896
rect 142436 69844 142488 69896
rect 142712 69844 142764 69896
rect 147036 69844 147088 69896
rect 179420 69844 179472 69896
rect 46204 69776 46256 69828
rect 103336 69776 103388 69828
rect 134708 69776 134760 69828
rect 147864 69776 147916 69828
rect 196624 69776 196676 69828
rect 41420 69708 41472 69760
rect 102140 69708 102192 69760
rect 122564 69708 122616 69760
rect 153292 69708 153344 69760
rect 153844 69708 153896 69760
rect 160192 69708 160244 69760
rect 354680 69708 354732 69760
rect 18604 69640 18656 69692
rect 103428 69640 103480 69692
rect 113548 69640 113600 69692
rect 142160 69640 142212 69692
rect 142988 69640 143040 69692
rect 143724 69640 143776 69692
rect 147036 69640 147088 69692
rect 147220 69640 147272 69692
rect 182824 69640 182876 69692
rect 192760 69640 192812 69692
rect 430580 69640 430632 69692
rect 116308 69572 116360 69624
rect 128452 69572 128504 69624
rect 141608 69572 141660 69624
rect 166540 69572 166592 69624
rect 188436 69572 188488 69624
rect 133696 69504 133748 69556
rect 199568 69028 199620 69080
rect 561680 69028 561732 69080
rect 109040 68960 109092 69012
rect 110972 68960 111024 69012
rect 104532 68892 104584 68944
rect 104808 68892 104860 68944
rect 135444 68960 135496 69012
rect 145380 68960 145432 69012
rect 147128 68960 147180 69012
rect 164332 68960 164384 69012
rect 199108 68960 199160 69012
rect 199660 68960 199712 69012
rect 161480 68892 161532 68944
rect 195244 68892 195296 68944
rect 180340 68824 180392 68876
rect 182180 68824 182232 68876
rect 176752 68756 176804 68808
rect 196256 68824 196308 68876
rect 195244 68416 195296 68468
rect 367100 68416 367152 68468
rect 199108 68348 199160 68400
rect 412640 68348 412692 68400
rect 48320 68280 48372 68332
rect 104808 68280 104860 68332
rect 167736 68280 167788 68332
rect 453304 68280 453356 68332
rect 196256 67600 196308 67652
rect 574744 67600 574796 67652
rect 110052 67532 110104 67584
rect 144000 67532 144052 67584
rect 155132 67532 155184 67584
rect 189264 67532 189316 67584
rect 108948 67464 109000 67516
rect 135444 67464 135496 67516
rect 135812 67464 135864 67516
rect 163044 67464 163096 67516
rect 195152 67464 195204 67516
rect 175648 67396 175700 67448
rect 200856 67396 200908 67448
rect 201408 67396 201460 67448
rect 78680 67056 78732 67108
rect 108488 67056 108540 67108
rect 120080 67056 120132 67108
rect 141976 67056 142028 67108
rect 75920 66988 75972 67040
rect 107108 66988 107160 67040
rect 113180 66988 113232 67040
rect 141056 66988 141108 67040
rect 150624 66988 150676 67040
rect 242900 66988 242952 67040
rect 80060 66920 80112 66972
rect 113456 66920 113508 66972
rect 117320 66920 117372 66972
rect 140964 66920 141016 66972
rect 189264 66920 189316 66972
rect 295340 66920 295392 66972
rect 60740 66852 60792 66904
rect 137284 66852 137336 66904
rect 195152 66852 195204 66904
rect 402980 66852 403032 66904
rect 140780 66240 140832 66292
rect 142160 66240 142212 66292
rect 201408 66240 201460 66292
rect 557540 66240 557592 66292
rect 102140 66172 102192 66224
rect 103244 66172 103296 66224
rect 137192 66172 137244 66224
rect 144368 66172 144420 66224
rect 147220 66172 147272 66224
rect 159180 66172 159232 66224
rect 192024 66172 192076 66224
rect 193128 66172 193180 66224
rect 109132 66104 109184 66156
rect 109960 66104 110012 66156
rect 139952 66104 140004 66156
rect 173164 66104 173216 66156
rect 194048 66104 194100 66156
rect 194508 66104 194560 66156
rect 104808 66036 104860 66088
rect 134340 66036 134392 66088
rect 98000 65696 98052 65748
rect 109132 65696 109184 65748
rect 93124 65628 93176 65680
rect 116584 65968 116636 66020
rect 139860 65968 139912 66020
rect 148416 65628 148468 65680
rect 207020 65628 207072 65680
rect 57244 65560 57296 65612
rect 102140 65560 102192 65612
rect 153752 65560 153804 65612
rect 274640 65560 274692 65612
rect 35992 65492 36044 65544
rect 104808 65492 104860 65544
rect 146392 65492 146444 65544
rect 183560 65492 183612 65544
rect 193128 65492 193180 65544
rect 346400 65492 346452 65544
rect 139400 64880 139452 64932
rect 142252 64948 142304 65000
rect 194508 64880 194560 64932
rect 529940 64880 529992 64932
rect 106188 64812 106240 64864
rect 137100 64812 137152 64864
rect 160192 64812 160244 64864
rect 194876 64812 194928 64864
rect 168656 64744 168708 64796
rect 203248 64744 203300 64796
rect 149888 64268 149940 64320
rect 224960 64268 225012 64320
rect 62120 64200 62172 64252
rect 106188 64200 106240 64252
rect 194876 64200 194928 64252
rect 358820 64200 358872 64252
rect 4160 64132 4212 64184
rect 133420 64132 133472 64184
rect 147404 64132 147456 64184
rect 187700 64132 187752 64184
rect 203248 64132 203300 64184
rect 472624 64132 472676 64184
rect 104624 63452 104676 63504
rect 132776 63452 132828 63504
rect 159088 63452 159140 63504
rect 193496 63452 193548 63504
rect 75184 62908 75236 62960
rect 104164 62908 104216 62960
rect 88340 62840 88392 62892
rect 139216 62840 139268 62892
rect 178868 62840 178920 62892
rect 227720 62840 227772 62892
rect 10324 62772 10376 62824
rect 104624 62772 104676 62824
rect 193496 62772 193548 62824
rect 340880 62772 340932 62824
rect 197452 62160 197504 62212
rect 197728 62160 197780 62212
rect 104532 62024 104584 62076
rect 104716 62024 104768 62076
rect 135996 62024 136048 62076
rect 162952 62024 163004 62076
rect 197452 62024 197504 62076
rect 197636 62024 197688 62076
rect 167184 61956 167236 62008
rect 199016 61956 199068 62008
rect 52552 61412 52604 61464
rect 104532 61412 104584 61464
rect 197452 61412 197504 61464
rect 394700 61412 394752 61464
rect 42800 61344 42852 61396
rect 135720 61344 135772 61396
rect 199016 61344 199068 61396
rect 459560 61344 459612 61396
rect 135260 61208 135312 61260
rect 142528 61208 142580 61260
rect 99380 60664 99432 60716
rect 100392 60664 100444 60716
rect 134432 60664 134484 60716
rect 162860 60664 162912 60716
rect 197452 60664 197504 60716
rect 197728 60664 197780 60716
rect 99472 60596 99524 60648
rect 100576 60596 100628 60648
rect 132684 60596 132736 60648
rect 166264 60596 166316 60648
rect 194232 60596 194284 60648
rect 194508 60596 194560 60648
rect 107476 60528 107528 60580
rect 137376 60528 137428 60580
rect 69020 60120 69072 60172
rect 107476 60120 107528 60172
rect 23480 60052 23532 60104
rect 99380 60052 99432 60104
rect 197452 60052 197504 60104
rect 398840 60052 398892 60104
rect 17960 59984 18012 60036
rect 99472 59984 99524 60036
rect 147312 59984 147364 60036
rect 186320 59984 186372 60036
rect 194508 59984 194560 60036
rect 396080 59984 396132 60036
rect 110512 59304 110564 59356
rect 114928 59304 114980 59356
rect 144276 59304 144328 59356
rect 148416 59304 148468 59356
rect 167092 59304 167144 59356
rect 201960 59304 202012 59356
rect 202788 59304 202840 59356
rect 148968 58760 149020 58812
rect 209872 58760 209924 58812
rect 202788 58692 202840 58744
rect 448520 58692 448572 58744
rect 169944 58624 169996 58676
rect 489920 58624 489972 58676
rect 168564 57876 168616 57928
rect 203432 57876 203484 57928
rect 204168 57876 204220 57928
rect 158996 57808 159048 57860
rect 193312 57808 193364 57860
rect 194508 57808 194560 57860
rect 151268 57332 151320 57384
rect 236000 57332 236052 57384
rect 194508 57264 194560 57316
rect 345020 57264 345072 57316
rect 77392 57196 77444 57248
rect 112536 57196 112588 57248
rect 147772 57196 147824 57248
rect 197452 57196 197504 57248
rect 204168 57196 204220 57248
rect 473452 57196 473504 57248
rect 99380 56516 99432 56568
rect 100668 56516 100720 56568
rect 133604 56516 133656 56568
rect 167828 56516 167880 56568
rect 201868 56516 201920 56568
rect 202788 56516 202840 56568
rect 158904 56448 158956 56500
rect 193404 56448 193456 56500
rect 194508 56448 194560 56500
rect 176936 56380 176988 56432
rect 200672 56380 200724 56432
rect 201408 56380 201460 56432
rect 63500 55904 63552 55956
rect 136824 55904 136876 55956
rect 194508 55904 194560 55956
rect 349160 55904 349212 55956
rect 12440 55836 12492 55888
rect 99380 55836 99432 55888
rect 145748 55836 145800 55888
rect 162124 55836 162176 55888
rect 202788 55836 202840 55888
rect 450544 55836 450596 55888
rect 138664 55224 138716 55276
rect 142252 55224 142304 55276
rect 201408 55224 201460 55276
rect 560944 55224 560996 55276
rect 169024 55156 169076 55208
rect 203064 55156 203116 55208
rect 152832 54612 152884 54664
rect 253940 54612 253992 54664
rect 84200 54544 84252 54596
rect 115204 54544 115256 54596
rect 158076 54544 158128 54596
rect 333980 54544 334032 54596
rect 99380 54476 99432 54528
rect 139768 54476 139820 54528
rect 203064 54476 203116 54528
rect 468484 54476 468536 54528
rect 100484 53728 100536 53780
rect 133052 53728 133104 53780
rect 147680 53116 147732 53168
rect 204260 53116 204312 53168
rect 9680 53048 9732 53100
rect 100484 53048 100536 53100
rect 176108 53048 176160 53100
rect 556160 53048 556212 53100
rect 143816 52844 143868 52896
rect 148508 52844 148560 52896
rect 168380 52368 168432 52420
rect 201500 52368 201552 52420
rect 202788 52368 202840 52420
rect 149796 51824 149848 51876
rect 215300 51824 215352 51876
rect 202788 51756 202840 51808
rect 464344 51756 464396 51808
rect 176660 51688 176712 51740
rect 578240 51688 578292 51740
rect 100760 51008 100812 51060
rect 101864 51008 101916 51060
rect 134248 51008 134300 51060
rect 93952 50396 94004 50448
rect 105544 50396 105596 50448
rect 30380 50328 30432 50380
rect 100760 50328 100812 50380
rect 155592 50328 155644 50380
rect 293960 50328 294012 50380
rect 148784 49104 148836 49156
rect 201500 49104 201552 49156
rect 149980 49036 150032 49088
rect 218152 49036 218204 49088
rect 170680 48968 170732 49020
rect 486424 48968 486476 49020
rect 149244 47676 149296 47728
rect 222200 47676 222252 47728
rect 151912 47608 151964 47660
rect 267740 47608 267792 47660
rect 144184 47540 144236 47592
rect 149244 47540 149296 47592
rect 173900 47540 173952 47592
rect 542360 47540 542412 47592
rect 155408 46316 155460 46368
rect 285680 46316 285732 46368
rect 165068 46248 165120 46300
rect 418160 46248 418212 46300
rect 145196 46180 145248 46232
rect 168380 46180 168432 46232
rect 169208 46180 169260 46232
rect 463700 46180 463752 46232
rect 148692 44888 148744 44940
rect 201592 44888 201644 44940
rect 60832 44820 60884 44872
rect 136640 44820 136692 44872
rect 154304 44820 154356 44872
rect 273260 44820 273312 44872
rect 146116 43596 146168 43648
rect 167000 43596 167052 43648
rect 151176 43528 151228 43580
rect 233240 43528 233292 43580
rect 162032 43460 162084 43512
rect 361580 43460 361632 43512
rect 74540 43392 74592 43444
rect 112444 43392 112496 43444
rect 164884 43392 164936 43444
rect 426440 43392 426492 43444
rect 155316 42236 155368 42288
rect 292672 42236 292724 42288
rect 156972 42168 157024 42220
rect 307852 42168 307904 42220
rect 171508 42100 171560 42152
rect 498292 42100 498344 42152
rect 174820 42032 174872 42084
rect 538864 42032 538916 42084
rect 138020 41624 138072 41676
rect 142620 41624 142672 41676
rect 154396 40944 154448 40996
rect 276020 40944 276072 40996
rect 158260 40876 158312 40928
rect 322940 40876 322992 40928
rect 166356 40808 166408 40860
rect 427820 40808 427872 40860
rect 173440 40740 173492 40792
rect 516140 40740 516192 40792
rect 13820 40672 13872 40724
rect 132868 40672 132920 40724
rect 177304 40672 177356 40724
rect 554780 40672 554832 40724
rect 144460 39992 144512 40044
rect 145104 39992 145156 40044
rect 152740 39584 152792 39636
rect 251180 39584 251232 39636
rect 160652 39516 160704 39568
rect 357532 39516 357584 39568
rect 169484 39448 169536 39500
rect 477500 39448 477552 39500
rect 170772 39380 170824 39432
rect 484400 39380 484452 39432
rect 31760 39312 31812 39364
rect 133880 39312 133932 39364
rect 145656 39312 145708 39364
rect 168472 39312 168524 39364
rect 174728 39312 174780 39364
rect 534080 39312 534132 39364
rect 154212 38156 154264 38208
rect 267832 38156 267884 38208
rect 164976 38088 165028 38140
rect 368480 38088 368532 38140
rect 170036 38020 170088 38072
rect 488540 38020 488592 38072
rect 173532 37952 173584 38004
rect 527824 37952 527876 38004
rect 38660 37884 38712 37936
rect 135628 37884 135680 37936
rect 175372 37884 175424 37936
rect 552020 37884 552072 37936
rect 135352 37272 135404 37324
rect 142436 37272 142488 37324
rect 147496 36864 147548 36916
rect 191840 36864 191892 36916
rect 148600 36796 148652 36848
rect 205640 36796 205692 36848
rect 156788 36728 156840 36780
rect 303620 36728 303672 36780
rect 170864 36660 170916 36712
rect 490012 36660 490064 36712
rect 171416 36592 171468 36644
rect 502340 36592 502392 36644
rect 145564 36524 145616 36576
rect 170404 36524 170456 36576
rect 176200 36524 176252 36576
rect 558920 36524 558972 36576
rect 152004 35368 152056 35420
rect 266360 35368 266412 35420
rect 158352 35300 158404 35352
rect 321560 35300 321612 35352
rect 169852 35232 169904 35284
rect 491300 35232 491352 35284
rect 53840 35164 53892 35216
rect 135444 35164 135496 35216
rect 177396 35164 177448 35216
rect 576216 35164 576268 35216
rect 155684 34008 155736 34060
rect 299572 34008 299624 34060
rect 163412 33940 163464 33992
rect 340972 33940 341024 33992
rect 162216 33872 162268 33924
rect 385040 33872 385092 33924
rect 167920 33804 167972 33856
rect 460940 33804 460992 33856
rect 170496 33736 170548 33788
rect 495440 33736 495492 33788
rect 147588 32648 147640 32700
rect 194600 32648 194652 32700
rect 154120 32580 154172 32632
rect 278780 32580 278832 32632
rect 160928 32512 160980 32564
rect 356704 32512 356756 32564
rect 166448 32444 166500 32496
rect 431960 32444 432012 32496
rect 172612 32376 172664 32428
rect 531412 32376 531464 32428
rect 157156 31288 157208 31340
rect 317420 31288 317472 31340
rect 159916 31220 159968 31272
rect 350540 31220 350592 31272
rect 164240 31152 164292 31204
rect 420920 31152 420972 31204
rect 169668 31084 169720 31136
rect 474740 31084 474792 31136
rect 44272 31016 44324 31068
rect 135536 31016 135588 31068
rect 177672 31016 177724 31068
rect 571984 31016 572036 31068
rect 158444 29792 158496 29844
rect 332692 29792 332744 29844
rect 162308 29724 162360 29776
rect 378784 29724 378836 29776
rect 168012 29656 168064 29708
rect 452660 29656 452712 29708
rect 171324 29588 171376 29640
rect 506572 29588 506624 29640
rect 152648 28500 152700 28552
rect 258080 28500 258132 28552
rect 159824 28432 159876 28484
rect 339500 28432 339552 28484
rect 163872 28364 163924 28416
rect 397460 28364 397512 28416
rect 169576 28296 169628 28348
rect 470600 28296 470652 28348
rect 171232 28228 171284 28280
rect 509240 28228 509292 28280
rect 165160 27072 165212 27124
rect 409880 27072 409932 27124
rect 180708 27004 180760 27056
rect 429200 27004 429252 27056
rect 171876 26936 171928 26988
rect 513380 26936 513432 26988
rect 174912 26868 174964 26920
rect 535460 26868 535512 26920
rect 156696 25780 156748 25832
rect 310520 25780 310572 25832
rect 181628 25712 181680 25764
rect 436100 25712 436152 25764
rect 173716 25644 173768 25696
rect 520280 25644 520332 25696
rect 175004 25576 175056 25628
rect 546500 25576 546552 25628
rect 145012 25508 145064 25560
rect 171784 25508 171836 25560
rect 177764 25508 177816 25560
rect 571340 25508 571392 25560
rect 154028 24352 154080 24404
rect 284392 24352 284444 24404
rect 157340 24284 157392 24336
rect 328460 24284 328512 24336
rect 168196 24216 168248 24268
rect 449900 24216 449952 24268
rect 172520 24148 172572 24200
rect 527180 24148 527232 24200
rect 176292 24080 176344 24132
rect 564532 24080 564584 24132
rect 150072 22992 150124 23044
rect 219440 22992 219492 23044
rect 161112 22924 161164 22976
rect 365812 22924 365864 22976
rect 165252 22856 165304 22908
rect 416780 22856 416832 22908
rect 173992 22788 174044 22840
rect 538220 22788 538272 22840
rect 177856 22720 177908 22772
rect 580264 22720 580316 22772
rect 158536 21632 158588 21684
rect 329104 21632 329156 21684
rect 158168 21564 158220 21616
rect 336740 21564 336792 21616
rect 337384 21564 337436 21616
rect 471980 21564 472032 21616
rect 158812 21496 158864 21548
rect 342904 21496 342956 21548
rect 178776 21428 178828 21480
rect 415492 21428 415544 21480
rect 166632 21360 166684 21412
rect 440332 21360 440384 21412
rect 3424 20612 3476 20664
rect 187884 20612 187936 20664
rect 485044 20612 485096 20664
rect 579988 20612 580040 20664
rect 154488 20204 154540 20256
rect 280160 20204 280212 20256
rect 155776 20136 155828 20188
rect 291200 20136 291252 20188
rect 155224 20068 155276 20120
rect 287060 20068 287112 20120
rect 287704 20068 287756 20120
rect 465172 20068 465224 20120
rect 161204 20000 161256 20052
rect 372620 20000 372672 20052
rect 143632 19932 143684 19984
rect 154580 19932 154632 19984
rect 182916 19932 182968 19984
rect 443000 19932 443052 19984
rect 149060 18844 149112 18896
rect 226340 18844 226392 18896
rect 155868 18776 155920 18828
rect 300860 18776 300912 18828
rect 176384 18708 176436 18760
rect 529204 18708 529256 18760
rect 175924 18640 175976 18692
rect 567200 18640 567252 18692
rect 177948 18572 178000 18624
rect 574100 18572 574152 18624
rect 151636 17484 151688 17536
rect 241520 17484 241572 17536
rect 165344 17416 165396 17468
rect 425060 17416 425112 17468
rect 166540 17348 166592 17400
rect 441620 17348 441672 17400
rect 168104 17280 168156 17332
rect 445760 17280 445812 17332
rect 146208 17212 146260 17264
rect 165620 17212 165672 17264
rect 170956 17212 171008 17264
rect 492680 17212 492732 17264
rect 152556 16056 152608 16108
rect 252376 16056 252428 16108
rect 161296 15988 161348 16040
rect 361120 15988 361172 16040
rect 161020 15920 161072 15972
rect 364616 15920 364668 15972
rect 400864 15920 400916 15972
rect 478880 15920 478932 15972
rect 166816 15852 166868 15904
rect 432052 15852 432104 15904
rect 153936 14696 153988 14748
rect 272432 14696 272484 14748
rect 155960 14628 156012 14680
rect 314660 14628 314712 14680
rect 163964 14560 164016 14612
rect 398932 14560 398984 14612
rect 164148 14492 164200 14544
rect 404360 14492 404412 14544
rect 172244 14424 172296 14476
rect 503720 14424 503772 14476
rect 157984 13200 158036 13252
rect 324412 13200 324464 13252
rect 164056 13132 164108 13184
rect 407212 13132 407264 13184
rect 172336 13064 172388 13116
rect 511264 13064 511316 13116
rect 151452 11976 151504 12028
rect 245200 11976 245252 12028
rect 160008 11908 160060 11960
rect 342904 11908 342956 11960
rect 162492 11840 162544 11892
rect 390652 11840 390704 11892
rect 166724 11772 166776 11824
rect 435088 11772 435140 11824
rect 174544 11704 174596 11756
rect 548616 11704 548668 11756
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 151084 10480 151136 10532
rect 234620 10480 234672 10532
rect 159640 10412 159692 10464
rect 349252 10412 349304 10464
rect 166908 10344 166960 10396
rect 439136 10344 439188 10396
rect 105728 10276 105780 10328
rect 139584 10276 139636 10328
rect 175280 10276 175332 10328
rect 563060 10276 563112 10328
rect 142804 9596 142856 9648
rect 143540 9596 143592 9648
rect 150348 9188 150400 9240
rect 227536 9188 227588 9240
rect 161388 9120 161440 9172
rect 371700 9120 371752 9172
rect 162584 9052 162636 9104
rect 387156 9052 387208 9104
rect 168288 8984 168340 9036
rect 456892 8984 456944 9036
rect 87972 8916 88024 8968
rect 138204 8916 138256 8968
rect 176568 8916 176620 8968
rect 556160 8916 556212 8968
rect 157248 7760 157300 7812
rect 316224 7760 316276 7812
rect 162400 7692 162452 7744
rect 378876 7692 378928 7744
rect 118700 7624 118752 7676
rect 119896 7624 119948 7676
rect 169760 7624 169812 7676
rect 482836 7624 482888 7676
rect 30104 7556 30156 7608
rect 134156 7556 134208 7608
rect 175096 7556 175148 7608
rect 545488 7556 545540 7608
rect 3424 6808 3476 6860
rect 13084 6808 13136 6860
rect 576124 6808 576176 6860
rect 580172 6808 580224 6860
rect 153844 6332 153896 6384
rect 276020 6332 276072 6384
rect 165528 6264 165580 6316
rect 411904 6264 411956 6316
rect 165436 6196 165488 6248
rect 414296 6196 414348 6248
rect 103336 6128 103388 6180
rect 140320 6128 140372 6180
rect 173808 6128 173860 6180
rect 525432 6128 525484 6180
rect 152372 5040 152424 5092
rect 259552 5040 259604 5092
rect 162676 4972 162728 5024
rect 382372 4972 382424 5024
rect 180156 4904 180208 4956
rect 422576 4904 422628 4956
rect 171048 4836 171100 4888
rect 486332 4836 486384 4888
rect 144828 4768 144880 4820
rect 158904 4768 158956 4820
rect 175188 4768 175240 4820
rect 541992 4768 542044 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 118792 4088 118844 4140
rect 121460 4088 121512 4140
rect 123484 4088 123536 4140
rect 124956 4088 125008 4140
rect 1676 4020 1728 4072
rect 8944 4020 8996 4072
rect 122288 4020 122340 4072
rect 124864 4020 124916 4072
rect 131856 4088 131908 4140
rect 301596 4088 301648 4140
rect 309048 4088 309100 4140
rect 315304 4088 315356 4140
rect 317328 4088 317380 4140
rect 450544 4088 450596 4140
rect 451004 4088 451056 4140
rect 527916 4088 527968 4140
rect 529020 4088 529072 4140
rect 576216 4088 576268 4140
rect 577412 4088 577464 4140
rect 125876 4020 125928 4072
rect 129924 4020 129976 4072
rect 203616 4020 203668 4072
rect 45928 3884 45980 3936
rect 46204 3884 46256 3936
rect 106924 3748 106976 3800
rect 134524 3952 134576 4004
rect 184204 3952 184256 4004
rect 210976 3952 211028 4004
rect 85672 3680 85724 3732
rect 131028 3884 131080 3936
rect 144736 3884 144788 3936
rect 148508 3884 148560 3936
rect 151820 3884 151872 3936
rect 181444 3884 181496 3936
rect 190828 3884 190880 3936
rect 193864 3884 193916 3936
rect 196808 3884 196860 3936
rect 196900 3884 196952 3936
rect 203892 3884 203944 3936
rect 211804 3884 211856 3936
rect 247684 4020 247736 4072
rect 248788 4020 248840 4072
rect 224224 3952 224276 4004
rect 247592 3952 247644 4004
rect 124680 3816 124732 3868
rect 140872 3816 140924 3868
rect 149704 3816 149756 3868
rect 212172 3816 212224 3868
rect 231032 3884 231084 3936
rect 261484 3884 261536 3936
rect 262956 3884 263008 3936
rect 240508 3816 240560 3868
rect 242164 3816 242216 3868
rect 298468 3816 298520 3868
rect 299572 3816 299624 3868
rect 300768 3816 300820 3868
rect 311164 3816 311216 3868
rect 312636 3816 312688 3868
rect 146944 3748 146996 3800
rect 156604 3748 156656 3800
rect 156696 3748 156748 3800
rect 170772 3748 170824 3800
rect 172428 3748 172480 3800
rect 328000 3748 328052 3800
rect 357532 3748 357584 3800
rect 358728 3748 358780 3800
rect 147128 3680 147180 3732
rect 162768 3680 162820 3732
rect 377680 3680 377732 3732
rect 66720 3612 66772 3664
rect 72424 3612 72476 3664
rect 83280 3612 83332 3664
rect 138112 3612 138164 3664
rect 163688 3612 163740 3664
rect 168380 3612 168432 3664
rect 169576 3612 169628 3664
rect 178684 3612 178736 3664
rect 408408 3612 408460 3664
rect 454684 3612 454736 3664
rect 500592 3612 500644 3664
rect 19432 3544 19484 3596
rect 21364 3544 21416 3596
rect 44180 3544 44232 3596
rect 45100 3544 45152 3596
rect 51356 3544 51408 3596
rect 54484 3544 54536 3596
rect 59636 3544 59688 3596
rect 64144 3544 64196 3596
rect 69112 3544 69164 3596
rect 6460 3476 6512 3528
rect 120724 3476 120776 3528
rect 8760 3408 8812 3460
rect 10324 3408 10376 3460
rect 17040 3408 17092 3460
rect 18604 3408 18656 3460
rect 27620 3408 27672 3460
rect 28540 3408 28592 3460
rect 33600 3408 33652 3460
rect 45928 3408 45980 3460
rect 52460 3408 52512 3460
rect 53380 3408 53432 3460
rect 56048 3408 56100 3460
rect 57244 3408 57296 3460
rect 60740 3408 60792 3460
rect 61660 3408 61712 3460
rect 65524 3408 65576 3460
rect 128176 3544 128228 3596
rect 130384 3544 130436 3596
rect 135260 3544 135312 3596
rect 136456 3544 136508 3596
rect 137652 3544 137704 3596
rect 138664 3544 138716 3596
rect 141424 3544 141476 3596
rect 147128 3544 147180 3596
rect 152464 3544 152516 3596
rect 175464 3544 175516 3596
rect 180064 3544 180116 3596
rect 180340 3544 180392 3596
rect 468300 3544 468352 3596
rect 468484 3544 468536 3596
rect 469864 3544 469916 3596
rect 472624 3544 472676 3596
rect 473452 3544 473504 3596
rect 475384 3544 475436 3596
rect 518348 3544 518400 3596
rect 525064 3544 525116 3596
rect 533712 3544 533764 3596
rect 538864 3544 538916 3596
rect 539600 3544 539652 3596
rect 545764 3544 545816 3596
rect 551468 3544 551520 3596
rect 126980 3476 127032 3528
rect 128452 3476 128504 3528
rect 131212 3476 131264 3528
rect 134156 3476 134208 3528
rect 136916 3476 136968 3528
rect 148324 3476 148376 3528
rect 15936 3340 15988 3392
rect 17224 3340 17276 3392
rect 77300 3340 77352 3392
rect 78220 3340 78272 3392
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 101036 3340 101088 3392
rect 102784 3340 102836 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 130936 3408 130988 3460
rect 162492 3408 162544 3460
rect 129924 3340 129976 3392
rect 132960 3340 133012 3392
rect 141516 3340 141568 3392
rect 162124 3340 162176 3392
rect 164884 3340 164936 3392
rect 171784 3476 171836 3528
rect 173164 3476 173216 3528
rect 176660 3340 176712 3392
rect 120724 3272 120776 3324
rect 131764 3272 131816 3324
rect 147036 3272 147088 3324
rect 150624 3272 150676 3324
rect 170404 3272 170456 3324
rect 174268 3272 174320 3324
rect 181536 3476 181588 3528
rect 186136 3476 186188 3528
rect 182088 3340 182140 3392
rect 259460 3340 259512 3392
rect 260656 3340 260708 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 329104 3340 329156 3392
rect 330392 3340 330444 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 342996 3340 343048 3392
rect 344560 3340 344612 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 356704 3340 356756 3392
rect 357532 3340 357584 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 378784 3340 378836 3392
rect 379980 3340 380032 3392
rect 382924 3340 382976 3392
rect 384764 3340 384816 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 414664 3340 414716 3392
rect 416688 3340 416740 3392
rect 418804 3340 418856 3392
rect 420184 3340 420236 3392
rect 431960 3340 432012 3392
rect 433248 3340 433300 3392
rect 446404 3340 446456 3392
rect 447416 3340 447468 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 453396 3340 453448 3392
rect 454500 3340 454552 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 486424 3340 486476 3392
rect 487620 3340 487672 3392
rect 324964 3272 325016 3324
rect 326804 3272 326856 3324
rect 382280 3272 382332 3324
rect 383568 3272 383620 3324
rect 451004 3272 451056 3324
rect 452108 3272 452160 3324
rect 496084 3408 496136 3460
rect 497096 3408 497148 3460
rect 504364 3476 504416 3528
rect 507676 3476 507728 3528
rect 529204 3476 529256 3528
rect 560852 3476 560904 3528
rect 560944 3476 560996 3528
rect 572720 3544 572772 3596
rect 574744 3544 574796 3596
rect 576308 3544 576360 3596
rect 567844 3476 567896 3528
rect 569132 3476 569184 3528
rect 580264 3476 580316 3528
rect 581000 3476 581052 3528
rect 505376 3340 505428 3392
rect 583392 3408 583444 3460
rect 192484 3204 192536 3256
rect 193220 3204 193272 3256
rect 400956 3204 401008 3256
rect 402520 3204 402572 3256
rect 520924 3204 520976 3256
rect 524236 3204 524288 3256
rect 38384 3136 38436 3188
rect 39304 3136 39356 3188
rect 511356 3136 511408 3188
rect 514760 3136 514812 3188
rect 20628 3000 20680 3052
rect 22744 3000 22796 3052
rect 23020 3000 23072 3052
rect 25504 3000 25556 3052
rect 147220 3000 147272 3052
rect 148324 3000 148376 3052
rect 148416 3000 148468 3052
rect 154212 3000 154264 3052
rect 175924 3000 175976 3052
rect 177856 3000 177908 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 563704 3000 563756 3052
rect 565636 3000 565688 3052
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 12348 2932 12400 2984
rect 14464 2932 14516 2984
rect 182824 2932 182876 2984
rect 189724 2932 189776 2984
rect 423680 2864 423732 2916
rect 424968 2864 425020 2916
rect 440240 2592 440292 2644
rect 441528 2592 441580 2644
rect 390560 2456 390612 2508
rect 391848 2456 391900 2508
rect 340880 1776 340932 1828
rect 342168 1776 342220 1828
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700534 8156 703520
rect 24320 700602 24348 703520
rect 24308 700596 24360 700602
rect 24308 700538 24360 700544
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 7564 514820 7616 514826
rect 3424 514762 3476 514768
rect 7564 514762 7616 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 2778 371376 2834 371385
rect 2778 371311 2780 371320
rect 2832 371311 2834 371320
rect 2780 371282 2832 371288
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3436 265674 3464 475623
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 4804 371340 4856 371346
rect 4804 371282 4856 371288
rect 3514 358456 3570 358465
rect 3514 358391 3516 358400
rect 3568 358391 3570 358400
rect 3516 358362 3568 358368
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4816 268462 4844 371282
rect 7576 271250 7604 514762
rect 8944 358420 8996 358426
rect 8944 358362 8996 358368
rect 8956 273970 8984 358362
rect 40052 279478 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 279472 40092 279478
rect 40040 279414 40092 279420
rect 8944 273964 8996 273970
rect 8944 273906 8996 273912
rect 7564 271244 7616 271250
rect 7564 271186 7616 271192
rect 71792 269822 71820 702986
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 105464 699718 105492 703520
rect 137848 700874 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700868 137888 700874
rect 137836 700810 137888 700816
rect 152464 700392 152516 700398
rect 152464 700334 152516 700340
rect 148324 700324 148376 700330
rect 148324 700266 148376 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 71780 269816 71832 269822
rect 71780 269758 71832 269764
rect 4804 268456 4856 268462
rect 4804 268398 4856 268404
rect 3424 265668 3476 265674
rect 3424 265610 3476 265616
rect 106936 264246 106964 699654
rect 146300 696992 146352 696998
rect 146300 696934 146352 696940
rect 143632 616888 143684 616894
rect 143632 616830 143684 616836
rect 142344 590708 142396 590714
rect 142344 590650 142396 590656
rect 139400 484424 139452 484430
rect 139400 484366 139452 484372
rect 138664 430636 138716 430642
rect 138664 430578 138716 430584
rect 135260 351960 135312 351966
rect 135260 351902 135312 351908
rect 134524 324352 134576 324358
rect 134524 324294 134576 324300
rect 133144 271924 133196 271930
rect 133144 271866 133196 271872
rect 119988 269816 120040 269822
rect 119988 269758 120040 269764
rect 120000 269142 120028 269758
rect 119988 269136 120040 269142
rect 119988 269078 120040 269084
rect 106924 264240 106976 264246
rect 106924 264182 106976 264188
rect 116952 264104 117004 264110
rect 116952 264046 117004 264052
rect 114192 263696 114244 263702
rect 114192 263638 114244 263644
rect 3516 263084 3568 263090
rect 3516 263026 3568 263032
rect 3424 262880 3476 262886
rect 3424 262822 3476 262828
rect 2780 215280 2832 215286
rect 2780 215222 2832 215228
rect 2792 214985 2820 215222
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 3436 201929 3464 262822
rect 3528 254153 3556 263026
rect 114008 262676 114060 262682
rect 114008 262618 114060 262624
rect 113916 262336 113968 262342
rect 113916 262278 113968 262284
rect 14464 260976 14516 260982
rect 14464 260918 14516 260924
rect 4804 260432 4856 260438
rect 4804 260374 4856 260380
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 4816 215286 4844 260374
rect 14476 241466 14504 260918
rect 14464 241460 14516 241466
rect 14464 241402 14516 241408
rect 4804 215280 4856 215286
rect 4804 215222 4856 215228
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 104806 201104 104862 201113
rect 104806 201039 104862 201048
rect 103336 198144 103388 198150
rect 103336 198086 103388 198092
rect 102876 198008 102928 198014
rect 102876 197950 102928 197956
rect 100576 194064 100628 194070
rect 100576 194006 100628 194012
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3436 151814 3464 162823
rect 3436 151786 3556 151814
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 149122 3464 149767
rect 3424 149116 3476 149122
rect 3424 149058 3476 149064
rect 3528 145586 3556 151786
rect 100208 151224 100260 151230
rect 100208 151166 100260 151172
rect 9588 149116 9640 149122
rect 9588 149058 9640 149064
rect 9600 148374 9628 149058
rect 9588 148368 9640 148374
rect 9588 148310 9640 148316
rect 3516 145580 3568 145586
rect 3516 145522 3568 145528
rect 3424 142180 3476 142186
rect 3424 142122 3476 142128
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2872 78056 2924 78062
rect 2872 77998 2924 78004
rect 2780 77988 2832 77994
rect 2780 77930 2832 77936
rect 2792 6914 2820 77930
rect 2884 16574 2912 77998
rect 3436 45529 3464 142122
rect 8944 140956 8996 140962
rect 8944 140898 8996 140904
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 6920 78124 6972 78130
rect 6920 78066 6972 78072
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 3568 71632 3570 71641
rect 3514 71567 3570 71576
rect 4160 64184 4212 64190
rect 4160 64126 4212 64132
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 64126
rect 6932 16574 6960 78066
rect 7562 75168 7618 75177
rect 7562 75103 7618 75112
rect 2884 16546 3648 16574
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 2792 6886 2912 6914
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1688 480 1716 4014
rect 2884 480 2912 6886
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 7484 3482 7512 16546
rect 7576 4146 7604 75103
rect 8956 71670 8984 140898
rect 31024 139528 31076 139534
rect 31024 139470 31076 139476
rect 13084 139460 13136 139466
rect 13084 139402 13136 139408
rect 8944 71664 8996 71670
rect 8944 71606 8996 71612
rect 8942 68232 8998 68241
rect 8942 68167 8998 68176
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 8956 4078 8984 68167
rect 11058 66872 11114 66881
rect 11058 66807 11114 66816
rect 10324 62824 10376 62830
rect 10324 62766 10376 62772
rect 9680 53100 9732 53106
rect 9680 53042 9732 53048
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 6472 480 6500 3470
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8772 480 8800 3402
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 53042
rect 10336 3466 10364 62766
rect 11072 16574 11100 66807
rect 12440 55888 12492 55894
rect 12440 55830 12492 55836
rect 12452 16574 12480 55830
rect 11072 16546 11192 16574
rect 12452 16546 13032 16574
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11164 480 11192 16546
rect 13004 3482 13032 16546
rect 13096 6866 13124 139402
rect 31036 111790 31064 139470
rect 31024 111784 31076 111790
rect 31024 111726 31076 111732
rect 77298 81560 77354 81569
rect 77298 81495 77354 81504
rect 71780 80708 71832 80714
rect 71780 80650 71832 80656
rect 46940 78396 46992 78402
rect 46940 78338 46992 78344
rect 20720 78192 20772 78198
rect 20720 78134 20772 78140
rect 14462 73808 14518 73817
rect 14462 73743 14518 73752
rect 13820 40724 13872 40730
rect 13820 40666 13872 40672
rect 13832 16574 13860 40666
rect 13832 16546 14320 16574
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13004 3454 13584 3482
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 480 12388 2926
rect 13556 480 13584 3454
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 2990 14504 73743
rect 18604 69692 18656 69698
rect 18604 69634 18656 69640
rect 17960 60036 18012 60042
rect 17960 59978 18012 59984
rect 17222 36544 17278 36553
rect 17222 36479 17278 36488
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 15948 480 15976 3334
rect 17052 480 17080 3402
rect 17236 3398 17264 36479
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 59978
rect 18616 3466 18644 69634
rect 20732 16574 20760 78134
rect 34520 76696 34572 76702
rect 34520 76638 34572 76644
rect 22742 75304 22798 75313
rect 22742 75239 22798 75248
rect 21364 72548 21416 72554
rect 21364 72490 21416 72496
rect 20732 16546 21312 16574
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 19444 480 19472 3538
rect 21284 3482 21312 16546
rect 21376 3602 21404 72490
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21284 3454 21864 3482
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20640 480 20668 2994
rect 21836 480 21864 3454
rect 22756 3058 22784 75239
rect 26238 73944 26294 73953
rect 26238 73879 26294 73888
rect 23480 60104 23532 60110
rect 23480 60046 23532 60052
rect 23492 16574 23520 60046
rect 25502 57216 25558 57225
rect 25502 57151 25558 57160
rect 24858 33824 24914 33833
rect 24858 33759 24914 33768
rect 24872 16574 24900 33759
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23032 480 23060 2994
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 25516 3058 25544 57151
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 73879
rect 27620 71052 27672 71058
rect 27620 70994 27672 71000
rect 27632 3466 27660 70994
rect 27710 51776 27766 51785
rect 27710 51711 27766 51720
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27724 480 27752 51711
rect 30380 50380 30432 50386
rect 30380 50322 30432 50328
rect 30392 16574 30420 50322
rect 31760 39364 31812 39370
rect 31760 39306 31812 39312
rect 31772 16574 31800 39306
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 30104 7608 30156 7614
rect 30104 7550 30156 7556
rect 28540 3460 28592 3466
rect 28540 3402 28592 3408
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3402
rect 30116 480 30144 7550
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33612 480 33640 3402
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 76638
rect 35900 76560 35952 76566
rect 35900 76502 35952 76508
rect 35912 6914 35940 76502
rect 45560 72480 45612 72486
rect 45560 72422 45612 72428
rect 41420 69760 41472 69766
rect 41420 69702 41472 69708
rect 40038 67008 40094 67017
rect 40038 66943 40094 66952
rect 35992 65544 36044 65550
rect 35992 65486 36044 65492
rect 36004 16574 36032 65486
rect 39302 48920 39358 48929
rect 39302 48855 39358 48864
rect 38660 37936 38712 37942
rect 38660 37878 38712 37884
rect 38672 16574 38700 37878
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 480 38424 3130
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3194 39344 48855
rect 40052 16574 40080 66943
rect 41432 16574 41460 69702
rect 42800 61396 42852 61402
rect 42800 61338 42852 61344
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 61338
rect 44178 47560 44234 47569
rect 44178 47495 44234 47504
rect 44192 3602 44220 47495
rect 44272 31068 44324 31074
rect 44272 31010 44324 31016
rect 44180 3596 44232 3602
rect 44180 3538 44232 3544
rect 44284 480 44312 31010
rect 45572 16574 45600 72422
rect 46204 69828 46256 69834
rect 46204 69770 46256 69776
rect 45572 16546 46152 16574
rect 45928 3936 45980 3942
rect 45928 3878 45980 3884
rect 45100 3596 45152 3602
rect 45100 3538 45152 3544
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3538
rect 45940 3466 45968 3878
rect 46124 3482 46152 16546
rect 46216 3942 46244 69770
rect 46952 16574 46980 78338
rect 57980 78328 58032 78334
rect 57980 78270 58032 78276
rect 52460 76628 52512 76634
rect 52460 76570 52512 76576
rect 48320 68332 48372 68338
rect 48320 68274 48372 68280
rect 48332 16574 48360 68274
rect 49698 58576 49754 58585
rect 49698 58511 49754 58520
rect 49712 16574 49740 58511
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 3936 46256 3942
rect 46204 3878 46256 3884
rect 45928 3460 45980 3466
rect 46124 3454 46704 3482
rect 45928 3402 45980 3408
rect 46676 480 46704 3454
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 51368 480 51396 3538
rect 52472 3466 52500 76570
rect 54484 73840 54536 73846
rect 54484 73782 54536 73788
rect 52552 61464 52604 61470
rect 52552 61406 52604 61412
rect 52460 3460 52512 3466
rect 52460 3402 52512 3408
rect 52564 480 52592 61406
rect 53840 35216 53892 35222
rect 53840 35158 53892 35164
rect 53852 16574 53880 35158
rect 53852 16546 54432 16574
rect 54404 3482 54432 16546
rect 54496 3602 54524 73782
rect 57244 65612 57296 65618
rect 57244 65554 57296 65560
rect 56598 46200 56654 46209
rect 56598 46135 56654 46144
rect 56612 16574 56640 46135
rect 56612 16546 56824 16574
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 53380 3460 53432 3466
rect 54404 3454 54984 3482
rect 53380 3402 53432 3408
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3402
rect 54956 480 54984 3454
rect 56048 3460 56100 3466
rect 56048 3402 56100 3408
rect 56060 480 56088 3402
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3466 57284 65554
rect 57992 16574 58020 78270
rect 64144 76764 64196 76770
rect 64144 76706 64196 76712
rect 60740 66904 60792 66910
rect 60740 66846 60792 66852
rect 57992 16546 58480 16574
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 58452 480 58480 16546
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59648 480 59676 3538
rect 60752 3466 60780 66846
rect 62120 64252 62172 64258
rect 62120 64194 62172 64200
rect 60832 44872 60884 44878
rect 60832 44814 60884 44820
rect 60740 3460 60792 3466
rect 60740 3402 60792 3408
rect 60844 480 60872 44814
rect 62132 16574 62160 64194
rect 63500 55956 63552 55962
rect 63500 55898 63552 55904
rect 63512 16574 63540 55898
rect 62132 16546 63264 16574
rect 63512 16546 64092 16574
rect 61660 3460 61712 3466
rect 61660 3402 61712 3408
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61672 354 61700 3402
rect 63236 480 63264 16546
rect 64064 3482 64092 16546
rect 64156 3602 64184 76706
rect 67640 75200 67692 75206
rect 67640 75142 67692 75148
rect 66720 3664 66772 3670
rect 66720 3606 66772 3612
rect 64144 3596 64196 3602
rect 64144 3538 64196 3544
rect 64064 3454 64368 3482
rect 64340 480 64368 3454
rect 65524 3460 65576 3466
rect 65524 3402 65576 3408
rect 65536 480 65564 3402
rect 66732 480 66760 3606
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 75142
rect 70400 72616 70452 72622
rect 70400 72558 70452 72564
rect 69020 60172 69072 60178
rect 69020 60114 69072 60120
rect 69032 16574 69060 60114
rect 70412 16574 70440 72558
rect 71792 16574 71820 80650
rect 72424 76832 72476 76838
rect 72424 76774 72476 76780
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72372 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 69124 480 69152 3538
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72344 3482 72372 16546
rect 72436 3670 72464 76774
rect 75920 67040 75972 67046
rect 75920 66982 75972 66988
rect 75184 62960 75236 62966
rect 75184 62902 75236 62908
rect 74540 43444 74592 43450
rect 74540 43386 74592 43392
rect 74552 16574 74580 43386
rect 74552 16546 75040 16574
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 72424 3664 72476 3670
rect 72424 3606 72476 3612
rect 72344 3454 72648 3482
rect 72620 480 72648 3454
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 62902
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 66982
rect 77312 3398 77340 81495
rect 85580 80776 85632 80782
rect 85580 80718 85632 80724
rect 81440 75268 81492 75274
rect 81440 75210 81492 75216
rect 78680 67108 78732 67114
rect 78680 67050 78732 67056
rect 77392 57248 77444 57254
rect 77392 57190 77444 57196
rect 77300 3392 77352 3398
rect 77300 3334 77352 3340
rect 77404 480 77432 57190
rect 78692 16574 78720 67050
rect 80060 66972 80112 66978
rect 80060 66914 80112 66920
rect 80072 16574 80100 66914
rect 81452 16574 81480 75210
rect 84200 54596 84252 54602
rect 84200 54538 84252 54544
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 78220 3392 78272 3398
rect 78220 3334 78272 3340
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3334
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 3664 83332 3670
rect 83280 3606 83332 3612
rect 83292 480 83320 3606
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 54538
rect 85592 16574 85620 80718
rect 100116 79348 100168 79354
rect 100116 79290 100168 79296
rect 96620 75744 96672 75750
rect 96620 75686 96672 75692
rect 95240 73908 95292 73914
rect 95240 73850 95292 73856
rect 89720 69896 89772 69902
rect 89720 69838 89772 69844
rect 88340 62892 88392 62898
rect 88340 62834 88392 62840
rect 88352 16574 88380 62834
rect 89732 16574 89760 69838
rect 93858 67144 93914 67153
rect 93858 67079 93914 67088
rect 93124 65680 93176 65686
rect 93124 65622 93176 65628
rect 92478 64152 92534 64161
rect 92478 64087 92534 64096
rect 85592 16546 86448 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 85672 3732 85724 3738
rect 85672 3674 85724 3680
rect 85684 480 85712 3674
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87972 8968 88024 8974
rect 87972 8910 88024 8916
rect 87984 480 88012 8910
rect 89180 480 89208 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 86838 -960 86950 326
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 91572 480 91600 3334
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 64087
rect 93136 3398 93164 65622
rect 93872 3398 93900 67079
rect 93952 50448 94004 50454
rect 93952 50390 94004 50396
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 50390
rect 95252 16574 95280 73850
rect 96632 16574 96660 75686
rect 100128 71602 100156 79290
rect 100220 72962 100248 151166
rect 100300 151156 100352 151162
rect 100300 151098 100352 151104
rect 100312 79354 100340 151098
rect 100392 151088 100444 151094
rect 100392 151030 100444 151036
rect 100300 79348 100352 79354
rect 100300 79290 100352 79296
rect 100208 72956 100260 72962
rect 100208 72898 100260 72904
rect 100220 72554 100248 72898
rect 100208 72548 100260 72554
rect 100208 72490 100260 72496
rect 100116 71596 100168 71602
rect 100116 71538 100168 71544
rect 100128 71058 100156 71538
rect 100116 71052 100168 71058
rect 100116 70994 100168 71000
rect 98000 65748 98052 65754
rect 98000 65690 98052 65696
rect 98012 16574 98040 65690
rect 100404 60722 100432 151030
rect 100482 148336 100538 148345
rect 100482 148271 100538 148280
rect 99380 60716 99432 60722
rect 99380 60658 99432 60664
rect 100392 60716 100444 60722
rect 100392 60658 100444 60664
rect 99392 60110 99420 60658
rect 99472 60648 99524 60654
rect 99472 60590 99524 60596
rect 99380 60104 99432 60110
rect 99380 60046 99432 60052
rect 99484 60042 99512 60590
rect 99472 60036 99524 60042
rect 99472 59978 99524 59984
rect 99380 56568 99432 56574
rect 99380 56510 99432 56516
rect 99392 55894 99420 56510
rect 99380 55888 99432 55894
rect 99380 55830 99432 55836
rect 99380 54528 99432 54534
rect 99380 54470 99432 54476
rect 99392 16574 99420 54470
rect 100496 53786 100524 148271
rect 100588 60654 100616 194006
rect 101680 193996 101732 194002
rect 101680 193938 101732 193944
rect 100666 193896 100722 193905
rect 100666 193831 100722 193840
rect 100576 60648 100628 60654
rect 100576 60590 100628 60596
rect 100680 56574 100708 193831
rect 101588 189916 101640 189922
rect 101588 189858 101640 189864
rect 101600 77042 101628 189858
rect 100760 77036 100812 77042
rect 100760 76978 100812 76984
rect 101588 77036 101640 77042
rect 101588 76978 101640 76984
rect 100772 76702 100800 76978
rect 100760 76696 100812 76702
rect 100760 76638 100812 76644
rect 101692 57905 101720 193938
rect 102784 192568 102836 192574
rect 102784 192510 102836 192516
rect 101772 190120 101824 190126
rect 101772 190062 101824 190068
rect 100758 57896 100814 57905
rect 100758 57831 100814 57840
rect 101678 57896 101734 57905
rect 101678 57831 101734 57840
rect 100772 57225 100800 57831
rect 100758 57216 100814 57225
rect 100758 57151 100814 57160
rect 100668 56568 100720 56574
rect 100668 56510 100720 56516
rect 100484 53780 100536 53786
rect 100484 53722 100536 53728
rect 100496 53106 100524 53722
rect 100484 53100 100536 53106
rect 100484 53042 100536 53048
rect 101784 52465 101812 190062
rect 101864 190052 101916 190058
rect 101864 189994 101916 190000
rect 100758 52456 100814 52465
rect 100758 52391 100814 52400
rect 101770 52456 101826 52465
rect 101770 52391 101826 52400
rect 100772 51785 100800 52391
rect 100758 51776 100814 51785
rect 100758 51711 100814 51720
rect 101876 51066 101904 189994
rect 102048 189848 102100 189854
rect 102048 189790 102100 189796
rect 101956 189780 102008 189786
rect 101956 189722 102008 189728
rect 100760 51060 100812 51066
rect 100760 51002 100812 51008
rect 101864 51060 101916 51066
rect 101864 51002 101916 51008
rect 100772 50386 100800 51002
rect 100760 50380 100812 50386
rect 100760 50322 100812 50328
rect 101968 49609 101996 189722
rect 100758 49600 100814 49609
rect 100758 49535 100814 49544
rect 101954 49600 102010 49609
rect 101954 49535 102010 49544
rect 100772 48929 100800 49535
rect 100758 48920 100814 48929
rect 100758 48855 100814 48864
rect 102060 48249 102088 189790
rect 102692 148776 102744 148782
rect 102692 148718 102744 148724
rect 102140 78668 102192 78674
rect 102140 78610 102192 78616
rect 102152 78198 102180 78610
rect 102140 78192 102192 78198
rect 102140 78134 102192 78140
rect 102140 70032 102192 70038
rect 102140 69974 102192 69980
rect 102152 69766 102180 69974
rect 102140 69760 102192 69766
rect 102140 69702 102192 69708
rect 102138 67416 102194 67425
rect 102138 67351 102194 67360
rect 102152 67017 102180 67351
rect 102138 67008 102194 67017
rect 102138 66943 102194 66952
rect 102140 66224 102192 66230
rect 102140 66166 102192 66172
rect 102152 65618 102180 66166
rect 102140 65612 102192 65618
rect 102140 65554 102192 65560
rect 102138 53136 102194 53145
rect 102138 53071 102194 53080
rect 100758 48240 100814 48249
rect 100758 48175 100814 48184
rect 102046 48240 102102 48249
rect 102046 48175 102102 48184
rect 100772 47569 100800 48175
rect 100758 47560 100814 47569
rect 100758 47495 100814 47504
rect 102152 16574 102180 53071
rect 102704 46889 102732 148718
rect 102796 77178 102824 192510
rect 102888 78674 102916 197950
rect 103060 195764 103112 195770
rect 103060 195706 103112 195712
rect 102968 189984 103020 189990
rect 102968 189926 103020 189932
rect 102876 78668 102928 78674
rect 102876 78610 102928 78616
rect 102784 77172 102836 77178
rect 102784 77114 102836 77120
rect 102784 71052 102836 71058
rect 102784 70994 102836 71000
rect 102230 46880 102286 46889
rect 102230 46815 102286 46824
rect 102690 46880 102746 46889
rect 102690 46815 102746 46824
rect 102244 46209 102272 46815
rect 102230 46200 102286 46209
rect 102230 46135 102286 46144
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 102152 16546 102272 16574
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 101048 480 101076 3334
rect 102244 480 102272 16546
rect 102796 3398 102824 70994
rect 102980 70038 103008 189926
rect 103072 73953 103100 195706
rect 103152 193928 103204 193934
rect 103152 193870 103204 193876
rect 103058 73944 103114 73953
rect 103058 73879 103114 73888
rect 102968 70032 103020 70038
rect 102968 69974 103020 69980
rect 103164 67425 103192 193870
rect 103242 192536 103298 192545
rect 103242 192471 103298 192480
rect 103150 67416 103206 67425
rect 103150 67351 103206 67360
rect 103256 66230 103284 192471
rect 103348 69834 103376 198086
rect 103428 198076 103480 198082
rect 103428 198018 103480 198024
rect 103336 69828 103388 69834
rect 103336 69770 103388 69776
rect 103440 69698 103468 198018
rect 104438 196888 104494 196897
rect 104438 196823 104494 196832
rect 104164 194472 104216 194478
rect 104164 194414 104216 194420
rect 104072 148640 104124 148646
rect 104072 148582 104124 148588
rect 103520 69964 103572 69970
rect 103520 69906 103572 69912
rect 103428 69692 103480 69698
rect 103428 69634 103480 69640
rect 103244 66224 103296 66230
rect 103244 66166 103296 66172
rect 103532 16574 103560 69906
rect 104084 58585 104112 148582
rect 104176 80322 104204 194414
rect 104348 194200 104400 194206
rect 104348 194142 104400 194148
rect 104256 192704 104308 192710
rect 104256 192646 104308 192652
rect 104268 80442 104296 192646
rect 104256 80436 104308 80442
rect 104256 80378 104308 80384
rect 104176 80294 104296 80322
rect 104164 80232 104216 80238
rect 104164 80174 104216 80180
rect 104176 77217 104204 80174
rect 104268 78606 104296 80294
rect 104256 78600 104308 78606
rect 104256 78542 104308 78548
rect 104268 78062 104296 78542
rect 104256 78056 104308 78062
rect 104256 77998 104308 78004
rect 104162 77208 104218 77217
rect 104162 77143 104218 77152
rect 104176 62966 104204 77143
rect 104360 72826 104388 194142
rect 104348 72820 104400 72826
rect 104348 72762 104400 72768
rect 104452 71398 104480 196823
rect 104716 194268 104768 194274
rect 104716 194210 104768 194216
rect 104622 194168 104678 194177
rect 104532 194132 104584 194138
rect 104622 194103 104678 194112
rect 104532 194074 104584 194080
rect 104440 71392 104492 71398
rect 104440 71334 104492 71340
rect 104544 68950 104572 194074
rect 104532 68944 104584 68950
rect 104532 68886 104584 68892
rect 104636 63510 104664 194103
rect 104624 63504 104676 63510
rect 104624 63446 104676 63452
rect 104164 62960 104216 62966
rect 104164 62902 104216 62908
rect 104636 62830 104664 63446
rect 104624 62824 104676 62830
rect 104624 62766 104676 62772
rect 104728 62082 104756 194210
rect 104820 69034 104848 201039
rect 111708 200660 111760 200666
rect 111708 200602 111760 200608
rect 107290 200424 107346 200433
rect 107200 200388 107252 200394
rect 107290 200359 107346 200368
rect 107200 200330 107252 200336
rect 106924 198280 106976 198286
rect 106924 198222 106976 198228
rect 106832 196784 106884 196790
rect 106832 196726 106884 196732
rect 106096 196648 106148 196654
rect 106096 196590 106148 196596
rect 105636 195424 105688 195430
rect 105636 195366 105688 195372
rect 105648 80782 105676 195366
rect 105820 195356 105872 195362
rect 105820 195298 105872 195304
rect 105728 193180 105780 193186
rect 105728 193122 105780 193128
rect 105636 80776 105688 80782
rect 105636 80718 105688 80724
rect 105740 76906 105768 193122
rect 105728 76900 105780 76906
rect 105728 76842 105780 76848
rect 105832 75750 105860 195298
rect 105912 193860 105964 193866
rect 105912 193802 105964 193808
rect 105820 75744 105872 75750
rect 105820 75686 105872 75692
rect 105924 73166 105952 193802
rect 106004 192840 106056 192846
rect 106004 192782 106056 192788
rect 105912 73160 105964 73166
rect 105912 73102 105964 73108
rect 105542 71904 105598 71913
rect 105542 71839 105598 71848
rect 104820 69006 104940 69034
rect 104808 68944 104860 68950
rect 104808 68886 104860 68892
rect 104820 68338 104848 68886
rect 104808 68332 104860 68338
rect 104808 68274 104860 68280
rect 104912 68218 104940 69006
rect 104820 68190 104940 68218
rect 104820 66094 104848 68190
rect 104808 66088 104860 66094
rect 104808 66030 104860 66036
rect 104820 65550 104848 66030
rect 104808 65544 104860 65550
rect 104808 65486 104860 65492
rect 104532 62076 104584 62082
rect 104532 62018 104584 62024
rect 104716 62076 104768 62082
rect 104716 62018 104768 62024
rect 104544 61470 104572 62018
rect 104532 61464 104584 61470
rect 104532 61406 104584 61412
rect 104806 59256 104862 59265
rect 104806 59191 104862 59200
rect 104820 58585 104848 59191
rect 104070 58576 104126 58585
rect 104070 58511 104126 58520
rect 104806 58576 104862 58585
rect 104806 58511 104862 58520
rect 105556 50454 105584 71839
rect 106016 70174 106044 192782
rect 106108 72729 106136 196590
rect 106186 192672 106242 192681
rect 106186 192607 106242 192616
rect 106094 72720 106150 72729
rect 106094 72655 106150 72664
rect 106108 71913 106136 72655
rect 106094 71904 106150 71913
rect 106094 71839 106150 71848
rect 106004 70168 106056 70174
rect 106004 70110 106056 70116
rect 106016 69970 106044 70110
rect 106004 69964 106056 69970
rect 106004 69906 106056 69912
rect 106200 64870 106228 192607
rect 106844 79626 106872 196726
rect 106832 79620 106884 79626
rect 106832 79562 106884 79568
rect 106844 71058 106872 79562
rect 106936 78266 106964 198222
rect 107106 196616 107162 196625
rect 107106 196551 107162 196560
rect 107016 195696 107068 195702
rect 107016 195638 107068 195644
rect 106924 78260 106976 78266
rect 106924 78202 106976 78208
rect 107028 75614 107056 195638
rect 107120 75721 107148 196551
rect 107212 78282 107240 200330
rect 107304 78470 107332 200359
rect 107382 200152 107438 200161
rect 107382 200087 107438 200096
rect 107292 78464 107344 78470
rect 107292 78406 107344 78412
rect 107292 78328 107344 78334
rect 107212 78276 107292 78282
rect 107212 78270 107344 78276
rect 107212 78254 107332 78270
rect 107304 77790 107332 78254
rect 107292 77784 107344 77790
rect 107292 77726 107344 77732
rect 107106 75712 107162 75721
rect 107106 75647 107162 75656
rect 107016 75608 107068 75614
rect 107016 75550 107068 75556
rect 106832 71052 106884 71058
rect 106832 70994 106884 71000
rect 107028 69902 107056 75550
rect 107016 69896 107068 69902
rect 107016 69838 107068 69844
rect 107120 67046 107148 75647
rect 107396 73846 107424 200087
rect 111248 199708 111300 199714
rect 111248 199650 111300 199656
rect 108856 199232 108908 199238
rect 108856 199174 108908 199180
rect 108946 199200 109002 199209
rect 108672 198552 108724 198558
rect 108672 198494 108724 198500
rect 108396 198416 108448 198422
rect 108396 198358 108448 198364
rect 108210 197024 108266 197033
rect 108210 196959 108266 196968
rect 107476 192432 107528 192438
rect 107476 192374 107528 192380
rect 107384 73840 107436 73846
rect 107384 73782 107436 73788
rect 107396 73642 107424 73782
rect 107384 73636 107436 73642
rect 107384 73578 107436 73584
rect 107108 67040 107160 67046
rect 107108 66982 107160 66988
rect 106188 64864 106240 64870
rect 106188 64806 106240 64812
rect 106200 64258 106228 64806
rect 106188 64252 106240 64258
rect 106188 64194 106240 64200
rect 107488 60586 107516 192374
rect 107568 190188 107620 190194
rect 107568 190130 107620 190136
rect 107476 60580 107528 60586
rect 107476 60522 107528 60528
rect 107488 60178 107516 60522
rect 107476 60172 107528 60178
rect 107476 60114 107528 60120
rect 107580 53825 107608 190130
rect 108224 80850 108252 196959
rect 108304 193112 108356 193118
rect 108304 193054 108356 193060
rect 108212 80844 108264 80850
rect 108212 80786 108264 80792
rect 108224 80714 108252 80786
rect 108212 80708 108264 80714
rect 108212 80650 108264 80656
rect 108316 74322 108344 193054
rect 108408 77994 108436 198358
rect 108486 196752 108542 196761
rect 108486 196687 108542 196696
rect 108396 77988 108448 77994
rect 108396 77930 108448 77936
rect 108500 75449 108528 196687
rect 108580 192500 108632 192506
rect 108580 192442 108632 192448
rect 108486 75440 108542 75449
rect 108486 75375 108542 75384
rect 108304 74316 108356 74322
rect 108304 74258 108356 74264
rect 108316 73234 108344 74258
rect 107660 73228 107712 73234
rect 107660 73170 107712 73176
rect 108304 73228 108356 73234
rect 108304 73170 108356 73176
rect 107566 53816 107622 53825
rect 107566 53751 107622 53760
rect 107580 53145 107608 53751
rect 107566 53136 107622 53145
rect 107566 53071 107622 53080
rect 105544 50448 105596 50454
rect 105544 50390 105596 50396
rect 107672 16574 107700 73170
rect 108500 67114 108528 75375
rect 108592 71330 108620 192442
rect 108684 73817 108712 198494
rect 108764 194336 108816 194342
rect 108764 194278 108816 194284
rect 108670 73808 108726 73817
rect 108670 73743 108726 73752
rect 108580 71324 108632 71330
rect 108580 71266 108632 71272
rect 108776 67153 108804 194278
rect 108868 71262 108896 199174
rect 108946 199135 109002 199144
rect 108856 71256 108908 71262
rect 108856 71198 108908 71204
rect 108960 67522 108988 199135
rect 110328 196920 110380 196926
rect 110328 196862 110380 196868
rect 109776 196716 109828 196722
rect 109776 196658 109828 196664
rect 109788 76673 109816 196658
rect 110236 195628 110288 195634
rect 110236 195570 110288 195576
rect 110144 193044 110196 193050
rect 110144 192986 110196 192992
rect 110052 192908 110104 192914
rect 110052 192850 110104 192856
rect 109868 192636 109920 192642
rect 109868 192578 109920 192584
rect 109774 76664 109830 76673
rect 109774 76599 109830 76608
rect 109880 71777 109908 192578
rect 109960 190324 110012 190330
rect 109960 190266 110012 190272
rect 109866 71768 109922 71777
rect 109866 71703 109922 71712
rect 109040 69012 109092 69018
rect 109040 68954 109092 68960
rect 108948 67516 109000 67522
rect 108948 67458 109000 67464
rect 108762 67144 108818 67153
rect 108488 67108 108540 67114
rect 108762 67079 108818 67088
rect 108488 67050 108540 67056
rect 103532 16546 104112 16574
rect 107672 16546 108160 16574
rect 103336 6180 103388 6186
rect 103336 6122 103388 6128
rect 102784 3392 102836 3398
rect 102784 3334 102836 3340
rect 103348 480 103376 6122
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 10328 105780 10334
rect 105728 10270 105780 10276
rect 105740 480 105768 10270
rect 106924 3800 106976 3806
rect 106924 3742 106976 3748
rect 106936 480 106964 3742
rect 108132 480 108160 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 68954
rect 109972 66162 110000 190266
rect 110064 67590 110092 192850
rect 110052 67584 110104 67590
rect 110156 67561 110184 192986
rect 110248 69970 110276 195570
rect 110236 69964 110288 69970
rect 110236 69906 110288 69912
rect 110340 69902 110368 196862
rect 111064 194404 111116 194410
rect 111064 194346 111116 194352
rect 110972 190392 111024 190398
rect 110972 190334 111024 190340
rect 110880 146940 110932 146946
rect 110880 146882 110932 146888
rect 110328 69896 110380 69902
rect 110328 69838 110380 69844
rect 110052 67526 110104 67532
rect 110142 67552 110198 67561
rect 110142 67487 110198 67496
rect 110418 67008 110474 67017
rect 110418 66943 110474 66952
rect 109132 66156 109184 66162
rect 109132 66098 109184 66104
rect 109960 66156 110012 66162
rect 109960 66098 110012 66104
rect 109144 65754 109172 66098
rect 109132 65748 109184 65754
rect 109132 65690 109184 65696
rect 110432 3398 110460 66943
rect 110892 64841 110920 146882
rect 110984 80102 111012 190334
rect 110972 80096 111024 80102
rect 110972 80038 111024 80044
rect 110984 69018 111012 80038
rect 111076 79490 111104 194346
rect 111156 192976 111208 192982
rect 111156 192918 111208 192924
rect 111064 79484 111116 79490
rect 111064 79426 111116 79432
rect 111168 74526 111196 192918
rect 111260 79422 111288 199650
rect 111524 199640 111576 199646
rect 111524 199582 111576 199588
rect 111340 196852 111392 196858
rect 111340 196794 111392 196800
rect 111248 79416 111300 79422
rect 111248 79358 111300 79364
rect 111352 76770 111380 196794
rect 111432 195900 111484 195906
rect 111432 195842 111484 195848
rect 111340 76764 111392 76770
rect 111340 76706 111392 76712
rect 111156 74520 111208 74526
rect 111156 74462 111208 74468
rect 111444 72758 111472 195842
rect 111536 75886 111564 199582
rect 111616 197124 111668 197130
rect 111616 197066 111668 197072
rect 111524 75880 111576 75886
rect 111524 75822 111576 75828
rect 111432 72752 111484 72758
rect 111432 72694 111484 72700
rect 111628 72690 111656 197066
rect 111720 74458 111748 200602
rect 112996 200456 113048 200462
rect 112996 200398 113048 200404
rect 112812 199504 112864 199510
rect 112812 199446 112864 199452
rect 112720 196988 112772 196994
rect 112720 196930 112772 196936
rect 112442 195392 112498 195401
rect 112442 195327 112498 195336
rect 112352 190256 112404 190262
rect 112352 190198 112404 190204
rect 112260 147076 112312 147082
rect 112260 147018 112312 147024
rect 111798 76936 111854 76945
rect 111798 76871 111854 76880
rect 111708 74452 111760 74458
rect 111708 74394 111760 74400
rect 111616 72684 111668 72690
rect 111616 72626 111668 72632
rect 110972 69012 111024 69018
rect 110972 68954 111024 68960
rect 110878 64832 110934 64841
rect 110878 64767 110934 64776
rect 110892 64161 110920 64767
rect 110878 64152 110934 64161
rect 110878 64087 110934 64096
rect 110512 59356 110564 59362
rect 110512 59298 110564 59304
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 59298
rect 111812 16574 111840 76871
rect 112272 74534 112300 147018
rect 112364 76945 112392 190198
rect 112456 79354 112484 195327
rect 112628 195288 112680 195294
rect 112628 195230 112680 195236
rect 112536 193792 112588 193798
rect 112536 193734 112588 193740
rect 112444 79348 112496 79354
rect 112444 79290 112496 79296
rect 112350 76936 112406 76945
rect 112350 76871 112406 76880
rect 112548 76498 112576 193734
rect 112640 77246 112668 195230
rect 112628 77240 112680 77246
rect 112628 77182 112680 77188
rect 112536 76492 112588 76498
rect 112536 76434 112588 76440
rect 112272 74506 112484 74534
rect 112456 71233 112484 74506
rect 112442 71224 112498 71233
rect 112442 71159 112498 71168
rect 112456 43450 112484 71159
rect 112548 57254 112576 76434
rect 112732 74186 112760 196930
rect 112824 75857 112852 199446
rect 112904 197260 112956 197266
rect 112904 197202 112956 197208
rect 112810 75848 112866 75857
rect 112810 75783 112866 75792
rect 112720 74180 112772 74186
rect 112720 74122 112772 74128
rect 112916 72554 112944 197202
rect 113008 74050 113036 200398
rect 113088 200320 113140 200326
rect 113088 200262 113140 200268
rect 113100 74497 113128 200262
rect 113824 190460 113876 190466
rect 113824 190402 113876 190408
rect 113364 148980 113416 148986
rect 113364 148922 113416 148928
rect 113086 74488 113142 74497
rect 113086 74423 113142 74432
rect 112996 74044 113048 74050
rect 112996 73986 113048 73992
rect 112904 72548 112956 72554
rect 112904 72490 112956 72496
rect 113376 71194 113404 148922
rect 113548 148300 113600 148306
rect 113548 148242 113600 148248
rect 113454 146976 113510 146985
rect 113454 146911 113510 146920
rect 113468 73982 113496 146911
rect 113456 73976 113508 73982
rect 113456 73918 113508 73924
rect 113364 71188 113416 71194
rect 113364 71130 113416 71136
rect 113180 67040 113232 67046
rect 113180 66982 113232 66988
rect 112536 57248 112588 57254
rect 112536 57190 112588 57196
rect 112444 43444 112496 43450
rect 112444 43386 112496 43392
rect 113192 16574 113220 66982
rect 113468 66978 113496 73918
rect 113560 69698 113588 148242
rect 113732 143540 113784 143546
rect 113732 143482 113784 143488
rect 113640 141772 113692 141778
rect 113640 141714 113692 141720
rect 113652 78062 113680 141714
rect 113640 78056 113692 78062
rect 113640 77998 113692 78004
rect 113744 77994 113772 143482
rect 113836 79558 113864 190402
rect 113928 147286 113956 262278
rect 113916 147280 113968 147286
rect 113916 147222 113968 147228
rect 114020 143206 114048 262618
rect 114100 195832 114152 195838
rect 114100 195774 114152 195780
rect 114008 143200 114060 143206
rect 114008 143142 114060 143148
rect 113824 79552 113876 79558
rect 113824 79494 113876 79500
rect 113732 77988 113784 77994
rect 113732 77930 113784 77936
rect 114112 74254 114140 195774
rect 114204 141642 114232 263638
rect 116860 262812 116912 262818
rect 116860 262754 116912 262760
rect 116768 262744 116820 262750
rect 116768 262686 116820 262692
rect 115296 261044 115348 261050
rect 115296 260986 115348 260992
rect 114376 199164 114428 199170
rect 114376 199106 114428 199112
rect 114284 195560 114336 195566
rect 114284 195502 114336 195508
rect 114192 141636 114244 141642
rect 114192 141578 114244 141584
rect 114100 74248 114152 74254
rect 114100 74190 114152 74196
rect 114296 73098 114324 195502
rect 114388 75585 114416 199106
rect 114468 198960 114520 198966
rect 114468 198902 114520 198908
rect 114374 75576 114430 75585
rect 114374 75511 114430 75520
rect 114480 75070 114508 198902
rect 115202 192808 115258 192817
rect 115202 192743 115258 192752
rect 115020 147212 115072 147218
rect 115020 147154 115072 147160
rect 114928 147144 114980 147150
rect 114928 147086 114980 147092
rect 114560 77104 114612 77110
rect 114560 77046 114612 77052
rect 114468 75064 114520 75070
rect 114468 75006 114520 75012
rect 114284 73092 114336 73098
rect 114284 73034 114336 73040
rect 113548 69692 113600 69698
rect 113548 69634 113600 69640
rect 113456 66972 113508 66978
rect 113456 66914 113508 66920
rect 114572 16574 114600 77046
rect 114940 67153 114968 147086
rect 115032 74534 115060 147154
rect 115112 143336 115164 143342
rect 115112 143278 115164 143284
rect 115124 77858 115152 143278
rect 115112 77852 115164 77858
rect 115112 77794 115164 77800
rect 115216 77110 115244 192743
rect 115308 144294 115336 260986
rect 115572 260908 115624 260914
rect 115572 260850 115624 260856
rect 115480 260092 115532 260098
rect 115480 260034 115532 260040
rect 115388 192772 115440 192778
rect 115388 192714 115440 192720
rect 115296 144288 115348 144294
rect 115296 144230 115348 144236
rect 115296 141908 115348 141914
rect 115296 141850 115348 141856
rect 115204 77104 115256 77110
rect 115204 77046 115256 77052
rect 115216 76702 115244 77046
rect 115204 76696 115256 76702
rect 115204 76638 115256 76644
rect 115032 74506 115244 74534
rect 115216 73846 115244 74506
rect 115204 73840 115256 73846
rect 115204 73782 115256 73788
rect 114926 67144 114982 67153
rect 114926 67079 114982 67088
rect 114940 59362 114968 67079
rect 114928 59356 114980 59362
rect 114928 59298 114980 59304
rect 115216 54602 115244 73782
rect 115308 71126 115336 141850
rect 115400 75818 115428 192714
rect 115492 141982 115520 260034
rect 115584 143070 115612 260850
rect 116676 259480 116728 259486
rect 116676 259422 116728 259428
rect 115848 200592 115900 200598
rect 115848 200534 115900 200540
rect 115664 199572 115716 199578
rect 115664 199514 115716 199520
rect 115572 143064 115624 143070
rect 115572 143006 115624 143012
rect 115480 141976 115532 141982
rect 115480 141918 115532 141924
rect 115676 77110 115704 199514
rect 115756 199096 115808 199102
rect 115756 199038 115808 199044
rect 115664 77104 115716 77110
rect 115768 77081 115796 199038
rect 115664 77046 115716 77052
rect 115754 77072 115810 77081
rect 115754 77007 115810 77016
rect 115388 75812 115440 75818
rect 115388 75754 115440 75760
rect 115860 73001 115888 200534
rect 116306 151056 116362 151065
rect 116306 150991 116362 151000
rect 116216 148436 116268 148442
rect 116216 148378 116268 148384
rect 116124 148232 116176 148238
rect 116124 148174 116176 148180
rect 115940 75132 115992 75138
rect 115940 75074 115992 75080
rect 115846 72992 115902 73001
rect 115846 72927 115902 72936
rect 115296 71120 115348 71126
rect 115296 71062 115348 71068
rect 115204 54596 115256 54602
rect 115204 54538 115256 54544
rect 115952 16574 115980 75074
rect 116136 71058 116164 148174
rect 116228 71641 116256 148378
rect 116214 71632 116270 71641
rect 116214 71567 116270 71576
rect 116124 71052 116176 71058
rect 116124 70994 116176 71000
rect 116320 69630 116348 150991
rect 116400 145716 116452 145722
rect 116400 145658 116452 145664
rect 116412 79801 116440 145658
rect 116492 144628 116544 144634
rect 116492 144570 116544 144576
rect 116398 79792 116454 79801
rect 116398 79727 116454 79736
rect 116504 75138 116532 144570
rect 116688 144226 116716 259422
rect 116780 146198 116808 262686
rect 116872 146266 116900 262754
rect 116860 146260 116912 146266
rect 116860 146202 116912 146208
rect 116768 146192 116820 146198
rect 116768 146134 116820 146140
rect 116858 145752 116914 145761
rect 116858 145687 116914 145696
rect 116768 145512 116820 145518
rect 116768 145454 116820 145460
rect 116676 144220 116728 144226
rect 116676 144162 116728 144168
rect 116584 141840 116636 141846
rect 116584 141782 116636 141788
rect 116492 75132 116544 75138
rect 116492 75074 116544 75080
rect 116308 69624 116360 69630
rect 116308 69566 116360 69572
rect 116596 66026 116624 141782
rect 116780 70378 116808 145454
rect 116872 144362 116900 145687
rect 116964 145450 116992 264046
rect 118332 264036 118384 264042
rect 118332 263978 118384 263984
rect 118056 262472 118108 262478
rect 118056 262414 118108 262420
rect 117962 261216 118018 261225
rect 117962 261151 118018 261160
rect 117976 260953 118004 261151
rect 117962 260944 118018 260953
rect 117962 260879 118018 260888
rect 117228 199300 117280 199306
rect 117228 199242 117280 199248
rect 117136 197192 117188 197198
rect 117136 197134 117188 197140
rect 117044 197056 117096 197062
rect 117044 196998 117096 197004
rect 116952 145444 117004 145450
rect 116952 145386 117004 145392
rect 116860 144356 116912 144362
rect 116860 144298 116912 144304
rect 117056 76974 117084 196998
rect 117044 76968 117096 76974
rect 117044 76910 117096 76916
rect 117148 75041 117176 197134
rect 117240 75546 117268 199242
rect 117320 197396 117372 197402
rect 117320 197338 117372 197344
rect 117332 195430 117360 197338
rect 117686 195936 117742 195945
rect 117686 195871 117742 195880
rect 117320 195424 117372 195430
rect 117320 195366 117372 195372
rect 117700 193798 117728 195871
rect 117688 193792 117740 193798
rect 117688 193734 117740 193740
rect 117686 151192 117742 151201
rect 117686 151127 117742 151136
rect 117596 148504 117648 148510
rect 117596 148446 117648 148452
rect 117504 147008 117556 147014
rect 117504 146950 117556 146956
rect 117228 75540 117280 75546
rect 117228 75482 117280 75488
rect 117134 75032 117190 75041
rect 117134 74967 117190 74976
rect 116768 70372 116820 70378
rect 116768 70314 116820 70320
rect 117516 70242 117544 146950
rect 117608 71738 117636 148446
rect 117700 73778 117728 151127
rect 118068 144770 118096 262414
rect 118240 260840 118292 260846
rect 118240 260782 118292 260788
rect 118148 260024 118200 260030
rect 118148 259966 118200 259972
rect 118056 144764 118108 144770
rect 118056 144706 118108 144712
rect 118160 141710 118188 259966
rect 118148 141704 118200 141710
rect 118148 141646 118200 141652
rect 118252 141302 118280 260782
rect 118344 143138 118372 263978
rect 119712 263968 119764 263974
rect 119712 263910 119764 263916
rect 118424 262948 118476 262954
rect 118424 262890 118476 262896
rect 118332 143132 118384 143138
rect 118332 143074 118384 143080
rect 118436 142050 118464 262890
rect 119620 262404 119672 262410
rect 119620 262346 119672 262352
rect 119528 259956 119580 259962
rect 119528 259898 119580 259904
rect 119436 259752 119488 259758
rect 119436 259694 119488 259700
rect 118608 198756 118660 198762
rect 118608 198698 118660 198704
rect 118516 195220 118568 195226
rect 118516 195162 118568 195168
rect 118424 142044 118476 142050
rect 118424 141986 118476 141992
rect 118240 141296 118292 141302
rect 118240 141238 118292 141244
rect 117780 141024 117832 141030
rect 117780 140966 117832 140972
rect 117792 85542 117820 140966
rect 118148 140616 118200 140622
rect 118148 140558 118200 140564
rect 117872 140548 117924 140554
rect 117872 140490 117924 140496
rect 117780 85536 117832 85542
rect 117780 85478 117832 85484
rect 117884 78878 117912 140490
rect 117964 140276 118016 140282
rect 117964 140218 118016 140224
rect 117872 78872 117924 78878
rect 117872 78814 117924 78820
rect 117976 74118 118004 140218
rect 118056 140208 118108 140214
rect 118056 140150 118108 140156
rect 117964 74112 118016 74118
rect 118068 74089 118096 140150
rect 117964 74054 118016 74060
rect 118054 74080 118110 74089
rect 118054 74015 118110 74024
rect 117688 73772 117740 73778
rect 117688 73714 117740 73720
rect 117596 71732 117648 71738
rect 117596 71674 117648 71680
rect 118160 71534 118188 140558
rect 118528 72593 118556 195162
rect 118620 75342 118648 198698
rect 118884 195492 118936 195498
rect 118884 195434 118936 195440
rect 118792 145988 118844 145994
rect 118792 145930 118844 145936
rect 118700 139664 118752 139670
rect 118700 139606 118752 139612
rect 118712 137970 118740 139606
rect 118700 137964 118752 137970
rect 118700 137906 118752 137912
rect 118804 79150 118832 145930
rect 118896 138145 118924 195434
rect 118976 145920 119028 145926
rect 118976 145862 119028 145868
rect 118882 138136 118938 138145
rect 118882 138071 118938 138080
rect 118792 79144 118844 79150
rect 118792 79086 118844 79092
rect 118988 79082 119016 145862
rect 119068 145852 119120 145858
rect 119068 145794 119120 145800
rect 119080 80986 119108 145794
rect 119448 141438 119476 259694
rect 119540 141506 119568 259898
rect 119632 142798 119660 262346
rect 119724 144702 119752 263910
rect 119804 262608 119856 262614
rect 119804 262550 119856 262556
rect 119712 144696 119764 144702
rect 119712 144638 119764 144644
rect 119712 144424 119764 144430
rect 119712 144366 119764 144372
rect 119620 142792 119672 142798
rect 119620 142734 119672 142740
rect 119528 141500 119580 141506
rect 119528 141442 119580 141448
rect 119436 141432 119488 141438
rect 119436 141374 119488 141380
rect 119252 140412 119304 140418
rect 119252 140354 119304 140360
rect 119068 80980 119120 80986
rect 119068 80922 119120 80928
rect 119264 79694 119292 140354
rect 119344 140072 119396 140078
rect 119344 140014 119396 140020
rect 119252 79688 119304 79694
rect 119252 79630 119304 79636
rect 118976 79076 119028 79082
rect 118976 79018 119028 79024
rect 119356 78946 119384 140014
rect 119344 78940 119396 78946
rect 119344 78882 119396 78888
rect 119724 76838 119752 144366
rect 119816 143478 119844 262550
rect 119896 199436 119948 199442
rect 119896 199378 119948 199384
rect 119804 143472 119856 143478
rect 119804 143414 119856 143420
rect 119802 138952 119858 138961
rect 119802 138887 119858 138896
rect 119712 76832 119764 76838
rect 119712 76774 119764 76780
rect 118608 75336 118660 75342
rect 118608 75278 118660 75284
rect 118514 72584 118570 72593
rect 118514 72519 118570 72528
rect 119816 72418 119844 138887
rect 119908 76809 119936 199378
rect 120000 145654 120028 269078
rect 133156 264110 133184 271866
rect 133144 264104 133196 264110
rect 133144 264046 133196 264052
rect 133328 264104 133380 264110
rect 133328 264046 133380 264052
rect 120908 263900 120960 263906
rect 120908 263842 120960 263848
rect 120816 261112 120868 261118
rect 120816 261054 120868 261060
rect 120632 259616 120684 259622
rect 120632 259558 120684 259564
rect 120448 197464 120500 197470
rect 120448 197406 120500 197412
rect 120460 197198 120488 197406
rect 120448 197192 120500 197198
rect 120448 197134 120500 197140
rect 120644 189038 120672 259558
rect 120724 259548 120776 259554
rect 120724 259490 120776 259496
rect 120632 189032 120684 189038
rect 120632 188974 120684 188980
rect 120448 148572 120500 148578
rect 120448 148514 120500 148520
rect 120356 145784 120408 145790
rect 120356 145726 120408 145732
rect 119988 145648 120040 145654
rect 119988 145590 120040 145596
rect 119986 144800 120042 144809
rect 119986 144735 120042 144744
rect 120000 143614 120028 144735
rect 119988 143608 120040 143614
rect 119988 143550 120040 143556
rect 119988 141568 120040 141574
rect 119988 141510 120040 141516
rect 120000 80714 120028 141510
rect 119988 80708 120040 80714
rect 119988 80650 120040 80656
rect 119894 76800 119950 76809
rect 119894 76735 119950 76744
rect 120368 74390 120396 145726
rect 120356 74384 120408 74390
rect 120356 74326 120408 74332
rect 119804 72412 119856 72418
rect 119804 72354 119856 72360
rect 119816 71806 119844 72354
rect 118700 71800 118752 71806
rect 118700 71742 118752 71748
rect 119804 71800 119856 71806
rect 119804 71742 119856 71748
rect 118148 71528 118200 71534
rect 118148 71470 118200 71476
rect 117504 70236 117556 70242
rect 117504 70178 117556 70184
rect 117320 66972 117372 66978
rect 117320 66914 117372 66920
rect 116584 66020 116636 66026
rect 116584 65962 116636 65968
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 66914
rect 118712 7682 118740 71742
rect 120460 71466 120488 148514
rect 120736 143449 120764 259490
rect 120722 143440 120778 143449
rect 120828 143410 120856 261054
rect 120722 143375 120778 143384
rect 120816 143404 120868 143410
rect 120816 143346 120868 143352
rect 120920 143002 120948 263842
rect 121736 263832 121788 263838
rect 121736 263774 121788 263780
rect 121000 263764 121052 263770
rect 121000 263706 121052 263712
rect 120908 142996 120960 143002
rect 120908 142938 120960 142944
rect 121012 142934 121040 263706
rect 121092 263628 121144 263634
rect 121092 263570 121144 263576
rect 121000 142928 121052 142934
rect 121000 142870 121052 142876
rect 121104 142866 121132 263570
rect 121184 259820 121236 259826
rect 121184 259762 121236 259768
rect 121196 259593 121224 259762
rect 121182 259584 121238 259593
rect 121182 259519 121238 259528
rect 121274 199744 121330 199753
rect 121274 199679 121330 199688
rect 121184 199368 121236 199374
rect 121184 199310 121236 199316
rect 121092 142860 121144 142866
rect 121092 142802 121144 142808
rect 121000 141364 121052 141370
rect 121000 141306 121052 141312
rect 120632 140684 120684 140690
rect 120632 140626 120684 140632
rect 120540 140344 120592 140350
rect 120540 140286 120592 140292
rect 120552 80209 120580 140286
rect 120538 80200 120594 80209
rect 120538 80135 120594 80144
rect 120644 79014 120672 140626
rect 120724 140480 120776 140486
rect 120724 140422 120776 140428
rect 120632 79008 120684 79014
rect 120632 78950 120684 78956
rect 120736 73953 120764 140422
rect 120814 138816 120870 138825
rect 120814 138751 120870 138760
rect 120722 73944 120778 73953
rect 120722 73879 120778 73888
rect 120828 71670 120856 138751
rect 120816 71664 120868 71670
rect 120816 71606 120868 71612
rect 120448 71460 120500 71466
rect 120448 71402 120500 71408
rect 121012 70310 121040 141306
rect 121196 75478 121224 199310
rect 121184 75472 121236 75478
rect 121184 75414 121236 75420
rect 121288 73030 121316 199679
rect 121368 198892 121420 198898
rect 121368 198834 121420 198840
rect 121276 73024 121328 73030
rect 121276 72966 121328 72972
rect 121380 72350 121408 198834
rect 121748 143313 121776 263774
rect 129830 263256 129886 263265
rect 129830 263191 129886 263200
rect 125968 262948 126020 262954
rect 125968 262890 126020 262896
rect 122380 262540 122432 262546
rect 122380 262482 122432 262488
rect 122196 260160 122248 260166
rect 122196 260102 122248 260108
rect 121920 259888 121972 259894
rect 121920 259830 121972 259836
rect 121932 146130 121960 259830
rect 122104 194540 122156 194546
rect 122104 194482 122156 194488
rect 122012 193724 122064 193730
rect 122012 193666 122064 193672
rect 121920 146124 121972 146130
rect 121920 146066 121972 146072
rect 121828 146056 121880 146062
rect 121828 145998 121880 146004
rect 121734 143304 121790 143313
rect 121734 143239 121790 143248
rect 121368 72344 121420 72350
rect 121368 72286 121420 72292
rect 121840 71369 121868 145998
rect 121920 140140 121972 140146
rect 121920 140082 121972 140088
rect 121932 71505 121960 140082
rect 122024 78334 122052 193666
rect 122116 78402 122144 194482
rect 122208 143274 122236 260102
rect 122288 198212 122340 198218
rect 122288 198154 122340 198160
rect 122196 143268 122248 143274
rect 122196 143210 122248 143216
rect 122194 139088 122250 139097
rect 122194 139023 122250 139032
rect 122104 78396 122156 78402
rect 122104 78338 122156 78344
rect 122012 78328 122064 78334
rect 122012 78270 122064 78276
rect 121918 71496 121974 71505
rect 121918 71431 121974 71440
rect 121826 71360 121882 71369
rect 121460 71324 121512 71330
rect 121826 71295 121882 71304
rect 121460 71266 121512 71272
rect 121472 70990 121500 71266
rect 121460 70984 121512 70990
rect 121460 70926 121512 70932
rect 121000 70304 121052 70310
rect 121000 70246 121052 70252
rect 120080 67108 120132 67114
rect 120080 67050 120132 67056
rect 120092 16574 120120 67050
rect 120092 16546 120672 16574
rect 118700 7676 118752 7682
rect 118700 7618 118752 7624
rect 119896 7676 119948 7682
rect 119896 7618 119948 7624
rect 118792 4140 118844 4146
rect 118792 4082 118844 4088
rect 118804 480 118832 4082
rect 119908 480 119936 7618
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 121472 4146 121500 70926
rect 122208 70106 122236 139023
rect 122300 80918 122328 198154
rect 122392 144566 122420 262482
rect 124312 260840 124364 260846
rect 124312 260782 124364 260788
rect 124324 259978 124352 260782
rect 124862 260536 124918 260545
rect 124862 260471 124918 260480
rect 124876 259978 124904 260471
rect 125980 259978 126008 262890
rect 128728 262676 128780 262682
rect 128728 262618 128780 262624
rect 127716 262404 127768 262410
rect 127716 262346 127768 262352
rect 127072 262336 127124 262342
rect 127072 262278 127124 262284
rect 126842 260092 126894 260098
rect 126842 260034 126894 260040
rect 124324 259950 124660 259978
rect 124876 259950 125212 259978
rect 125980 259950 126316 259978
rect 126854 259964 126882 260034
rect 127084 259978 127112 262278
rect 127622 261216 127678 261225
rect 127622 261151 127678 261160
rect 127636 260953 127664 261151
rect 127622 260944 127678 260953
rect 127622 260879 127678 260888
rect 127728 259978 127756 262346
rect 128740 259978 128768 262618
rect 129280 262472 129332 262478
rect 129280 262414 129332 262420
rect 129292 259978 129320 262414
rect 129844 261458 129872 263191
rect 132040 263016 132092 263022
rect 132040 262958 132092 262964
rect 131120 262948 131172 262954
rect 131120 262890 131172 262896
rect 131764 262948 131816 262954
rect 131764 262890 131816 262896
rect 131132 262818 131160 262890
rect 131120 262812 131172 262818
rect 131120 262754 131172 262760
rect 131120 262608 131172 262614
rect 131120 262550 131172 262556
rect 129832 261452 129884 261458
rect 129832 261394 129884 261400
rect 129844 259978 129872 261394
rect 131132 261322 131160 262550
rect 131120 261316 131172 261322
rect 131120 261258 131172 261264
rect 130384 261044 130436 261050
rect 130384 260986 130436 260992
rect 130396 259978 130424 260986
rect 131132 259978 131160 261258
rect 131776 259978 131804 262890
rect 132052 260914 132080 262958
rect 133236 261112 133288 261118
rect 133236 261054 133288 261060
rect 132040 260908 132092 260914
rect 132040 260850 132092 260856
rect 132052 259978 132080 260850
rect 133248 260370 133276 261054
rect 133236 260364 133288 260370
rect 133236 260306 133288 260312
rect 133248 259978 133276 260306
rect 127084 259950 127420 259978
rect 127728 259950 127972 259978
rect 128740 259950 129076 259978
rect 129292 259950 129628 259978
rect 129844 259950 130180 259978
rect 130396 259950 130732 259978
rect 131132 259950 131284 259978
rect 131776 259950 131836 259978
rect 132052 259950 132388 259978
rect 132940 259950 133276 259978
rect 133340 259978 133368 264046
rect 134248 264036 134300 264042
rect 134248 263978 134300 263984
rect 133970 261080 134026 261089
rect 133970 261015 134026 261024
rect 133984 259978 134012 261015
rect 134260 259978 134288 263978
rect 134536 262750 134564 324294
rect 134616 298172 134668 298178
rect 134616 298114 134668 298120
rect 134628 264042 134656 298114
rect 134616 264036 134668 264042
rect 134616 263978 134668 263984
rect 134524 262744 134576 262750
rect 134524 262686 134576 262692
rect 134800 262744 134852 262750
rect 134800 262686 134852 262692
rect 134812 259978 134840 262686
rect 135272 260234 135300 351902
rect 135904 311908 135956 311914
rect 135904 311850 135956 311856
rect 135916 265169 135944 311850
rect 137284 286340 137336 286346
rect 137284 286282 137336 286288
rect 137296 267734 137324 286282
rect 137204 267706 137324 267734
rect 135902 265160 135958 265169
rect 135902 265095 135958 265104
rect 135260 260228 135312 260234
rect 135260 260170 135312 260176
rect 135916 259978 135944 265095
rect 137204 263702 137232 267706
rect 137836 267028 137888 267034
rect 137836 266970 137888 266976
rect 137848 263974 137876 266970
rect 137836 263968 137888 263974
rect 137836 263910 137888 263916
rect 137192 263696 137244 263702
rect 137192 263638 137244 263644
rect 136226 260228 136278 260234
rect 136226 260170 136278 260176
rect 133340 259950 133492 259978
rect 133984 259964 134044 259978
rect 133984 259950 134058 259964
rect 134260 259950 134596 259978
rect 134812 259950 135148 259978
rect 135700 259950 135944 259978
rect 136238 259964 136266 260170
rect 137204 259978 137232 263638
rect 137468 263560 137520 263566
rect 137468 263502 137520 263508
rect 137480 260953 137508 263502
rect 137466 260944 137522 260953
rect 137466 260879 137522 260888
rect 136804 259950 137232 259978
rect 134030 259706 134058 259950
rect 137480 259842 137508 260879
rect 137356 259814 137508 259842
rect 137848 259842 137876 263910
rect 138676 262993 138704 430578
rect 138756 418192 138808 418198
rect 138756 418134 138808 418140
rect 138768 265033 138796 418134
rect 139412 267734 139440 484366
rect 140044 470620 140096 470626
rect 140044 470562 140096 470568
rect 140056 267734 140084 470562
rect 140780 280832 140832 280838
rect 140780 280774 140832 280780
rect 139412 267706 139716 267734
rect 140056 267706 140360 267734
rect 138754 265024 138810 265033
rect 138754 264959 138810 264968
rect 138662 262984 138718 262993
rect 138662 262919 138718 262928
rect 138676 259978 138704 262919
rect 138460 259950 138704 259978
rect 138768 259978 138796 264959
rect 139400 264308 139452 264314
rect 139400 264250 139452 264256
rect 139412 263906 139440 264250
rect 139400 263900 139452 263906
rect 139400 263842 139452 263848
rect 139412 259978 139440 263842
rect 139688 260030 139716 267706
rect 140332 262857 140360 267706
rect 140318 262848 140374 262857
rect 140318 262783 140374 262792
rect 139676 260024 139728 260030
rect 138768 259950 139012 259978
rect 139412 259950 139564 259978
rect 140332 259978 140360 262783
rect 139728 259972 140116 259978
rect 139676 259966 140116 259972
rect 139688 259950 140116 259966
rect 140332 259950 140668 259978
rect 140792 259962 140820 280774
rect 142356 267734 142384 590650
rect 142804 563100 142856 563106
rect 142804 563042 142856 563048
rect 142816 267734 142844 563042
rect 142896 524476 142948 524482
rect 142896 524418 142948 524424
rect 142264 267706 142384 267734
rect 142632 267706 142844 267734
rect 140964 265736 141016 265742
rect 140964 265678 141016 265684
rect 140976 263770 141004 265678
rect 140964 263764 141016 263770
rect 140964 263706 141016 263712
rect 140976 259978 141004 263706
rect 142158 262440 142214 262449
rect 142158 262375 142214 262384
rect 142172 259978 142200 262375
rect 142264 260137 142292 267706
rect 142632 263838 142660 267706
rect 142620 263832 142672 263838
rect 142620 263774 142672 263780
rect 142250 260128 142306 260137
rect 142250 260063 142306 260072
rect 142632 259978 142660 263774
rect 142908 262449 142936 524418
rect 142894 262440 142950 262449
rect 142894 262375 142950 262384
rect 143644 260273 143672 616830
rect 144184 576904 144236 576910
rect 144184 576846 144236 576852
rect 144196 262585 144224 576846
rect 145564 289128 145616 289134
rect 145564 289070 145616 289076
rect 144920 282192 144972 282198
rect 144920 282134 144972 282140
rect 144182 262576 144238 262585
rect 144182 262511 144238 262520
rect 143630 260264 143686 260273
rect 143630 260199 143686 260208
rect 143400 260128 143456 260137
rect 143400 260063 143456 260072
rect 140780 259956 140832 259962
rect 139688 259901 139716 259950
rect 140976 259950 141220 259978
rect 141436 259962 141772 259978
rect 141424 259956 141772 259962
rect 140780 259898 140832 259904
rect 141476 259950 141772 259956
rect 142172 259950 142324 259978
rect 142632 259950 142876 259978
rect 143414 259964 143442 260063
rect 144196 259978 144224 262511
rect 144504 260264 144560 260273
rect 144504 260199 144560 260208
rect 143980 259950 144224 259978
rect 144518 259964 144546 260199
rect 144932 260001 144960 282134
rect 145576 263809 145604 289070
rect 146208 268388 146260 268394
rect 146208 268330 146260 268336
rect 146220 263945 146248 268330
rect 146206 263936 146262 263945
rect 146206 263871 146262 263880
rect 145562 263800 145618 263809
rect 145562 263735 145618 263744
rect 144918 259992 144974 260001
rect 145576 259978 145604 263735
rect 146220 260250 146248 263871
rect 146174 260222 146248 260250
rect 144974 259950 145084 259978
rect 145576 259950 145636 259978
rect 146174 259964 146202 260222
rect 146312 259978 146340 696934
rect 146944 683188 146996 683194
rect 146944 683130 146996 683136
rect 146956 262721 146984 683130
rect 147680 283620 147732 283626
rect 147680 283562 147732 283568
rect 146942 262712 146998 262721
rect 146942 262647 146998 262656
rect 146956 259978 146984 262647
rect 147692 260273 147720 283562
rect 147772 269816 147824 269822
rect 147772 269758 147824 269764
rect 147678 260264 147734 260273
rect 147678 260199 147734 260208
rect 147784 259978 147812 269758
rect 148336 267734 148364 700266
rect 149704 345092 149756 345098
rect 149704 345034 149756 345040
rect 149060 287700 149112 287706
rect 149060 287642 149112 287648
rect 148336 267706 148640 267734
rect 148612 263673 148640 267706
rect 148598 263664 148654 263673
rect 148598 263599 148654 263608
rect 148368 260264 148424 260273
rect 148368 260199 148424 260208
rect 146312 259950 146740 259978
rect 146956 259950 147292 259978
rect 147784 259950 147844 259978
rect 144918 259927 144974 259936
rect 141424 259898 141476 259904
rect 144932 259867 144960 259927
rect 146312 259894 146340 259950
rect 146300 259888 146352 259894
rect 137848 259814 137908 259842
rect 147784 259842 147812 259950
rect 146300 259830 146352 259836
rect 147692 259826 147812 259842
rect 147680 259820 147812 259826
rect 147732 259814 147812 259820
rect 147680 259762 147732 259768
rect 148138 259720 148194 259729
rect 134030 259692 134380 259706
rect 134044 259690 134380 259692
rect 134044 259684 134392 259690
rect 134044 259678 134340 259684
rect 148382 259706 148410 260199
rect 148612 259978 148640 263599
rect 149072 260273 149100 287642
rect 149152 271176 149204 271182
rect 149152 271118 149204 271124
rect 149058 260264 149114 260273
rect 149058 260199 149114 260208
rect 149164 259978 149192 271118
rect 149716 264382 149744 345034
rect 150438 284336 150494 284345
rect 150438 284271 150494 284280
rect 149704 264376 149756 264382
rect 149704 264318 149756 264324
rect 150452 263498 150480 284271
rect 151084 275324 151136 275330
rect 151084 275266 151136 275272
rect 151096 263634 151124 275266
rect 151912 273284 151964 273290
rect 151912 273226 151964 273232
rect 151924 267734 151952 273226
rect 151924 267706 152412 267734
rect 151084 263628 151136 263634
rect 151084 263570 151136 263576
rect 150440 263492 150492 263498
rect 150440 263434 150492 263440
rect 150530 263120 150586 263129
rect 150530 263055 150586 263064
rect 150024 260264 150080 260273
rect 150024 260199 150080 260208
rect 148612 259950 148948 259978
rect 149164 259950 149500 259978
rect 150038 259964 150066 260199
rect 150544 259978 150572 263055
rect 151096 259978 151124 263570
rect 151360 263492 151412 263498
rect 151360 263434 151412 263440
rect 151372 259978 151400 263434
rect 152188 262540 152240 262546
rect 152188 262482 152240 262488
rect 152200 259978 152228 262482
rect 152384 259978 152412 267706
rect 152476 262546 152504 700334
rect 153212 262750 153240 702406
rect 157340 700868 157392 700874
rect 157340 700810 157392 700816
rect 155960 700800 156012 700806
rect 155960 700742 156012 700748
rect 154580 700664 154632 700670
rect 154580 700606 154632 700612
rect 153292 700460 153344 700466
rect 153292 700402 153344 700408
rect 153200 262744 153252 262750
rect 153200 262686 153252 262692
rect 152464 262540 152516 262546
rect 152464 262482 152516 262488
rect 153304 259978 153332 700402
rect 153382 276040 153438 276049
rect 153382 275975 153438 275984
rect 153396 267734 153424 275975
rect 153396 267706 154068 267734
rect 153844 262676 153896 262682
rect 153844 262618 153896 262624
rect 153856 259978 153884 262618
rect 154040 259978 154068 267706
rect 154592 259978 154620 700606
rect 155868 262608 155920 262614
rect 155868 262550 155920 262556
rect 155880 259978 155908 262550
rect 155972 260273 156000 700742
rect 156050 277536 156106 277545
rect 156050 277471 156106 277480
rect 155958 260264 156014 260273
rect 155958 260199 156014 260208
rect 150544 259950 150604 259978
rect 151096 259950 151156 259978
rect 151372 259950 151708 259978
rect 152200 259950 152260 259978
rect 152384 259950 152812 259978
rect 153304 259950 153364 259978
rect 153856 259950 153916 259978
rect 154040 259950 154468 259978
rect 154592 259950 155264 259978
rect 155572 259950 155908 259978
rect 156064 259978 156092 277471
rect 157156 262540 157208 262546
rect 157156 262482 157208 262488
rect 156648 260264 156704 260273
rect 156648 260199 156704 260208
rect 156064 259950 156124 259978
rect 149256 259865 149284 259950
rect 149242 259856 149298 259865
rect 153304 259842 153332 259950
rect 149242 259791 149298 259800
rect 153212 259814 153332 259842
rect 153212 259758 153240 259814
rect 148194 259692 148410 259706
rect 153200 259752 153252 259758
rect 153200 259694 153252 259700
rect 148194 259678 148396 259692
rect 148138 259655 148194 259664
rect 134340 259626 134392 259632
rect 155236 259593 155264 259950
rect 156662 259706 156690 260199
rect 157168 259978 157196 262482
rect 157352 260234 157380 700810
rect 160744 700732 160796 700738
rect 160744 700674 160796 700680
rect 157432 450560 157484 450566
rect 157432 450502 157484 450508
rect 157340 260228 157392 260234
rect 157340 260170 157392 260176
rect 157444 259978 157472 450502
rect 160100 279472 160152 279478
rect 160100 279414 160152 279420
rect 158720 269136 158772 269142
rect 158720 269078 158772 269084
rect 158732 267734 158760 269078
rect 158732 267706 159588 267734
rect 158720 264240 158772 264246
rect 158720 264182 158772 264188
rect 158732 263634 158760 264182
rect 158720 263628 158772 263634
rect 158720 263570 158772 263576
rect 159364 263628 159416 263634
rect 159364 263570 159416 263576
rect 158720 262744 158772 262750
rect 158720 262686 158772 262692
rect 158732 260953 158760 262686
rect 158718 260944 158774 260953
rect 158718 260879 158774 260888
rect 158306 260228 158358 260234
rect 158306 260170 158358 260176
rect 158318 259978 158346 260170
rect 158732 259978 158760 260879
rect 159376 259978 159404 263570
rect 159560 259978 159588 267706
rect 160112 260273 160140 279414
rect 160756 267734 160784 700674
rect 162216 700596 162268 700602
rect 162216 700538 162268 700544
rect 162124 700528 162176 700534
rect 162124 700470 162176 700476
rect 161480 683256 161532 683262
rect 161480 683198 161532 683204
rect 160756 267706 160876 267734
rect 160848 265305 160876 267706
rect 160834 265296 160890 265305
rect 160834 265231 160890 265240
rect 160098 260264 160154 260273
rect 160098 260199 160154 260208
rect 160848 259978 160876 265231
rect 161492 260273 161520 683198
rect 162136 267734 162164 700470
rect 162044 267706 162164 267734
rect 162044 262721 162072 267706
rect 162228 265169 162256 700538
rect 163504 670744 163556 670750
rect 163504 670686 163556 670692
rect 162214 265160 162270 265169
rect 162214 265095 162270 265104
rect 162030 262712 162086 262721
rect 162030 262647 162086 262656
rect 161064 260264 161120 260273
rect 161064 260199 161120 260208
rect 161478 260264 161534 260273
rect 161478 260199 161534 260208
rect 157168 259950 157228 259978
rect 157444 259950 158116 259978
rect 158318 259964 158668 259978
rect 158332 259950 158668 259964
rect 158732 259950 158884 259978
rect 159376 259950 159436 259978
rect 159560 259950 159988 259978
rect 160540 259950 160876 259978
rect 158088 259826 158116 259950
rect 158076 259820 158128 259826
rect 158076 259762 158128 259768
rect 158640 259758 158668 259950
rect 161078 259842 161106 260199
rect 162044 259978 162072 262647
rect 162228 260250 162256 265095
rect 163516 264994 163544 670686
rect 163596 656940 163648 656946
rect 163596 656882 163648 656888
rect 163504 264988 163556 264994
rect 163504 264930 163556 264936
rect 163410 263120 163466 263129
rect 163410 263055 163466 263064
rect 163424 262449 163452 263055
rect 163410 262440 163466 262449
rect 163410 262375 163466 262384
rect 161644 259950 162072 259978
rect 162182 260222 162256 260250
rect 162720 260264 162776 260273
rect 162182 259964 162210 260222
rect 162720 260199 162776 260208
rect 162734 259978 162762 260199
rect 162858 259992 162914 260001
rect 162734 259964 162858 259978
rect 162748 259950 162858 259964
rect 163424 259978 163452 262375
rect 163300 259950 163452 259978
rect 163516 259978 163544 264930
rect 163608 263129 163636 656882
rect 164240 632120 164292 632126
rect 164240 632062 164292 632068
rect 163594 263120 163650 263129
rect 163594 263055 163650 263064
rect 164252 259978 164280 632062
rect 164884 618316 164936 618322
rect 164884 618258 164936 618264
rect 164896 265033 164924 618258
rect 164976 605872 165028 605878
rect 164976 605814 165028 605820
rect 164882 265024 164938 265033
rect 164882 264959 164938 264968
rect 164988 262585 165016 605814
rect 165620 579692 165672 579698
rect 165620 579634 165672 579640
rect 165158 265024 165214 265033
rect 165158 264959 165214 264968
rect 164974 262576 165030 262585
rect 164974 262511 165030 262520
rect 164988 260250 165016 262511
rect 164942 260222 165016 260250
rect 163516 259950 163852 259978
rect 164252 259962 164740 259978
rect 164942 259964 164970 260222
rect 165172 259978 165200 264959
rect 165632 259978 165660 579634
rect 167644 565888 167696 565894
rect 167644 565830 167696 565836
rect 166264 553444 166316 553450
rect 166264 553386 166316 553392
rect 166276 262750 166304 553386
rect 167000 527196 167052 527202
rect 167000 527138 167052 527144
rect 166264 262744 166316 262750
rect 166264 262686 166316 262692
rect 166276 259978 166304 262686
rect 167012 260234 167040 527138
rect 167656 267734 167684 565830
rect 167736 501016 167788 501022
rect 167736 500958 167788 500964
rect 167564 267706 167684 267734
rect 167748 267734 167776 500958
rect 169772 450566 169800 702406
rect 202800 700806 202828 703520
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 182824 643136 182876 643142
rect 182824 643078 182876 643084
rect 181444 536852 181496 536858
rect 181444 536794 181496 536800
rect 180064 510672 180116 510678
rect 180064 510614 180116 510620
rect 170404 462392 170456 462398
rect 170404 462334 170456 462340
rect 169760 450560 169812 450566
rect 169760 450502 169812 450508
rect 169760 422340 169812 422346
rect 169760 422282 169812 422288
rect 169024 271244 169076 271250
rect 169024 271186 169076 271192
rect 169036 267734 169064 271186
rect 167748 267706 167868 267734
rect 169036 267706 169156 267734
rect 167564 265441 167592 267706
rect 167550 265432 167606 265441
rect 167550 265367 167606 265376
rect 167000 260228 167052 260234
rect 167000 260170 167052 260176
rect 167564 259978 167592 265367
rect 167840 262818 167868 267706
rect 169128 265062 169156 267706
rect 169208 265668 169260 265674
rect 169208 265610 169260 265616
rect 169116 265056 169168 265062
rect 169116 264998 169168 265004
rect 167828 262812 167880 262818
rect 167828 262754 167880 262760
rect 167690 260228 167742 260234
rect 167690 260170 167742 260176
rect 167702 260098 167730 260170
rect 167690 260092 167742 260098
rect 167690 260034 167742 260040
rect 164252 259956 164752 259962
rect 164252 259950 164700 259956
rect 162858 259927 162914 259936
rect 165172 259950 165508 259978
rect 165632 259950 166212 259978
rect 166276 259950 166612 259978
rect 167164 259950 167592 259978
rect 167702 259964 167730 260034
rect 167840 259978 167868 262754
rect 169128 259978 169156 264998
rect 169220 260302 169248 265610
rect 169208 260296 169260 260302
rect 169208 260238 169260 260244
rect 167840 259950 168268 259978
rect 168820 259950 169156 259978
rect 169220 259978 169248 260238
rect 169772 260234 169800 422282
rect 170220 265396 170272 265402
rect 170220 265338 170272 265344
rect 169760 260228 169812 260234
rect 169760 260170 169812 260176
rect 170232 259978 170260 265338
rect 170416 265130 170444 462334
rect 178684 456816 178736 456822
rect 178684 456758 178736 456764
rect 170496 448588 170548 448594
rect 170496 448530 170548 448536
rect 170508 265402 170536 448530
rect 171784 409896 171836 409902
rect 171784 409838 171836 409844
rect 170496 265396 170548 265402
rect 170496 265338 170548 265344
rect 171692 265260 171744 265266
rect 171692 265202 171744 265208
rect 170404 265124 170456 265130
rect 170404 265066 170456 265072
rect 170680 265124 170732 265130
rect 170680 265066 170732 265072
rect 170692 259978 170720 265066
rect 171002 260228 171054 260234
rect 171002 260170 171054 260176
rect 169220 259950 169372 259978
rect 169924 259950 170260 259978
rect 170476 259950 170720 259978
rect 171014 259964 171042 260170
rect 171704 259978 171732 265202
rect 171796 265198 171824 409838
rect 171876 397520 171928 397526
rect 171876 397462 171928 397468
rect 171888 265266 171916 397462
rect 173900 318844 173952 318850
rect 173900 318786 173952 318792
rect 173164 273964 173216 273970
rect 173164 273906 173216 273912
rect 172704 268456 172756 268462
rect 172704 268398 172756 268404
rect 171876 265260 171928 265266
rect 171876 265202 171928 265208
rect 171784 265192 171836 265198
rect 171784 265134 171836 265140
rect 171580 259950 171732 259978
rect 171796 259978 171824 265134
rect 172716 263770 172744 268398
rect 173176 267734 173204 273906
rect 173176 267706 173480 267734
rect 173452 265470 173480 267706
rect 173440 265464 173492 265470
rect 173440 265406 173492 265412
rect 173256 264376 173308 264382
rect 173256 264318 173308 264324
rect 172704 263764 172756 263770
rect 172704 263706 172756 263712
rect 172716 260250 172744 263706
rect 173268 263702 173296 264318
rect 173256 263696 173308 263702
rect 173256 263638 173308 263644
rect 173268 260250 173296 263638
rect 172670 260222 172744 260250
rect 173222 260222 173296 260250
rect 171796 259950 172132 259978
rect 172670 259964 172698 260222
rect 173222 259964 173250 260222
rect 173452 259978 173480 265406
rect 173912 259978 173940 318786
rect 175924 305040 175976 305046
rect 175924 304982 175976 304988
rect 174544 292596 174596 292602
rect 174544 292538 174596 292544
rect 174556 265606 174584 292538
rect 175936 267734 175964 304982
rect 175844 267706 175964 267734
rect 174544 265600 174596 265606
rect 174544 265542 174596 265548
rect 174556 259978 174584 265542
rect 175844 265334 175872 267706
rect 175924 266416 175976 266422
rect 175924 266358 175976 266364
rect 175832 265328 175884 265334
rect 175832 265270 175884 265276
rect 175844 259978 175872 265270
rect 175936 260166 175964 266358
rect 178696 264314 178724 456758
rect 180076 265742 180104 510614
rect 181456 280838 181484 536794
rect 182836 282198 182864 643078
rect 188344 630692 188396 630698
rect 188344 630634 188396 630640
rect 185584 404388 185636 404394
rect 185584 404330 185636 404336
rect 182824 282192 182876 282198
rect 182824 282134 182876 282140
rect 181444 280832 181496 280838
rect 181444 280774 181496 280780
rect 185596 267034 185624 404330
rect 188356 289134 188384 630634
rect 196624 378208 196676 378214
rect 196624 378150 196676 378156
rect 188344 289128 188396 289134
rect 188344 289070 188396 289076
rect 196636 286346 196664 378150
rect 196624 286340 196676 286346
rect 196624 286282 196676 286288
rect 186688 273964 186740 273970
rect 186688 273906 186740 273912
rect 186700 273290 186728 273906
rect 186688 273284 186740 273290
rect 186688 273226 186740 273232
rect 187148 273284 187200 273290
rect 187148 273226 187200 273232
rect 185584 267028 185636 267034
rect 185584 266970 185636 266976
rect 180064 265736 180116 265742
rect 180064 265678 180116 265684
rect 178684 264308 178736 264314
rect 178684 264250 178736 264256
rect 177396 263084 177448 263090
rect 177396 263026 177448 263032
rect 177408 261118 177436 263026
rect 179052 262880 179104 262886
rect 179052 262822 179104 262828
rect 179236 262880 179288 262886
rect 179236 262822 179288 262828
rect 179064 261390 179092 262822
rect 179052 261384 179104 261390
rect 179052 261326 179104 261332
rect 177948 261248 178000 261254
rect 177948 261190 178000 261196
rect 177396 261112 177448 261118
rect 177396 261054 177448 261060
rect 176200 260976 176252 260982
rect 176200 260918 176252 260924
rect 175924 260160 175976 260166
rect 175924 260102 175976 260108
rect 173452 259950 173788 259978
rect 173912 259950 174492 259978
rect 174556 259950 174892 259978
rect 175444 259950 175872 259978
rect 175936 259978 175964 260102
rect 176212 259978 176240 260918
rect 177408 259978 177436 261054
rect 177960 260438 177988 261190
rect 177948 260432 178000 260438
rect 177948 260374 178000 260380
rect 178684 260432 178736 260438
rect 178684 260374 178736 260380
rect 177960 259978 177988 260374
rect 178696 260302 178724 260374
rect 178684 260296 178736 260302
rect 178684 260238 178736 260244
rect 178500 260024 178552 260030
rect 175936 259950 175996 259978
rect 176212 259950 176548 259978
rect 177100 259950 177436 259978
rect 177652 259950 177988 259978
rect 178204 259972 178500 259978
rect 179064 259978 179092 261326
rect 178204 259966 178552 259972
rect 178204 259964 178540 259966
rect 178190 259950 178540 259964
rect 178756 259950 179092 259978
rect 179248 259978 179276 262822
rect 181444 262472 181496 262478
rect 181444 262414 181496 262420
rect 181168 262268 181220 262274
rect 181168 262210 181220 262216
rect 180708 261180 180760 261186
rect 180708 261122 180760 261128
rect 179696 260500 179748 260506
rect 179696 260442 179748 260448
rect 179248 259950 179308 259978
rect 164700 259898 164752 259904
rect 166184 259894 166212 259950
rect 166172 259888 166224 259894
rect 161202 259856 161258 259865
rect 161078 259828 161202 259842
rect 161092 259814 161202 259828
rect 166172 259830 166224 259836
rect 161202 259791 161258 259800
rect 158628 259752 158680 259758
rect 156878 259720 156934 259729
rect 156662 259692 156878 259706
rect 156676 259678 156878 259692
rect 158628 259694 158680 259700
rect 156878 259655 156934 259664
rect 123298 259584 123354 259593
rect 123942 259584 123998 259593
rect 123354 259542 123556 259570
rect 123298 259519 123354 259528
rect 155222 259584 155278 259593
rect 123998 259542 124108 259570
rect 125612 259554 125764 259570
rect 125600 259548 125764 259554
rect 123942 259519 123998 259528
rect 125652 259542 125764 259548
rect 128372 259542 128524 259570
rect 125600 259490 125652 259496
rect 128372 259486 128400 259542
rect 174464 259554 174492 259950
rect 178190 259706 178218 259950
rect 179708 259758 179736 260442
rect 180720 259978 180748 261122
rect 181180 259978 181208 262210
rect 181260 260568 181312 260574
rect 181260 260510 181312 260516
rect 180412 259950 180748 259978
rect 180964 259950 181208 259978
rect 181272 259826 181300 260510
rect 181350 260128 181406 260137
rect 181350 260063 181406 260072
rect 181260 259820 181312 259826
rect 181260 259762 181312 259768
rect 178052 259692 178218 259706
rect 179696 259752 179748 259758
rect 180156 259752 180208 259758
rect 179696 259694 179748 259700
rect 179860 259700 180156 259706
rect 181364 259729 181392 260063
rect 181456 259978 181484 262414
rect 184756 262404 184808 262410
rect 184756 262346 184808 262352
rect 182916 262336 182968 262342
rect 182916 262278 182968 262284
rect 181996 261044 182048 261050
rect 181996 260986 182048 260992
rect 181628 260024 181680 260030
rect 181456 259950 181516 259978
rect 181628 259966 181680 259972
rect 181720 260024 181772 260030
rect 181720 259966 181772 259972
rect 182008 259978 182036 260986
rect 182928 259978 182956 262278
rect 184020 260908 184072 260914
rect 184020 260850 184072 260856
rect 184032 259978 184060 260850
rect 181640 259826 181668 259966
rect 181628 259820 181680 259826
rect 181628 259762 181680 259768
rect 179860 259694 180208 259700
rect 181350 259720 181406 259729
rect 178052 259678 178204 259692
rect 179860 259678 180196 259694
rect 178052 259622 178080 259678
rect 181350 259655 181406 259664
rect 181732 259622 181760 259966
rect 182008 259950 182068 259978
rect 182620 259950 182956 259978
rect 183724 259950 184060 259978
rect 184664 260024 184716 260030
rect 184664 259966 184716 259972
rect 184768 259978 184796 262346
rect 184572 259752 184624 259758
rect 184276 259700 184572 259706
rect 184276 259694 184624 259700
rect 184276 259678 184612 259694
rect 184676 259690 184704 259966
rect 184768 259950 184828 259978
rect 184664 259684 184716 259690
rect 184664 259626 184716 259632
rect 178040 259616 178092 259622
rect 178040 259558 178092 259564
rect 181720 259616 181772 259622
rect 185674 259584 185730 259593
rect 181720 259558 181772 259564
rect 183172 259554 183508 259570
rect 155222 259519 155278 259528
rect 174452 259548 174504 259554
rect 183172 259548 183520 259554
rect 183172 259542 183468 259548
rect 174452 259490 174504 259496
rect 185380 259542 185674 259570
rect 185674 259519 185730 259528
rect 183468 259490 183520 259496
rect 128360 259480 128412 259486
rect 122838 259448 122894 259457
rect 122894 259406 123004 259434
rect 128360 259422 128412 259428
rect 122838 259383 122894 259392
rect 122562 209672 122618 209681
rect 122562 209607 122618 209616
rect 122576 205601 122604 209607
rect 122562 205592 122618 205601
rect 122562 205527 122618 205536
rect 122562 201104 122618 201113
rect 122562 201039 122618 201048
rect 122576 200190 122604 201039
rect 124034 200696 124090 200705
rect 124034 200631 124090 200640
rect 131948 200660 132000 200666
rect 122748 200524 122800 200530
rect 122748 200466 122800 200472
rect 122564 200184 122616 200190
rect 122564 200126 122616 200132
rect 122472 198348 122524 198354
rect 122472 198290 122524 198296
rect 122380 144560 122432 144566
rect 122380 144502 122432 144508
rect 122378 140312 122434 140321
rect 122378 140247 122434 140256
rect 122392 132569 122420 140247
rect 122378 132560 122434 132569
rect 122378 132495 122434 132504
rect 122378 132424 122434 132433
rect 122378 132359 122434 132368
rect 122392 122913 122420 132359
rect 122378 122904 122434 122913
rect 122378 122839 122434 122848
rect 122378 122768 122434 122777
rect 122378 122703 122434 122712
rect 122392 113257 122420 122703
rect 122378 113248 122434 113257
rect 122378 113183 122434 113192
rect 122378 113112 122434 113121
rect 122378 113047 122434 113056
rect 122392 103601 122420 113047
rect 122378 103592 122434 103601
rect 122378 103527 122434 103536
rect 122378 103456 122434 103465
rect 122378 103391 122434 103400
rect 122392 93945 122420 103391
rect 122378 93936 122434 93945
rect 122378 93871 122434 93880
rect 122378 93800 122434 93809
rect 122378 93735 122434 93744
rect 122392 84289 122420 93735
rect 122378 84280 122434 84289
rect 122378 84215 122434 84224
rect 122378 84144 122434 84153
rect 122378 84079 122434 84088
rect 122288 80912 122340 80918
rect 122288 80854 122340 80860
rect 122392 74633 122420 84079
rect 122484 79218 122512 198290
rect 122562 196072 122618 196081
rect 122562 196007 122618 196016
rect 122576 190505 122604 196007
rect 122656 195968 122708 195974
rect 122656 195910 122708 195916
rect 122562 190496 122618 190505
rect 122562 190431 122618 190440
rect 122562 190360 122618 190369
rect 122562 190295 122618 190304
rect 122576 180849 122604 190295
rect 122562 180840 122618 180849
rect 122562 180775 122618 180784
rect 122564 144492 122616 144498
rect 122564 144434 122616 144440
rect 122472 79212 122524 79218
rect 122472 79154 122524 79160
rect 122378 74624 122434 74633
rect 122378 74559 122434 74568
rect 122196 70100 122248 70106
rect 122196 70042 122248 70048
rect 122576 69766 122604 144434
rect 122668 72894 122696 195910
rect 122760 75410 122788 200466
rect 123300 198484 123352 198490
rect 123300 198426 123352 198432
rect 123208 193656 123260 193662
rect 123208 193598 123260 193604
rect 122838 149016 122894 149025
rect 122838 148951 122894 148960
rect 122852 139602 122880 148951
rect 123116 148844 123168 148850
rect 123116 148786 123168 148792
rect 122840 139596 122892 139602
rect 122840 139538 122892 139544
rect 123024 81116 123076 81122
rect 123024 81058 123076 81064
rect 123036 80918 123064 81058
rect 123024 80912 123076 80918
rect 123024 80854 123076 80860
rect 123024 78532 123076 78538
rect 123024 78474 123076 78480
rect 123036 77994 123064 78474
rect 123024 77988 123076 77994
rect 123024 77930 123076 77936
rect 122748 75404 122800 75410
rect 122748 75346 122800 75352
rect 122656 72888 122708 72894
rect 122656 72830 122708 72836
rect 123128 71330 123156 148786
rect 123220 78130 123248 193598
rect 123312 79286 123340 198426
rect 123392 196512 123444 196518
rect 123392 196454 123444 196460
rect 123300 79280 123352 79286
rect 123300 79222 123352 79228
rect 123208 78124 123260 78130
rect 123208 78066 123260 78072
rect 123404 77926 123432 196454
rect 124048 143546 124076 200631
rect 131948 200602 132000 200608
rect 177856 200660 177908 200666
rect 177856 200602 177908 200608
rect 180064 200660 180116 200666
rect 180064 200602 180116 200608
rect 124126 200560 124182 200569
rect 124126 200495 124182 200504
rect 123852 143540 123904 143546
rect 123852 143482 123904 143488
rect 124036 143540 124088 143546
rect 124036 143482 124088 143488
rect 123864 143342 123892 143482
rect 123760 143336 123812 143342
rect 123760 143278 123812 143284
rect 123852 143336 123904 143342
rect 123852 143278 123904 143284
rect 123772 142730 123800 143278
rect 123760 142724 123812 142730
rect 123760 142666 123812 142672
rect 124140 142154 124168 200495
rect 131960 200433 131988 200602
rect 132038 200560 132094 200569
rect 132038 200495 132094 200504
rect 132052 200462 132080 200495
rect 132040 200456 132092 200462
rect 126610 200424 126666 200433
rect 126610 200359 126666 200368
rect 131946 200424 132002 200433
rect 132040 200398 132092 200404
rect 131946 200359 132002 200368
rect 125600 200116 125652 200122
rect 125600 200058 125652 200064
rect 125232 199980 125284 199986
rect 125232 199922 125284 199928
rect 124864 194812 124916 194818
rect 124864 194754 124916 194760
rect 124496 148708 124548 148714
rect 124496 148650 124548 148656
rect 124048 142126 124168 142154
rect 124048 141001 124076 142126
rect 124034 140992 124090 141001
rect 124034 140927 124090 140936
rect 124048 139890 124076 140927
rect 124048 139862 124108 139890
rect 123556 139602 123892 139618
rect 123556 139596 123904 139602
rect 123556 139590 123852 139596
rect 123852 139538 123904 139544
rect 124508 139369 124536 148650
rect 124588 143540 124640 143546
rect 124588 143482 124640 143488
rect 124600 140826 124628 143482
rect 124876 143342 124904 194754
rect 125244 194070 125272 199922
rect 125612 198014 125640 200058
rect 126624 199481 126652 200359
rect 130936 200320 130988 200326
rect 128910 200288 128966 200297
rect 130936 200262 130988 200268
rect 128910 200223 128966 200232
rect 127532 199912 127584 199918
rect 127532 199854 127584 199860
rect 126610 199472 126666 199481
rect 126610 199407 126666 199416
rect 126336 198824 126388 198830
rect 126336 198766 126388 198772
rect 125600 198008 125652 198014
rect 125600 197950 125652 197956
rect 126152 197804 126204 197810
rect 126152 197746 126204 197752
rect 125232 194064 125284 194070
rect 125232 194006 125284 194012
rect 125508 188420 125560 188426
rect 125508 188362 125560 188368
rect 125048 148912 125100 148918
rect 125048 148854 125100 148860
rect 124864 143336 124916 143342
rect 124864 143278 124916 143284
rect 124588 140820 124640 140826
rect 124588 140762 124640 140768
rect 124956 140820 125008 140826
rect 124956 140762 125008 140768
rect 124968 139890 124996 140762
rect 125060 139913 125088 148854
rect 125230 148608 125286 148617
rect 125230 148543 125286 148552
rect 125244 140321 125272 148543
rect 125416 141296 125468 141302
rect 125416 141238 125468 141244
rect 125428 140865 125456 141238
rect 125414 140856 125470 140865
rect 125414 140791 125470 140800
rect 125230 140312 125286 140321
rect 125230 140247 125286 140256
rect 124660 139862 124996 139890
rect 125046 139904 125102 139913
rect 125428 139890 125456 140791
rect 125212 139862 125456 139890
rect 125046 139839 125102 139848
rect 125520 139369 125548 188362
rect 125598 141672 125654 141681
rect 125598 141607 125654 141616
rect 125612 139754 125640 141607
rect 125968 140752 126020 140758
rect 125968 140694 126020 140700
rect 125612 139738 125916 139754
rect 125612 139732 125928 139738
rect 125612 139726 125876 139732
rect 125876 139674 125928 139680
rect 125980 139369 126008 140694
rect 126164 139369 126192 197746
rect 126244 187468 126296 187474
rect 126244 187410 126296 187416
rect 126256 140622 126284 187410
rect 126348 140690 126376 198766
rect 126704 198620 126756 198626
rect 126704 198562 126756 198568
rect 126428 189508 126480 189514
rect 126428 189450 126480 189456
rect 126336 140684 126388 140690
rect 126336 140626 126388 140632
rect 126244 140616 126296 140622
rect 126244 140558 126296 140564
rect 126440 140554 126468 189450
rect 126612 149048 126664 149054
rect 126612 148990 126664 148996
rect 126520 148164 126572 148170
rect 126520 148106 126572 148112
rect 126532 141370 126560 148106
rect 126520 141364 126572 141370
rect 126520 141306 126572 141312
rect 126624 140758 126652 148990
rect 126612 140752 126664 140758
rect 126612 140694 126664 140700
rect 126428 140548 126480 140554
rect 126428 140490 126480 140496
rect 126716 140321 126744 198562
rect 127544 198286 127572 199854
rect 128820 199708 128872 199714
rect 128820 199650 128872 199656
rect 128832 199617 128860 199650
rect 128818 199608 128874 199617
rect 128818 199543 128874 199552
rect 127532 198280 127584 198286
rect 127532 198222 127584 198228
rect 127624 182028 127676 182034
rect 127624 181970 127676 181976
rect 126980 147280 127032 147286
rect 126980 147222 127032 147228
rect 126992 146441 127020 147222
rect 126978 146432 127034 146441
rect 126978 146367 127034 146376
rect 126794 143440 126850 143449
rect 126794 143375 126850 143384
rect 126808 142225 126836 143375
rect 126794 142216 126850 142225
rect 126794 142151 126850 142160
rect 126702 140312 126758 140321
rect 126702 140247 126758 140256
rect 126808 140162 126836 142151
rect 126888 142044 126940 142050
rect 126888 141986 126940 141992
rect 126900 140894 126928 141986
rect 126888 140888 126940 140894
rect 126888 140830 126940 140836
rect 126716 140134 126836 140162
rect 126716 139754 126744 140134
rect 126900 140026 126928 140830
rect 126992 140758 127020 146367
rect 127348 141976 127400 141982
rect 127348 141918 127400 141924
rect 127360 141137 127388 141918
rect 127346 141128 127402 141137
rect 127346 141063 127402 141072
rect 126980 140752 127032 140758
rect 126980 140694 127032 140700
rect 126316 139726 126744 139754
rect 126808 139998 126928 140026
rect 126808 139754 126836 139998
rect 127360 139890 127388 141063
rect 127360 139862 127420 139890
rect 126808 139726 126868 139754
rect 127636 139369 127664 181970
rect 128452 142792 128504 142798
rect 128452 142734 128504 142740
rect 127716 140752 127768 140758
rect 127716 140694 127768 140700
rect 127728 139890 127756 140694
rect 127728 139862 127972 139890
rect 128464 139754 128492 142734
rect 128924 140185 128952 200223
rect 130198 200152 130254 200161
rect 130198 200087 130254 200096
rect 129646 199064 129702 199073
rect 129646 198999 129702 199008
rect 129186 197296 129242 197305
rect 129186 197231 129242 197240
rect 129096 183116 129148 183122
rect 129096 183058 129148 183064
rect 129108 142730 129136 183058
rect 129096 142724 129148 142730
rect 129096 142666 129148 142672
rect 128910 140176 128966 140185
rect 128910 140111 128966 140120
rect 129200 140049 129228 197231
rect 129280 180328 129332 180334
rect 129280 180270 129332 180276
rect 129292 140078 129320 180270
rect 129372 144220 129424 144226
rect 129372 144162 129424 144168
rect 129384 142798 129412 144162
rect 129556 143200 129608 143206
rect 129556 143142 129608 143148
rect 129372 142792 129424 142798
rect 129372 142734 129424 142740
rect 129280 140072 129332 140078
rect 129186 140040 129242 140049
rect 129280 140014 129332 140020
rect 129186 139975 129242 139984
rect 129384 139890 129412 142734
rect 129568 141098 129596 143142
rect 129556 141092 129608 141098
rect 129556 141034 129608 141040
rect 129076 139862 129412 139890
rect 129568 139890 129596 141034
rect 129660 140162 129688 198999
rect 130212 198937 130240 200087
rect 130198 198928 130254 198937
rect 130198 198863 130254 198872
rect 130948 198694 130976 200262
rect 131578 200152 131634 200161
rect 131578 200087 131634 200096
rect 132052 200110 132388 200138
rect 131592 199646 131620 200087
rect 131946 200016 132002 200025
rect 131946 199951 132002 199960
rect 131580 199640 131632 199646
rect 131580 199582 131632 199588
rect 131488 199232 131540 199238
rect 131488 199174 131540 199180
rect 131580 199232 131632 199238
rect 131580 199174 131632 199180
rect 131500 198801 131528 199174
rect 131486 198792 131542 198801
rect 131486 198727 131542 198736
rect 130936 198688 130988 198694
rect 130936 198630 130988 198636
rect 131028 197668 131080 197674
rect 131028 197610 131080 197616
rect 130568 197328 130620 197334
rect 130568 197270 130620 197276
rect 130474 197160 130530 197169
rect 130474 197095 130530 197104
rect 130384 188352 130436 188358
rect 130384 188294 130436 188300
rect 130290 146296 130346 146305
rect 130290 146231 130346 146240
rect 129830 146160 129886 146169
rect 129830 146095 129886 146104
rect 129740 145444 129792 145450
rect 129740 145386 129792 145392
rect 129752 142254 129780 145386
rect 129844 143206 129872 146095
rect 129922 146024 129978 146033
rect 129922 145959 129978 145968
rect 129832 143200 129884 143206
rect 129832 143142 129884 143148
rect 129936 142322 129964 145959
rect 130016 144764 130068 144770
rect 130016 144706 130068 144712
rect 130028 144226 130056 144706
rect 130016 144220 130068 144226
rect 130016 144162 130068 144168
rect 129924 142316 129976 142322
rect 129924 142258 129976 142264
rect 129740 142248 129792 142254
rect 129740 142190 129792 142196
rect 130028 142154 130056 144162
rect 130028 142126 130148 142154
rect 129660 140134 129780 140162
rect 129752 140078 129780 140134
rect 129740 140072 129792 140078
rect 129740 140014 129792 140020
rect 130016 140004 130068 140010
rect 130016 139946 130068 139952
rect 129568 139862 129628 139890
rect 128820 139800 128872 139806
rect 128464 139748 128820 139754
rect 128464 139742 128872 139748
rect 128464 139726 128860 139742
rect 130028 139369 130056 139946
rect 130120 139890 130148 142126
rect 130304 139890 130332 146231
rect 130396 141914 130424 188294
rect 130384 141908 130436 141914
rect 130384 141850 130436 141856
rect 130488 140010 130516 197095
rect 130580 145518 130608 197270
rect 130568 145512 130620 145518
rect 130568 145454 130620 145460
rect 130476 140004 130528 140010
rect 130476 139946 130528 139952
rect 130120 139862 130180 139890
rect 130304 139862 130732 139890
rect 131040 139369 131068 197610
rect 131592 192846 131620 199174
rect 131960 198734 131988 199951
rect 131868 198706 131988 198734
rect 131580 192840 131632 192846
rect 131580 192782 131632 192788
rect 131868 190454 131896 198706
rect 132052 195265 132080 200110
rect 132466 199968 132494 200124
rect 132328 199940 132494 199968
rect 132224 197872 132276 197878
rect 132224 197814 132276 197820
rect 132038 195256 132094 195265
rect 132038 195191 132094 195200
rect 131868 190426 131988 190454
rect 131764 188488 131816 188494
rect 131764 188430 131816 188436
rect 131304 146260 131356 146266
rect 131304 146202 131356 146208
rect 131212 146192 131264 146198
rect 131212 146134 131264 146140
rect 131118 145888 131174 145897
rect 131118 145823 131174 145832
rect 131132 143478 131160 145823
rect 131120 143472 131172 143478
rect 131120 143414 131172 143420
rect 131224 143342 131252 146134
rect 131212 143336 131264 143342
rect 131212 143278 131264 143284
rect 131212 142724 131264 142730
rect 131212 142666 131264 142672
rect 131224 139890 131252 142666
rect 131316 140758 131344 146202
rect 131396 144288 131448 144294
rect 131396 144230 131448 144236
rect 131408 142730 131436 144230
rect 131488 143540 131540 143546
rect 131488 143482 131540 143488
rect 131580 143540 131632 143546
rect 131580 143482 131632 143488
rect 131396 142724 131448 142730
rect 131396 142666 131448 142672
rect 131304 140752 131356 140758
rect 131304 140694 131356 140700
rect 131500 139890 131528 143482
rect 131592 142798 131620 143482
rect 131580 142792 131632 142798
rect 131580 142734 131632 142740
rect 131776 141846 131804 188430
rect 131960 176654 131988 190426
rect 131868 176626 131988 176654
rect 131868 148782 131896 176626
rect 131856 148776 131908 148782
rect 131856 148718 131908 148724
rect 131764 141840 131816 141846
rect 131764 141782 131816 141788
rect 131224 139862 131284 139890
rect 131500 139862 131836 139890
rect 132236 139369 132264 197814
rect 132328 188465 132356 199940
rect 132558 199866 132586 200124
rect 132512 199838 132586 199866
rect 132512 198422 132540 199838
rect 132650 199764 132678 200124
rect 132604 199736 132678 199764
rect 132742 199764 132770 200124
rect 132834 199889 132862 200124
rect 132926 199918 132954 200124
rect 132914 199912 132966 199918
rect 132820 199880 132876 199889
rect 132914 199854 132966 199860
rect 132820 199815 132876 199824
rect 132868 199776 132920 199782
rect 132742 199736 132816 199764
rect 132500 198416 132552 198422
rect 132500 198358 132552 198364
rect 132604 194478 132632 199736
rect 132788 197441 132816 199736
rect 133018 199764 133046 200124
rect 133110 199918 133138 200124
rect 133202 199918 133230 200124
rect 133098 199912 133150 199918
rect 133098 199854 133150 199860
rect 133190 199912 133242 199918
rect 133190 199854 133242 199860
rect 133294 199850 133322 200124
rect 133386 199889 133414 200124
rect 133478 199918 133506 200124
rect 133466 199912 133518 199918
rect 133372 199880 133428 199889
rect 133282 199844 133334 199850
rect 133466 199854 133518 199860
rect 133372 199815 133428 199824
rect 133282 199786 133334 199792
rect 133018 199736 133092 199764
rect 132868 199718 132920 199724
rect 132774 197432 132830 197441
rect 132774 197367 132830 197376
rect 132776 196988 132828 196994
rect 132776 196930 132828 196936
rect 132788 196314 132816 196930
rect 132776 196308 132828 196314
rect 132776 196250 132828 196256
rect 132592 194472 132644 194478
rect 132592 194414 132644 194420
rect 132880 191834 132908 199718
rect 132960 197192 133012 197198
rect 132960 197134 133012 197140
rect 132972 196858 133000 197134
rect 132960 196852 133012 196858
rect 132960 196794 133012 196800
rect 133064 194177 133092 199736
rect 133328 199708 133380 199714
rect 133328 199650 133380 199656
rect 133420 199708 133472 199714
rect 133570 199696 133598 200124
rect 133662 199764 133690 200124
rect 133754 199918 133782 200124
rect 133742 199912 133794 199918
rect 133742 199854 133794 199860
rect 133662 199736 133736 199764
rect 133570 199668 133644 199696
rect 133420 199650 133472 199656
rect 133144 199640 133196 199646
rect 133144 199582 133196 199588
rect 133156 199345 133184 199582
rect 133142 199336 133198 199345
rect 133142 199271 133198 199280
rect 133142 199064 133198 199073
rect 133142 198999 133144 199008
rect 133196 198999 133198 199008
rect 133144 198970 133196 198976
rect 133340 198558 133368 199650
rect 133328 198552 133380 198558
rect 133328 198494 133380 198500
rect 133144 196988 133196 196994
rect 133144 196930 133196 196936
rect 133156 196722 133184 196930
rect 133144 196716 133196 196722
rect 133144 196658 133196 196664
rect 133328 196512 133380 196518
rect 133328 196454 133380 196460
rect 133340 196314 133368 196454
rect 133328 196308 133380 196314
rect 133328 196250 133380 196256
rect 133050 194168 133106 194177
rect 133050 194103 133106 194112
rect 132880 191806 133092 191834
rect 132868 188964 132920 188970
rect 132868 188906 132920 188912
rect 132314 188456 132370 188465
rect 132314 188391 132370 188400
rect 132684 187536 132736 187542
rect 132684 187478 132736 187484
rect 132696 151230 132724 187478
rect 132684 151224 132736 151230
rect 132684 151166 132736 151172
rect 132592 143064 132644 143070
rect 132592 143006 132644 143012
rect 132316 140752 132368 140758
rect 132316 140694 132368 140700
rect 132328 139890 132356 140694
rect 132604 139890 132632 143006
rect 132880 141778 132908 188906
rect 133064 148345 133092 191806
rect 133432 188970 133460 199650
rect 133616 198529 133644 199668
rect 133602 198520 133658 198529
rect 133602 198455 133658 198464
rect 133708 198200 133736 199736
rect 133846 199696 133874 200124
rect 133938 199764 133966 200124
rect 134030 199918 134058 200124
rect 134122 199918 134150 200124
rect 134018 199912 134070 199918
rect 134018 199854 134070 199860
rect 134110 199912 134162 199918
rect 134110 199854 134162 199860
rect 133938 199736 134012 199764
rect 133846 199668 133920 199696
rect 133616 198172 133736 198200
rect 133616 198082 133644 198172
rect 133604 198076 133656 198082
rect 133604 198018 133656 198024
rect 133696 196036 133748 196042
rect 133696 195978 133748 195984
rect 133708 195906 133736 195978
rect 133696 195900 133748 195906
rect 133696 195842 133748 195848
rect 133420 188964 133472 188970
rect 133420 188906 133472 188912
rect 133892 187542 133920 199668
rect 133984 189145 134012 199736
rect 134064 199640 134116 199646
rect 134214 199628 134242 200124
rect 134306 199889 134334 200124
rect 134292 199880 134348 199889
rect 134292 199815 134348 199824
rect 134398 199764 134426 200124
rect 134490 199918 134518 200124
rect 134582 199918 134610 200124
rect 134674 199918 134702 200124
rect 134478 199912 134530 199918
rect 134478 199854 134530 199860
rect 134570 199912 134622 199918
rect 134570 199854 134622 199860
rect 134662 199912 134714 199918
rect 134662 199854 134714 199860
rect 134352 199736 134426 199764
rect 134524 199776 134576 199782
rect 134214 199600 134288 199628
rect 134064 199582 134116 199588
rect 134076 194002 134104 199582
rect 134156 196104 134208 196110
rect 134156 196046 134208 196052
rect 134064 193996 134116 194002
rect 134064 193938 134116 193944
rect 134168 191298 134196 196046
rect 134076 191270 134196 191298
rect 134076 190126 134104 191270
rect 134260 191162 134288 199600
rect 134352 195770 134380 199736
rect 134524 199718 134576 199724
rect 134616 199776 134668 199782
rect 134766 199764 134794 200124
rect 134858 199889 134886 200124
rect 134844 199880 134900 199889
rect 134844 199815 134900 199824
rect 134950 199764 134978 200124
rect 134766 199736 134840 199764
rect 134616 199718 134668 199724
rect 134340 195764 134392 195770
rect 134340 195706 134392 195712
rect 134168 191134 134288 191162
rect 134064 190120 134116 190126
rect 134064 190062 134116 190068
rect 134168 189718 134196 191134
rect 134536 189802 134564 199718
rect 134628 196897 134656 199718
rect 134708 199640 134760 199646
rect 134708 199582 134760 199588
rect 134614 196888 134670 196897
rect 134614 196823 134670 196832
rect 134720 196110 134748 199582
rect 134708 196104 134760 196110
rect 134708 196046 134760 196052
rect 134812 190058 134840 199736
rect 134904 199736 134978 199764
rect 134904 198150 134932 199736
rect 135042 199696 135070 200124
rect 135134 199764 135162 200124
rect 135226 199918 135254 200124
rect 135214 199912 135266 199918
rect 135214 199854 135266 199860
rect 135318 199764 135346 200124
rect 135134 199736 135208 199764
rect 134996 199668 135070 199696
rect 134892 198144 134944 198150
rect 134892 198086 134944 198092
rect 134800 190052 134852 190058
rect 134800 189994 134852 190000
rect 134996 189922 135024 199668
rect 135180 197441 135208 199736
rect 135272 199736 135346 199764
rect 135410 199764 135438 200124
rect 135502 199918 135530 200124
rect 135490 199912 135542 199918
rect 135594 199889 135622 200124
rect 135686 199918 135714 200124
rect 135674 199912 135726 199918
rect 135490 199854 135542 199860
rect 135580 199880 135636 199889
rect 135674 199854 135726 199860
rect 135580 199815 135636 199824
rect 135536 199776 135588 199782
rect 135410 199736 135484 199764
rect 135166 197432 135222 197441
rect 135166 197367 135222 197376
rect 134984 189916 135036 189922
rect 134984 189858 135036 189864
rect 134260 189774 134564 189802
rect 135272 189786 135300 199736
rect 135352 199640 135404 199646
rect 135352 199582 135404 199588
rect 135364 199481 135392 199582
rect 135350 199472 135406 199481
rect 135350 199407 135406 199416
rect 135260 189780 135312 189786
rect 134156 189712 134208 189718
rect 134156 189654 134208 189660
rect 133970 189136 134026 189145
rect 133970 189071 134026 189080
rect 133880 187536 133932 187542
rect 133880 187478 133932 187484
rect 134260 151162 134288 189774
rect 135260 189722 135312 189728
rect 134432 189712 134484 189718
rect 134432 189654 134484 189660
rect 134248 151156 134300 151162
rect 134248 151098 134300 151104
rect 134444 151094 134472 189654
rect 135456 187105 135484 199736
rect 135778 199764 135806 200124
rect 135536 199718 135588 199724
rect 135732 199736 135806 199764
rect 135548 193934 135576 199718
rect 135628 199708 135680 199714
rect 135628 199650 135680 199656
rect 135536 193928 135588 193934
rect 135536 193870 135588 193876
rect 135640 188465 135668 199650
rect 135732 194206 135760 199736
rect 135870 199594 135898 200124
rect 135962 199730 135990 200124
rect 136054 199918 136082 200124
rect 136042 199912 136094 199918
rect 136042 199854 136094 199860
rect 136146 199764 136174 200124
rect 136238 199889 136266 200124
rect 136330 199918 136358 200124
rect 136318 199912 136370 199918
rect 136224 199880 136280 199889
rect 136318 199854 136370 199860
rect 136224 199815 136280 199824
rect 136422 199764 136450 200124
rect 136514 199918 136542 200124
rect 136502 199912 136554 199918
rect 136502 199854 136554 199860
rect 136100 199736 136174 199764
rect 136376 199736 136450 199764
rect 136606 199764 136634 200124
rect 136698 199918 136726 200124
rect 136790 199923 136818 200124
rect 136686 199912 136738 199918
rect 136686 199854 136738 199860
rect 136776 199914 136832 199923
rect 136882 199918 136910 200124
rect 136776 199849 136832 199858
rect 136870 199912 136922 199918
rect 136870 199854 136922 199860
rect 136732 199776 136784 199782
rect 136606 199736 136680 199764
rect 135962 199702 136036 199730
rect 135870 199566 135944 199594
rect 135720 194200 135772 194206
rect 135720 194142 135772 194148
rect 135916 189854 135944 199566
rect 136008 196217 136036 199702
rect 135994 196208 136050 196217
rect 135994 196143 136050 196152
rect 135996 196036 136048 196042
rect 135996 195978 136048 195984
rect 136008 195770 136036 195978
rect 135996 195764 136048 195770
rect 135996 195706 136048 195712
rect 136100 194138 136128 199736
rect 136180 199640 136232 199646
rect 136180 199582 136232 199588
rect 136192 198937 136220 199582
rect 136178 198928 136234 198937
rect 136178 198863 136234 198872
rect 136178 196344 136234 196353
rect 136178 196279 136234 196288
rect 136088 194132 136140 194138
rect 136088 194074 136140 194080
rect 136192 189990 136220 196279
rect 136270 196072 136326 196081
rect 136270 196007 136326 196016
rect 136180 189984 136232 189990
rect 136180 189926 136232 189932
rect 135904 189848 135956 189854
rect 135904 189790 135956 189796
rect 135626 188456 135682 188465
rect 135626 188391 135682 188400
rect 136284 188290 136312 196007
rect 136376 194274 136404 199736
rect 136456 199640 136508 199646
rect 136456 199582 136508 199588
rect 136548 199640 136600 199646
rect 136548 199582 136600 199588
rect 136468 194993 136496 199582
rect 136560 199481 136588 199582
rect 136546 199472 136602 199481
rect 136546 199407 136602 199416
rect 136652 199209 136680 199736
rect 136732 199718 136784 199724
rect 136824 199776 136876 199782
rect 136974 199764 137002 200124
rect 137066 199918 137094 200124
rect 137054 199912 137106 199918
rect 137158 199889 137186 200124
rect 137054 199854 137106 199860
rect 137144 199880 137200 199889
rect 137250 199850 137278 200124
rect 137144 199815 137200 199824
rect 137238 199844 137290 199850
rect 137238 199786 137290 199792
rect 137342 199764 137370 200124
rect 137434 199918 137462 200124
rect 137422 199912 137474 199918
rect 137526 199889 137554 200124
rect 137422 199854 137474 199860
rect 137512 199880 137568 199889
rect 137512 199815 137568 199824
rect 137618 199764 137646 200124
rect 136974 199736 137048 199764
rect 137342 199736 137508 199764
rect 136824 199718 136876 199724
rect 136638 199200 136694 199209
rect 136638 199135 136694 199144
rect 136548 198280 136600 198286
rect 136548 198222 136600 198228
rect 136454 194984 136510 194993
rect 136454 194919 136510 194928
rect 136364 194268 136416 194274
rect 136364 194210 136416 194216
rect 136560 192710 136588 198222
rect 136548 192704 136600 192710
rect 136548 192646 136600 192652
rect 136744 192545 136772 199718
rect 136836 199238 136864 199718
rect 136824 199232 136876 199238
rect 136824 199174 136876 199180
rect 136914 199200 136970 199209
rect 136914 199135 136970 199144
rect 136822 198928 136878 198937
rect 136822 198863 136878 198872
rect 136836 192574 136864 198863
rect 136928 194342 136956 199135
rect 136916 194336 136968 194342
rect 136916 194278 136968 194284
rect 137020 193186 137048 199736
rect 137100 199708 137152 199714
rect 137100 199650 137152 199656
rect 137192 199708 137244 199714
rect 137192 199650 137244 199656
rect 137008 193180 137060 193186
rect 137008 193122 137060 193128
rect 136824 192568 136876 192574
rect 136730 192536 136786 192545
rect 136824 192510 136876 192516
rect 136730 192471 136786 192480
rect 137112 190454 137140 199650
rect 137204 195106 137232 199650
rect 137374 199472 137430 199481
rect 137374 199407 137430 199416
rect 137204 195078 137324 195106
rect 137190 194984 137246 194993
rect 137190 194919 137246 194928
rect 137020 190426 137140 190454
rect 137020 188465 137048 190426
rect 137006 188456 137062 188465
rect 137006 188391 137062 188400
rect 135628 188284 135680 188290
rect 135628 188226 135680 188232
rect 136272 188284 136324 188290
rect 136272 188226 136324 188232
rect 135442 187096 135498 187105
rect 135442 187031 135498 187040
rect 134432 151088 134484 151094
rect 134432 151030 134484 151036
rect 135640 148646 135668 188226
rect 137204 187649 137232 194919
rect 137296 192681 137324 195078
rect 137282 192672 137338 192681
rect 137282 192607 137338 192616
rect 137282 188048 137338 188057
rect 137282 187983 137338 187992
rect 137190 187640 137246 187649
rect 137190 187575 137246 187584
rect 135628 148640 135680 148646
rect 135628 148582 135680 148588
rect 133050 148336 133106 148345
rect 133050 148271 133106 148280
rect 137296 147218 137324 187983
rect 137388 183122 137416 199407
rect 137480 186289 137508 199736
rect 137572 199736 137646 199764
rect 137572 190454 137600 199736
rect 137710 199696 137738 200124
rect 137802 199918 137830 200124
rect 137894 199923 137922 200124
rect 137790 199912 137842 199918
rect 137790 199854 137842 199860
rect 137880 199914 137936 199923
rect 137880 199849 137936 199858
rect 137836 199776 137888 199782
rect 137986 199764 138014 200124
rect 137836 199718 137888 199724
rect 137940 199736 138014 199764
rect 137664 199668 137738 199696
rect 137664 194818 137692 199668
rect 137848 199424 137876 199718
rect 137756 199396 137876 199424
rect 137652 194812 137704 194818
rect 137652 194754 137704 194760
rect 137756 192438 137784 199396
rect 137940 199356 137968 199736
rect 138078 199696 138106 200124
rect 138170 199889 138198 200124
rect 138262 199918 138290 200124
rect 138354 199918 138382 200124
rect 138250 199912 138302 199918
rect 138156 199880 138212 199889
rect 138250 199854 138302 199860
rect 138342 199912 138394 199918
rect 138342 199854 138394 199860
rect 138156 199815 138212 199824
rect 138204 199776 138256 199782
rect 138446 199764 138474 200124
rect 138538 199918 138566 200124
rect 138526 199912 138578 199918
rect 138526 199854 138578 199860
rect 138630 199764 138658 200124
rect 138256 199736 138336 199764
rect 138204 199718 138256 199724
rect 137848 199328 137968 199356
rect 138032 199668 138106 199696
rect 137848 197033 137876 199328
rect 137926 199064 137982 199073
rect 137926 198999 137982 199008
rect 137834 197024 137890 197033
rect 137834 196959 137890 196968
rect 137940 195702 137968 198999
rect 138032 198286 138060 199668
rect 138204 199640 138256 199646
rect 138124 199600 138204 199628
rect 138020 198280 138072 198286
rect 138020 198222 138072 198228
rect 138124 198132 138152 199600
rect 138204 199582 138256 199588
rect 138202 199472 138258 199481
rect 138202 199407 138258 199416
rect 138032 198104 138152 198132
rect 138032 195945 138060 198104
rect 138216 198064 138244 199407
rect 138124 198036 138244 198064
rect 138018 195936 138074 195945
rect 138018 195871 138074 195880
rect 137928 195696 137980 195702
rect 137928 195638 137980 195644
rect 137744 192432 137796 192438
rect 137744 192374 137796 192380
rect 137572 190426 137692 190454
rect 137664 188465 137692 190426
rect 137650 188456 137706 188465
rect 137650 188391 137706 188400
rect 137466 186280 137522 186289
rect 137466 186215 137522 186224
rect 137376 183116 137428 183122
rect 137376 183058 137428 183064
rect 138124 176654 138152 198036
rect 138308 197962 138336 199736
rect 138216 197934 138336 197962
rect 138400 199736 138474 199764
rect 138584 199736 138658 199764
rect 138722 199764 138750 200124
rect 138814 199918 138842 200124
rect 138802 199912 138854 199918
rect 138802 199854 138854 199860
rect 138722 199736 138796 199764
rect 138216 196625 138244 197934
rect 138296 197872 138348 197878
rect 138296 197814 138348 197820
rect 138308 197674 138336 197814
rect 138296 197668 138348 197674
rect 138296 197610 138348 197616
rect 138202 196616 138258 196625
rect 138202 196551 138258 196560
rect 138400 194993 138428 199736
rect 138480 199640 138532 199646
rect 138480 199582 138532 199588
rect 138492 196761 138520 199582
rect 138478 196752 138534 196761
rect 138478 196687 138534 196696
rect 138386 194984 138442 194993
rect 138386 194919 138442 194928
rect 138584 194857 138612 199736
rect 138664 199640 138716 199646
rect 138664 199582 138716 199588
rect 138676 198801 138704 199582
rect 138662 198792 138718 198801
rect 138662 198727 138718 198736
rect 138664 195424 138716 195430
rect 138664 195366 138716 195372
rect 138570 194848 138626 194857
rect 138570 194783 138626 194792
rect 138676 190398 138704 195366
rect 138768 194342 138796 199736
rect 138906 199730 138934 200124
rect 138998 199764 139026 200124
rect 139090 199918 139118 200124
rect 139182 199918 139210 200124
rect 139274 199918 139302 200124
rect 139366 199918 139394 200124
rect 139078 199912 139130 199918
rect 139078 199854 139130 199860
rect 139170 199912 139222 199918
rect 139170 199854 139222 199860
rect 139262 199912 139314 199918
rect 139262 199854 139314 199860
rect 139354 199912 139406 199918
rect 139354 199854 139406 199860
rect 139124 199776 139176 199782
rect 138998 199736 139072 199764
rect 138860 199702 138934 199730
rect 138860 199481 138888 199702
rect 138940 199640 138992 199646
rect 138940 199582 138992 199588
rect 138846 199472 138902 199481
rect 138846 199407 138902 199416
rect 138848 199232 138900 199238
rect 138848 199174 138900 199180
rect 138756 194336 138808 194342
rect 138756 194278 138808 194284
rect 138664 190392 138716 190398
rect 138664 190334 138716 190340
rect 138860 188465 138888 199174
rect 138952 197402 138980 199582
rect 139044 199238 139072 199736
rect 139124 199718 139176 199724
rect 139032 199232 139084 199238
rect 139032 199174 139084 199180
rect 138940 197396 138992 197402
rect 138940 197338 138992 197344
rect 139136 194993 139164 199718
rect 139216 199708 139268 199714
rect 139458 199696 139486 200124
rect 139216 199650 139268 199656
rect 139412 199668 139486 199696
rect 139228 199073 139256 199650
rect 139308 199640 139360 199646
rect 139308 199582 139360 199588
rect 139320 199345 139348 199582
rect 139306 199336 139362 199345
rect 139306 199271 139362 199280
rect 139214 199064 139270 199073
rect 139214 198999 139270 199008
rect 139214 198384 139270 198393
rect 139214 198319 139270 198328
rect 139228 197713 139256 198319
rect 139214 197704 139270 197713
rect 139214 197639 139270 197648
rect 139214 196072 139270 196081
rect 139214 196007 139270 196016
rect 139122 194984 139178 194993
rect 139122 194919 139178 194928
rect 138940 194336 138992 194342
rect 138940 194278 138992 194284
rect 138952 188601 138980 194278
rect 139228 190454 139256 196007
rect 139228 190426 139348 190454
rect 138938 188592 138994 188601
rect 138938 188527 138994 188536
rect 138846 188456 138902 188465
rect 138846 188391 138902 188400
rect 139320 188358 139348 190426
rect 139412 188494 139440 199668
rect 139550 199628 139578 200124
rect 139504 199600 139578 199628
rect 139400 188488 139452 188494
rect 139400 188430 139452 188436
rect 139308 188352 139360 188358
rect 139308 188294 139360 188300
rect 139504 176654 139532 199600
rect 139642 199560 139670 200124
rect 139734 199696 139762 200124
rect 139826 199764 139854 200124
rect 139918 199918 139946 200124
rect 139906 199912 139958 199918
rect 139906 199854 139958 199860
rect 140010 199764 140038 200124
rect 140102 199918 140130 200124
rect 140090 199912 140142 199918
rect 140090 199854 140142 199860
rect 140194 199764 140222 200124
rect 140286 199918 140314 200124
rect 140274 199912 140326 199918
rect 140274 199854 140326 199860
rect 140378 199850 140406 200124
rect 140470 199918 140498 200124
rect 140458 199912 140510 199918
rect 140458 199854 140510 199860
rect 140366 199844 140418 199850
rect 140366 199786 140418 199792
rect 139826 199736 139900 199764
rect 140010 199736 140084 199764
rect 139734 199668 139808 199696
rect 139596 199532 139670 199560
rect 139596 196654 139624 199532
rect 139780 199492 139808 199668
rect 139688 199464 139808 199492
rect 139688 199209 139716 199464
rect 139872 199424 139900 199736
rect 139952 199640 140004 199646
rect 139952 199582 140004 199588
rect 139780 199396 139900 199424
rect 139674 199200 139730 199209
rect 139674 199135 139730 199144
rect 139584 196648 139636 196654
rect 139584 196590 139636 196596
rect 139780 188601 139808 199396
rect 139964 199356 139992 199582
rect 139872 199328 139992 199356
rect 139872 195362 139900 199328
rect 140056 199288 140084 199736
rect 139964 199260 140084 199288
rect 140148 199736 140222 199764
rect 139860 195356 139912 195362
rect 139860 195298 139912 195304
rect 139964 190330 139992 199260
rect 140042 199064 140098 199073
rect 140042 198999 140098 199008
rect 140056 197441 140084 198999
rect 140042 197432 140098 197441
rect 140042 197367 140098 197376
rect 140044 197192 140096 197198
rect 140044 197134 140096 197140
rect 140056 196790 140084 197134
rect 140148 196858 140176 199736
rect 140562 199730 140590 200124
rect 140654 199850 140682 200124
rect 140746 199850 140774 200124
rect 140838 199918 140866 200124
rect 140930 199918 140958 200124
rect 141022 199918 141050 200124
rect 141114 199918 141142 200124
rect 141206 199918 141234 200124
rect 141298 199918 141326 200124
rect 141390 199918 141418 200124
rect 140826 199912 140878 199918
rect 140826 199854 140878 199860
rect 140918 199912 140970 199918
rect 140918 199854 140970 199860
rect 141010 199912 141062 199918
rect 141010 199854 141062 199860
rect 141102 199912 141154 199918
rect 141102 199854 141154 199860
rect 141194 199912 141246 199918
rect 141194 199854 141246 199860
rect 141286 199912 141338 199918
rect 141286 199854 141338 199860
rect 141378 199912 141430 199918
rect 141378 199854 141430 199860
rect 140642 199844 140694 199850
rect 140642 199786 140694 199792
rect 140734 199844 140786 199850
rect 140734 199786 140786 199792
rect 140320 199708 140372 199714
rect 140320 199650 140372 199656
rect 140412 199708 140464 199714
rect 140412 199650 140464 199656
rect 140516 199702 140590 199730
rect 140918 199776 140970 199782
rect 141482 199764 141510 200124
rect 141574 199918 141602 200124
rect 141666 199918 141694 200124
rect 141758 199918 141786 200124
rect 141850 199918 141878 200124
rect 141562 199912 141614 199918
rect 141562 199854 141614 199860
rect 141654 199912 141706 199918
rect 141654 199854 141706 199860
rect 141746 199912 141798 199918
rect 141746 199854 141798 199860
rect 141838 199912 141890 199918
rect 141838 199854 141890 199860
rect 141608 199776 141660 199782
rect 141482 199736 141556 199764
rect 140918 199718 140970 199724
rect 140228 199640 140280 199646
rect 140228 199582 140280 199588
rect 140240 199073 140268 199582
rect 140332 199345 140360 199650
rect 140318 199336 140374 199345
rect 140318 199271 140374 199280
rect 140318 199200 140374 199209
rect 140318 199135 140374 199144
rect 140226 199064 140282 199073
rect 140226 198999 140282 199008
rect 140226 198928 140282 198937
rect 140332 198898 140360 199135
rect 140226 198863 140282 198872
rect 140320 198892 140372 198898
rect 140136 196852 140188 196858
rect 140136 196794 140188 196800
rect 140044 196784 140096 196790
rect 140044 196726 140096 196732
rect 139952 190324 140004 190330
rect 139952 190266 140004 190272
rect 140240 190194 140268 198863
rect 140320 198834 140372 198840
rect 140228 190188 140280 190194
rect 140228 190130 140280 190136
rect 139766 188592 139822 188601
rect 139766 188527 139822 188536
rect 140424 188465 140452 199650
rect 140516 193866 140544 199702
rect 140596 199640 140648 199646
rect 140596 199582 140648 199588
rect 140688 199640 140740 199646
rect 140688 199582 140740 199588
rect 140780 199640 140832 199646
rect 140780 199582 140832 199588
rect 140608 199345 140636 199582
rect 140594 199336 140650 199345
rect 140594 199271 140650 199280
rect 140504 193860 140556 193866
rect 140504 193802 140556 193808
rect 140700 193118 140728 199582
rect 140792 195430 140820 199582
rect 140930 199356 140958 199718
rect 141102 199708 141154 199714
rect 141102 199650 141154 199656
rect 141240 199708 141292 199714
rect 141292 199668 141372 199696
rect 141240 199650 141292 199656
rect 141010 199640 141062 199646
rect 141010 199582 141062 199588
rect 141022 199424 141050 199582
rect 141114 199492 141142 199650
rect 141114 199464 141280 199492
rect 141022 199396 141188 199424
rect 140930 199328 141096 199356
rect 140780 195424 140832 195430
rect 140780 195366 140832 195372
rect 140688 193112 140740 193118
rect 140688 193054 140740 193060
rect 140410 188456 140466 188465
rect 140410 188391 140466 188400
rect 141068 182174 141096 199328
rect 141160 185502 141188 199396
rect 141252 190262 141280 199464
rect 141240 190256 141292 190262
rect 141240 190198 141292 190204
rect 141148 185496 141200 185502
rect 141148 185438 141200 185444
rect 140976 182146 141096 182174
rect 141344 182174 141372 199668
rect 141424 199640 141476 199646
rect 141424 199582 141476 199588
rect 141436 190602 141464 199582
rect 141424 190596 141476 190602
rect 141424 190538 141476 190544
rect 141344 182146 141464 182174
rect 138124 176626 138520 176654
rect 139504 176626 139808 176654
rect 137284 147212 137336 147218
rect 137284 147154 137336 147160
rect 138492 147082 138520 176626
rect 138480 147076 138532 147082
rect 138480 147018 138532 147024
rect 139780 146946 139808 176626
rect 140976 147150 141004 182146
rect 140964 147144 141016 147150
rect 140964 147086 141016 147092
rect 139768 146940 139820 146946
rect 139768 146882 139820 146888
rect 138112 144696 138164 144702
rect 138112 144638 138164 144644
rect 140870 144664 140926 144673
rect 137560 143472 137612 143478
rect 137560 143414 137612 143420
rect 133144 143404 133196 143410
rect 133144 143346 133196 143352
rect 132868 141772 132920 141778
rect 132868 141714 132920 141720
rect 133156 139890 133184 143346
rect 135444 143336 135496 143342
rect 135444 143278 135496 143284
rect 134800 143132 134852 143138
rect 134800 143074 134852 143080
rect 134248 142316 134300 142322
rect 134248 142258 134300 142264
rect 133880 142248 133932 142254
rect 133880 142190 133932 142196
rect 133892 139890 133920 142190
rect 134260 139890 134288 142258
rect 134812 139890 134840 143074
rect 135456 139890 135484 143278
rect 136640 143268 136692 143274
rect 136640 143210 136692 143216
rect 135904 143200 135956 143206
rect 135904 143142 135956 143148
rect 135916 139890 135944 143142
rect 136652 139890 136680 143210
rect 137008 141636 137060 141642
rect 137008 141578 137060 141584
rect 137020 139890 137048 141578
rect 137572 139890 137600 143414
rect 138124 139890 138152 144638
rect 140870 144599 140926 144608
rect 138662 143984 138718 143993
rect 138662 143919 138718 143928
rect 138676 139890 138704 143919
rect 139398 143848 139454 143857
rect 139398 143783 139454 143792
rect 139412 139890 139440 143783
rect 139768 142996 139820 143002
rect 139768 142938 139820 142944
rect 139780 139890 139808 142938
rect 140320 141704 140372 141710
rect 140320 141646 140372 141652
rect 140332 139890 140360 141646
rect 140884 139890 140912 144599
rect 141436 141545 141464 182146
rect 141528 176654 141556 199736
rect 141608 199718 141660 199724
rect 141700 199776 141752 199782
rect 141942 199764 141970 200124
rect 141700 199718 141752 199724
rect 141896 199736 141970 199764
rect 142034 199764 142062 200124
rect 142126 199923 142154 200124
rect 142112 199914 142168 199923
rect 142112 199849 142168 199858
rect 142218 199764 142246 200124
rect 142034 199736 142108 199764
rect 141620 182034 141648 199718
rect 141712 190369 141740 199718
rect 141792 199708 141844 199714
rect 141792 199650 141844 199656
rect 141804 194410 141832 199650
rect 141792 194404 141844 194410
rect 141792 194346 141844 194352
rect 141896 190466 141924 199736
rect 141976 199640 142028 199646
rect 141976 199582 142028 199588
rect 141988 192506 142016 199582
rect 141976 192500 142028 192506
rect 141976 192442 142028 192448
rect 142080 191185 142108 199736
rect 142172 199736 142246 199764
rect 142310 199764 142338 200124
rect 142402 199918 142430 200124
rect 142494 199923 142522 200124
rect 142390 199912 142442 199918
rect 142390 199854 142442 199860
rect 142480 199914 142536 199923
rect 142586 199918 142614 200124
rect 142678 199918 142706 200124
rect 142770 199918 142798 200124
rect 142480 199849 142536 199858
rect 142574 199912 142626 199918
rect 142574 199854 142626 199860
rect 142666 199912 142718 199918
rect 142666 199854 142718 199860
rect 142758 199912 142810 199918
rect 142758 199854 142810 199860
rect 142436 199776 142488 199782
rect 142310 199736 142384 199764
rect 142066 191176 142122 191185
rect 142066 191111 142122 191120
rect 142172 191049 142200 199736
rect 142252 199640 142304 199646
rect 142252 199582 142304 199588
rect 142264 192817 142292 199582
rect 142356 195401 142384 199736
rect 142436 199718 142488 199724
rect 142712 199776 142764 199782
rect 142862 199764 142890 200124
rect 142954 199918 142982 200124
rect 142942 199912 142994 199918
rect 142942 199854 142994 199860
rect 142712 199718 142764 199724
rect 142816 199736 142890 199764
rect 142448 199617 142476 199718
rect 142528 199708 142580 199714
rect 142528 199650 142580 199656
rect 142620 199708 142672 199714
rect 142620 199650 142672 199656
rect 142434 199608 142490 199617
rect 142434 199543 142490 199552
rect 142540 196994 142568 199650
rect 142528 196988 142580 196994
rect 142528 196930 142580 196936
rect 142632 195974 142660 199650
rect 142448 195946 142660 195974
rect 142448 195770 142476 195946
rect 142436 195764 142488 195770
rect 142436 195706 142488 195712
rect 142342 195392 142398 195401
rect 142342 195327 142398 195336
rect 142724 195276 142752 199718
rect 142816 196926 142844 199736
rect 143046 199730 143074 200124
rect 143000 199702 143074 199730
rect 142896 199640 142948 199646
rect 142896 199582 142948 199588
rect 142908 197198 142936 199582
rect 142896 197192 142948 197198
rect 142896 197134 142948 197140
rect 142804 196920 142856 196926
rect 142804 196862 142856 196868
rect 142540 195248 142752 195276
rect 142250 192808 142306 192817
rect 142250 192743 142306 192752
rect 142158 191040 142214 191049
rect 142158 190975 142214 190984
rect 141884 190460 141936 190466
rect 141884 190402 141936 190408
rect 141698 190360 141754 190369
rect 141698 190295 141754 190304
rect 142068 185496 142120 185502
rect 142068 185438 142120 185444
rect 141608 182028 141660 182034
rect 141608 181970 141660 181976
rect 142080 180849 142108 185438
rect 142066 180840 142122 180849
rect 142066 180775 142122 180784
rect 142066 180704 142122 180713
rect 142066 180639 142122 180648
rect 141528 176626 141648 176654
rect 141516 142928 141568 142934
rect 141516 142870 141568 142876
rect 141422 141536 141478 141545
rect 141422 141471 141478 141480
rect 141528 139890 141556 142870
rect 141620 141273 141648 176626
rect 142080 171193 142108 180639
rect 142066 171184 142122 171193
rect 142066 171119 142122 171128
rect 142066 171048 142122 171057
rect 142066 170983 142122 170992
rect 142080 161537 142108 170983
rect 142066 161528 142122 161537
rect 142066 161463 142122 161472
rect 142066 161392 142122 161401
rect 142066 161327 142122 161336
rect 142080 151881 142108 161327
rect 142066 151872 142122 151881
rect 142066 151807 142122 151816
rect 142066 151736 142122 151745
rect 142066 151671 142122 151680
rect 142080 142361 142108 151671
rect 142540 148238 142568 195248
rect 143000 195140 143028 199702
rect 143138 199594 143166 200124
rect 143230 199730 143258 200124
rect 143322 199918 143350 200124
rect 143414 199918 143442 200124
rect 143506 199923 143534 200124
rect 143310 199912 143362 199918
rect 143310 199854 143362 199860
rect 143402 199912 143454 199918
rect 143402 199854 143454 199860
rect 143492 199914 143548 199923
rect 143492 199849 143548 199858
rect 143598 199730 143626 200124
rect 143230 199702 143304 199730
rect 143092 199566 143166 199594
rect 143092 195634 143120 199566
rect 143276 197130 143304 199702
rect 143356 199708 143408 199714
rect 143356 199650 143408 199656
rect 143448 199708 143500 199714
rect 143448 199650 143500 199656
rect 143552 199702 143626 199730
rect 143264 197124 143316 197130
rect 143264 197066 143316 197072
rect 143080 195628 143132 195634
rect 143080 195570 143132 195576
rect 142632 195112 143028 195140
rect 142632 148986 142660 195112
rect 143368 176654 143396 199650
rect 143460 196450 143488 199650
rect 143448 196444 143500 196450
rect 143448 196386 143500 196392
rect 143552 188426 143580 199702
rect 143690 199696 143718 200124
rect 143782 199764 143810 200124
rect 143874 199918 143902 200124
rect 143966 199918 143994 200124
rect 143862 199912 143914 199918
rect 143862 199854 143914 199860
rect 143954 199912 144006 199918
rect 143954 199854 144006 199860
rect 143782 199736 143856 199764
rect 143690 199668 143764 199696
rect 143632 199572 143684 199578
rect 143632 199514 143684 199520
rect 143644 199170 143672 199514
rect 143632 199164 143684 199170
rect 143632 199106 143684 199112
rect 143736 198490 143764 199668
rect 143724 198484 143776 198490
rect 143724 198426 143776 198432
rect 143828 198370 143856 199736
rect 144058 199730 144086 200124
rect 144150 199923 144178 200124
rect 144136 199914 144192 199923
rect 144136 199849 144192 199858
rect 144242 199730 144270 200124
rect 144334 199923 144362 200124
rect 144320 199914 144376 199923
rect 144320 199849 144376 199858
rect 144426 199764 144454 200124
rect 144518 199923 144546 200124
rect 144504 199914 144560 199923
rect 144610 199918 144638 200124
rect 144702 199918 144730 200124
rect 144504 199849 144560 199858
rect 144598 199912 144650 199918
rect 144598 199854 144650 199860
rect 144690 199912 144742 199918
rect 144690 199854 144742 199860
rect 144644 199776 144696 199782
rect 144426 199736 144500 199764
rect 144058 199714 144132 199730
rect 144058 199708 144144 199714
rect 144058 199702 144092 199708
rect 144242 199702 144316 199730
rect 144092 199650 144144 199656
rect 143908 199640 143960 199646
rect 143908 199582 143960 199588
rect 144000 199640 144052 199646
rect 144000 199582 144052 199588
rect 144182 199608 144238 199617
rect 143736 198342 143856 198370
rect 143736 196790 143764 198342
rect 143724 196784 143776 196790
rect 143724 196726 143776 196732
rect 143920 195129 143948 199582
rect 143906 195120 143962 195129
rect 143906 195055 143962 195064
rect 144012 192914 144040 199582
rect 144092 199572 144144 199578
rect 144182 199543 144238 199552
rect 144092 199514 144144 199520
rect 144104 196518 144132 199514
rect 144196 197470 144224 199543
rect 144184 197464 144236 197470
rect 144184 197406 144236 197412
rect 144092 196512 144144 196518
rect 144092 196454 144144 196460
rect 144288 196058 144316 199702
rect 144368 199640 144420 199646
rect 144368 199582 144420 199588
rect 144380 198762 144408 199582
rect 144368 198756 144420 198762
rect 144368 198698 144420 198704
rect 144288 196030 144408 196058
rect 144380 192982 144408 196030
rect 144368 192976 144420 192982
rect 144368 192918 144420 192924
rect 144000 192908 144052 192914
rect 144000 192850 144052 192856
rect 143816 190596 143868 190602
rect 143816 190538 143868 190544
rect 143540 188420 143592 188426
rect 143540 188362 143592 188368
rect 143000 176626 143396 176654
rect 142620 148980 142672 148986
rect 142620 148922 142672 148928
rect 143000 148306 143028 176626
rect 142988 148300 143040 148306
rect 142988 148242 143040 148248
rect 142528 148232 142580 148238
rect 142528 148174 142580 148180
rect 143828 144634 143856 190538
rect 144472 188329 144500 199736
rect 144550 199744 144606 199753
rect 144794 199764 144822 200124
rect 144886 199889 144914 200124
rect 144978 199918 145006 200124
rect 144966 199912 145018 199918
rect 144872 199880 144928 199889
rect 144966 199854 145018 199860
rect 144872 199815 144928 199824
rect 144644 199718 144696 199724
rect 144748 199736 144822 199764
rect 144550 199679 144606 199688
rect 144564 192642 144592 199679
rect 144552 192636 144604 192642
rect 144552 192578 144604 192584
rect 144458 188320 144514 188329
rect 144458 188255 144514 188264
rect 144656 183841 144684 199718
rect 144748 193050 144776 199736
rect 145070 199730 145098 200124
rect 145162 199764 145190 200124
rect 145254 199918 145282 200124
rect 145346 199918 145374 200124
rect 145438 199918 145466 200124
rect 145530 199923 145558 200124
rect 145242 199912 145294 199918
rect 145242 199854 145294 199860
rect 145334 199912 145386 199918
rect 145334 199854 145386 199860
rect 145426 199912 145478 199918
rect 145426 199854 145478 199860
rect 145516 199914 145572 199923
rect 145622 199918 145650 200124
rect 145516 199849 145572 199858
rect 145610 199912 145662 199918
rect 145610 199854 145662 199860
rect 145380 199776 145432 199782
rect 145162 199736 145236 199764
rect 144920 199708 144972 199714
rect 144920 199650 144972 199656
rect 145024 199702 145098 199730
rect 144828 199572 144880 199578
rect 144828 199514 144880 199520
rect 144840 198694 144868 199514
rect 144828 198688 144880 198694
rect 144828 198630 144880 198636
rect 144932 198064 144960 199650
rect 144840 198036 144960 198064
rect 144840 197810 144868 198036
rect 144828 197804 144880 197810
rect 144828 197746 144880 197752
rect 145024 195838 145052 199702
rect 145104 199572 145156 199578
rect 145104 199514 145156 199520
rect 145012 195832 145064 195838
rect 145012 195774 145064 195780
rect 145116 195294 145144 199514
rect 145208 199306 145236 199736
rect 145564 199776 145616 199782
rect 145380 199718 145432 199724
rect 145470 199744 145526 199753
rect 145288 199708 145340 199714
rect 145288 199650 145340 199656
rect 145196 199300 145248 199306
rect 145196 199242 145248 199248
rect 145300 197713 145328 199650
rect 145392 198257 145420 199718
rect 145714 199764 145742 200124
rect 145564 199718 145616 199724
rect 145668 199736 145742 199764
rect 145806 199764 145834 200124
rect 145898 199889 145926 200124
rect 145884 199880 145940 199889
rect 145884 199815 145940 199824
rect 145990 199764 146018 200124
rect 146082 199918 146110 200124
rect 146174 199918 146202 200124
rect 146070 199912 146122 199918
rect 146070 199854 146122 199860
rect 146162 199912 146214 199918
rect 146162 199854 146214 199860
rect 145806 199736 145880 199764
rect 145470 199679 145526 199688
rect 145378 198248 145434 198257
rect 145378 198183 145434 198192
rect 145286 197704 145342 197713
rect 145286 197639 145342 197648
rect 145484 197538 145512 199679
rect 145472 197532 145524 197538
rect 145472 197474 145524 197480
rect 145576 197354 145604 199718
rect 145668 199442 145696 199736
rect 145746 199472 145802 199481
rect 145656 199436 145708 199442
rect 145746 199407 145802 199416
rect 145656 199378 145708 199384
rect 145760 197554 145788 199407
rect 145484 197326 145604 197354
rect 145668 197526 145788 197554
rect 145104 195288 145156 195294
rect 145104 195230 145156 195236
rect 145484 194041 145512 197326
rect 145668 197282 145696 197526
rect 145576 197254 145696 197282
rect 145470 194032 145526 194041
rect 145470 193967 145526 193976
rect 144736 193044 144788 193050
rect 144736 192986 144788 192992
rect 144642 183832 144698 183841
rect 144642 183767 144698 183776
rect 143816 144628 143868 144634
rect 143816 144570 143868 144576
rect 142526 144528 142582 144537
rect 142526 144463 142582 144472
rect 142066 142352 142122 142361
rect 142066 142287 142122 142296
rect 142252 141500 142304 141506
rect 142252 141442 142304 141448
rect 141606 141264 141662 141273
rect 141606 141199 141662 141208
rect 142264 139890 142292 141442
rect 142540 139890 142568 144463
rect 144182 144392 144238 144401
rect 144182 144327 144238 144336
rect 143078 143304 143134 143313
rect 143078 143239 143134 143248
rect 143092 139890 143120 143239
rect 143630 141672 143686 141681
rect 143630 141607 143686 141616
rect 143644 139890 143672 141607
rect 144196 139890 144224 144327
rect 145288 143608 145340 143614
rect 145288 143550 145340 143556
rect 145010 143032 145066 143041
rect 145010 142967 145066 142976
rect 145024 139890 145052 142967
rect 145300 139890 145328 143550
rect 145576 140282 145604 197254
rect 145656 190868 145708 190874
rect 145656 190810 145708 190816
rect 145668 147014 145696 190810
rect 145748 185020 145800 185026
rect 145748 184962 145800 184968
rect 145760 148617 145788 184962
rect 145852 179178 145880 199736
rect 145944 199736 146018 199764
rect 146116 199776 146168 199782
rect 145944 199238 145972 199736
rect 146266 199764 146294 200124
rect 146116 199718 146168 199724
rect 146220 199736 146294 199764
rect 146024 199640 146076 199646
rect 146024 199582 146076 199588
rect 145932 199232 145984 199238
rect 145932 199174 145984 199180
rect 146036 193662 146064 199582
rect 146024 193656 146076 193662
rect 146024 193598 146076 193604
rect 146128 191185 146156 199718
rect 146220 199073 146248 199736
rect 146358 199696 146386 200124
rect 146450 199918 146478 200124
rect 146438 199912 146490 199918
rect 146438 199854 146490 199860
rect 146542 199764 146570 200124
rect 146634 199918 146662 200124
rect 146622 199912 146674 199918
rect 146622 199854 146674 199860
rect 146726 199764 146754 200124
rect 146312 199668 146386 199696
rect 146496 199736 146570 199764
rect 146680 199736 146754 199764
rect 146818 199764 146846 200124
rect 146910 199918 146938 200124
rect 146898 199912 146950 199918
rect 146898 199854 146950 199860
rect 147002 199764 147030 200124
rect 147094 199918 147122 200124
rect 147186 199918 147214 200124
rect 147082 199912 147134 199918
rect 147082 199854 147134 199860
rect 147174 199912 147226 199918
rect 147174 199854 147226 199860
rect 147278 199764 147306 200124
rect 147370 199918 147398 200124
rect 147358 199912 147410 199918
rect 147358 199854 147410 199860
rect 147462 199764 147490 200124
rect 146818 199736 146892 199764
rect 147002 199736 147168 199764
rect 146206 199064 146262 199073
rect 146206 198999 146262 199008
rect 146114 191176 146170 191185
rect 146114 191111 146170 191120
rect 146312 182174 146340 199668
rect 146496 197985 146524 199736
rect 146576 199640 146628 199646
rect 146576 199582 146628 199588
rect 146482 197976 146538 197985
rect 146482 197911 146538 197920
rect 146588 197577 146616 199582
rect 146680 198626 146708 199736
rect 146864 199442 146892 199736
rect 146944 199640 146996 199646
rect 146944 199582 146996 199588
rect 147036 199640 147088 199646
rect 147036 199582 147088 199588
rect 146852 199436 146904 199442
rect 146852 199378 146904 199384
rect 146668 198620 146720 198626
rect 146668 198562 146720 198568
rect 146574 197568 146630 197577
rect 146574 197503 146630 197512
rect 146956 195673 146984 199582
rect 147048 198966 147076 199582
rect 147036 198960 147088 198966
rect 147036 198902 147088 198908
rect 146942 195664 146998 195673
rect 146942 195599 146998 195608
rect 147140 195566 147168 199736
rect 147232 199736 147306 199764
rect 147416 199736 147490 199764
rect 147554 199764 147582 200124
rect 147646 199918 147674 200124
rect 147634 199912 147686 199918
rect 147634 199854 147686 199860
rect 147738 199764 147766 200124
rect 147830 199918 147858 200124
rect 147818 199912 147870 199918
rect 147818 199854 147870 199860
rect 147554 199753 147628 199764
rect 147554 199744 147642 199753
rect 147554 199736 147586 199744
rect 147128 195560 147180 195566
rect 147128 195502 147180 195508
rect 147232 191185 147260 199736
rect 147312 199640 147364 199646
rect 147312 199582 147364 199588
rect 147218 191176 147274 191185
rect 146760 191140 146812 191146
rect 147324 191146 147352 199582
rect 147218 191111 147274 191120
rect 147312 191140 147364 191146
rect 146760 191082 146812 191088
rect 147312 191082 147364 191088
rect 146312 182146 146524 182174
rect 145840 179172 145892 179178
rect 145840 179114 145892 179120
rect 145746 148608 145802 148617
rect 145746 148543 145802 148552
rect 145656 147008 145708 147014
rect 145656 146950 145708 146956
rect 146496 145926 146524 182146
rect 146576 179172 146628 179178
rect 146576 179114 146628 179120
rect 146588 145994 146616 179114
rect 146772 151814 146800 191082
rect 147416 180794 147444 199736
rect 147586 199679 147642 199688
rect 147692 199736 147766 199764
rect 147588 199572 147640 199578
rect 147588 199514 147640 199520
rect 147600 199102 147628 199514
rect 147588 199096 147640 199102
rect 147588 199038 147640 199044
rect 147692 198830 147720 199736
rect 147772 199640 147824 199646
rect 147922 199628 147950 200124
rect 148014 199923 148042 200124
rect 148000 199914 148056 199923
rect 148106 199918 148134 200124
rect 148000 199849 148056 199858
rect 148094 199912 148146 199918
rect 148094 199854 148146 199860
rect 148048 199776 148100 199782
rect 148198 199764 148226 200124
rect 148290 199918 148318 200124
rect 148278 199912 148330 199918
rect 148278 199854 148330 199860
rect 148382 199764 148410 200124
rect 148474 199918 148502 200124
rect 148462 199912 148514 199918
rect 148462 199854 148514 199860
rect 148566 199764 148594 200124
rect 148658 199923 148686 200124
rect 148644 199914 148700 199923
rect 148750 199918 148778 200124
rect 148842 199918 148870 200124
rect 148934 199918 148962 200124
rect 148644 199849 148700 199858
rect 148738 199912 148790 199918
rect 148738 199854 148790 199860
rect 148830 199912 148882 199918
rect 148830 199854 148882 199860
rect 148922 199912 148974 199918
rect 148922 199854 148974 199860
rect 148048 199718 148100 199724
rect 148152 199736 148226 199764
rect 148336 199736 148410 199764
rect 148520 199736 148594 199764
rect 148692 199776 148744 199782
rect 147922 199600 147996 199628
rect 147772 199582 147824 199588
rect 147680 198824 147732 198830
rect 147680 198766 147732 198772
rect 147784 197713 147812 199582
rect 147770 197704 147826 197713
rect 147770 197639 147826 197648
rect 147680 197532 147732 197538
rect 147680 197474 147732 197480
rect 147588 197124 147640 197130
rect 147588 197066 147640 197072
rect 147048 180766 147444 180794
rect 146772 151786 146984 151814
rect 146668 146124 146720 146130
rect 146668 146066 146720 146072
rect 146576 145988 146628 145994
rect 146576 145930 146628 145936
rect 146484 145920 146536 145926
rect 146484 145862 146536 145868
rect 146298 145752 146354 145761
rect 146298 145687 146354 145696
rect 145838 144256 145894 144265
rect 145838 144191 145894 144200
rect 145564 140276 145616 140282
rect 145564 140218 145616 140224
rect 145852 139890 145880 144191
rect 146312 143478 146340 145687
rect 146300 143472 146352 143478
rect 146300 143414 146352 143420
rect 146390 143168 146446 143177
rect 146390 143103 146446 143112
rect 146404 139890 146432 143103
rect 146680 140706 146708 146066
rect 146680 140678 146892 140706
rect 146864 139890 146892 140678
rect 146956 140418 146984 151786
rect 147048 140486 147076 180766
rect 147600 146985 147628 197066
rect 147586 146976 147642 146985
rect 147586 146911 147642 146920
rect 147692 145858 147720 197474
rect 147968 196246 147996 199600
rect 147956 196240 148008 196246
rect 147956 196182 148008 196188
rect 148060 195537 148088 199718
rect 148152 199374 148180 199736
rect 148232 199640 148284 199646
rect 148232 199582 148284 199588
rect 148140 199368 148192 199374
rect 148140 199310 148192 199316
rect 148244 198354 148272 199582
rect 148232 198348 148284 198354
rect 148232 198290 148284 198296
rect 148336 195974 148364 199736
rect 148416 199640 148468 199646
rect 148416 199582 148468 199588
rect 148428 199170 148456 199582
rect 148416 199164 148468 199170
rect 148416 199106 148468 199112
rect 148244 195946 148364 195974
rect 148046 195528 148102 195537
rect 148046 195463 148102 195472
rect 148244 195344 148272 195946
rect 147968 195316 148272 195344
rect 147968 193730 147996 195316
rect 148520 195276 148548 199736
rect 148692 199718 148744 199724
rect 148784 199776 148836 199782
rect 149026 199764 149054 200124
rect 149118 199918 149146 200124
rect 149106 199912 149158 199918
rect 149106 199854 149158 199860
rect 149210 199764 149238 200124
rect 148784 199718 148836 199724
rect 148980 199736 149054 199764
rect 149164 199736 149238 199764
rect 149302 199764 149330 200124
rect 149394 199918 149422 200124
rect 149382 199912 149434 199918
rect 149382 199854 149434 199860
rect 149486 199764 149514 200124
rect 149578 199918 149606 200124
rect 149566 199912 149618 199918
rect 149670 199889 149698 200124
rect 149566 199854 149618 199860
rect 149656 199880 149712 199889
rect 149656 199815 149712 199824
rect 149612 199776 149664 199782
rect 149302 199736 149376 199764
rect 149486 199736 149560 199764
rect 148704 198744 148732 199718
rect 148612 198716 148732 198744
rect 148612 197062 148640 198716
rect 148600 197056 148652 197062
rect 148600 196998 148652 197004
rect 148060 195248 148548 195276
rect 147956 193724 148008 193730
rect 147956 193666 148008 193672
rect 148060 151814 148088 195248
rect 148796 195158 148824 199718
rect 148876 199640 148928 199646
rect 148876 199582 148928 199588
rect 148888 198801 148916 199582
rect 148874 198792 148930 198801
rect 148874 198727 148930 198736
rect 148980 195226 149008 199736
rect 149164 198218 149192 199736
rect 149244 199504 149296 199510
rect 149244 199446 149296 199452
rect 149152 198212 149204 198218
rect 149152 198154 149204 198160
rect 149058 196072 149114 196081
rect 149058 196007 149114 196016
rect 148968 195220 149020 195226
rect 148968 195162 149020 195168
rect 148232 195152 148284 195158
rect 148232 195094 148284 195100
rect 148784 195152 148836 195158
rect 148784 195094 148836 195100
rect 147968 151786 148088 151814
rect 147680 145852 147732 145858
rect 147680 145794 147732 145800
rect 147678 145616 147734 145625
rect 147678 145551 147734 145560
rect 147036 140480 147088 140486
rect 147036 140422 147088 140428
rect 146944 140412 146996 140418
rect 146944 140354 146996 140360
rect 147692 139890 147720 145551
rect 147968 140214 147996 151786
rect 148046 142896 148102 142905
rect 148046 142831 148102 142840
rect 147956 140208 148008 140214
rect 147956 140150 148008 140156
rect 148060 139890 148088 142831
rect 148244 140350 148272 195094
rect 148692 185836 148744 185842
rect 148692 185778 148744 185784
rect 148704 180794 148732 185778
rect 149072 182174 149100 196007
rect 149256 195809 149284 199446
rect 149348 198801 149376 199736
rect 149334 198792 149390 198801
rect 149334 198727 149390 198736
rect 149532 198370 149560 199736
rect 149612 199718 149664 199724
rect 149762 199730 149790 200124
rect 149854 199918 149882 200124
rect 149946 199918 149974 200124
rect 149842 199912 149894 199918
rect 149842 199854 149894 199860
rect 149934 199912 149986 199918
rect 150038 199889 150066 200124
rect 150130 199918 150158 200124
rect 150118 199912 150170 199918
rect 149934 199854 149986 199860
rect 150024 199880 150080 199889
rect 150118 199854 150170 199860
rect 150024 199815 150080 199824
rect 149888 199776 149940 199782
rect 149440 198342 149560 198370
rect 149440 197878 149468 198342
rect 149428 197872 149480 197878
rect 149428 197814 149480 197820
rect 149624 197354 149652 199718
rect 149762 199702 149836 199730
rect 150072 199776 150124 199782
rect 149888 199718 149940 199724
rect 150070 199744 150072 199753
rect 150222 199764 150250 200124
rect 150314 199918 150342 200124
rect 150406 199918 150434 200124
rect 150498 199923 150526 200124
rect 150302 199912 150354 199918
rect 150302 199854 150354 199860
rect 150394 199912 150446 199918
rect 150394 199854 150446 199860
rect 150484 199914 150540 199923
rect 150484 199849 150540 199858
rect 150590 199764 150618 200124
rect 150682 199918 150710 200124
rect 150774 199918 150802 200124
rect 150866 199918 150894 200124
rect 150958 199918 150986 200124
rect 150670 199912 150722 199918
rect 150670 199854 150722 199860
rect 150762 199912 150814 199918
rect 150762 199854 150814 199860
rect 150854 199912 150906 199918
rect 150854 199854 150906 199860
rect 150946 199912 150998 199918
rect 150946 199854 150998 199860
rect 150124 199744 150126 199753
rect 149532 197326 149652 197354
rect 149242 195800 149298 195809
rect 149242 195735 149298 195744
rect 149532 195344 149560 197326
rect 149702 195528 149758 195537
rect 149702 195463 149758 195472
rect 149440 195316 149560 195344
rect 149440 194546 149468 195316
rect 149428 194540 149480 194546
rect 149428 194482 149480 194488
rect 149716 189514 149744 195463
rect 149808 192778 149836 199702
rect 149796 192772 149848 192778
rect 149796 192714 149848 192720
rect 149704 189508 149756 189514
rect 149704 189450 149756 189456
rect 149704 189372 149756 189378
rect 149704 189314 149756 189320
rect 149520 186380 149572 186386
rect 149520 186322 149572 186328
rect 148336 180766 148732 180794
rect 148980 182146 149100 182174
rect 148336 148170 148364 180766
rect 148980 149734 149008 182146
rect 148968 149728 149020 149734
rect 148968 149670 149020 149676
rect 148324 148164 148376 148170
rect 148324 148106 148376 148112
rect 149532 146062 149560 186322
rect 149716 151814 149744 189314
rect 149900 180334 149928 199718
rect 150070 199679 150126 199688
rect 150176 199736 150250 199764
rect 150544 199736 150618 199764
rect 150716 199776 150768 199782
rect 150072 199572 150124 199578
rect 150072 199514 150124 199520
rect 149978 195528 150034 195537
rect 149978 195463 150034 195472
rect 149992 188465 150020 195463
rect 149978 188456 150034 188465
rect 149978 188391 150034 188400
rect 150084 187474 150112 199514
rect 150072 187468 150124 187474
rect 150072 187410 150124 187416
rect 150176 186386 150204 199736
rect 150348 199708 150400 199714
rect 150348 199650 150400 199656
rect 150256 199640 150308 199646
rect 150256 199582 150308 199588
rect 150268 198830 150296 199582
rect 150256 198824 150308 198830
rect 150256 198766 150308 198772
rect 150360 195129 150388 199650
rect 150544 197334 150572 199736
rect 151050 199764 151078 200124
rect 151142 199889 151170 200124
rect 151234 199918 151262 200124
rect 151326 199918 151354 200124
rect 151418 199918 151446 200124
rect 151510 199923 151538 200124
rect 151222 199912 151274 199918
rect 151128 199880 151184 199889
rect 151222 199854 151274 199860
rect 151314 199912 151366 199918
rect 151314 199854 151366 199860
rect 151406 199912 151458 199918
rect 151406 199854 151458 199860
rect 151496 199914 151552 199923
rect 151496 199849 151552 199858
rect 151128 199815 151184 199824
rect 151602 199764 151630 200124
rect 150716 199718 150768 199724
rect 151004 199736 151078 199764
rect 151556 199736 151630 199764
rect 150532 197328 150584 197334
rect 150532 197270 150584 197276
rect 150728 195265 150756 199718
rect 150806 199608 150862 199617
rect 150806 199543 150862 199552
rect 150820 199374 150848 199543
rect 150808 199368 150860 199374
rect 150808 199310 150860 199316
rect 150714 195256 150770 195265
rect 150714 195191 150770 195200
rect 150346 195120 150402 195129
rect 150346 195055 150402 195064
rect 150532 191208 150584 191214
rect 150346 191176 150402 191185
rect 150532 191150 150584 191156
rect 150346 191111 150402 191120
rect 150164 186380 150216 186386
rect 150164 186322 150216 186328
rect 149888 180328 149940 180334
rect 149888 180270 149940 180276
rect 149624 151786 149744 151814
rect 149520 146056 149572 146062
rect 149520 145998 149572 146004
rect 148600 144356 148652 144362
rect 148600 144298 148652 144304
rect 148232 140344 148284 140350
rect 148232 140286 148284 140292
rect 148612 139890 148640 144298
rect 149152 143472 149204 143478
rect 149152 143414 149204 143420
rect 149164 139890 149192 143414
rect 132328 139862 132388 139890
rect 132604 139862 132940 139890
rect 133156 139862 133492 139890
rect 133892 139862 134044 139890
rect 134260 139862 134596 139890
rect 134812 139862 135148 139890
rect 135456 139862 135700 139890
rect 135916 139862 136252 139890
rect 136652 139862 136804 139890
rect 137020 139862 137356 139890
rect 137572 139862 137908 139890
rect 138124 139862 138460 139890
rect 138676 139862 139012 139890
rect 139412 139862 139564 139890
rect 139780 139862 140116 139890
rect 140332 139862 140668 139890
rect 140884 139862 141220 139890
rect 141528 139862 141772 139890
rect 142264 139862 142324 139890
rect 142540 139862 142876 139890
rect 143092 139862 143428 139890
rect 143644 139862 143980 139890
rect 144196 139862 144532 139890
rect 145024 139862 145084 139890
rect 145300 139862 145636 139890
rect 145852 139862 146188 139890
rect 146404 139862 146740 139890
rect 146864 139862 147292 139890
rect 147692 139862 147844 139890
rect 148060 139862 148396 139890
rect 148612 139862 148948 139890
rect 149164 139862 149500 139890
rect 149624 139369 149652 151786
rect 150360 149705 150388 191111
rect 150346 149696 150402 149705
rect 150346 149631 150402 149640
rect 150544 144430 150572 191150
rect 151004 190454 151032 199736
rect 151556 199730 151584 199736
rect 151176 199708 151228 199714
rect 151176 199650 151228 199656
rect 151464 199702 151584 199730
rect 151084 199640 151136 199646
rect 151084 199582 151136 199588
rect 151096 199306 151124 199582
rect 151084 199300 151136 199306
rect 151084 199242 151136 199248
rect 151188 197946 151216 199650
rect 151360 199572 151412 199578
rect 151360 199514 151412 199520
rect 151268 199504 151320 199510
rect 151268 199446 151320 199452
rect 151176 197940 151228 197946
rect 151176 197882 151228 197888
rect 151280 193866 151308 199446
rect 151268 193860 151320 193866
rect 151268 193802 151320 193808
rect 150912 190426 151032 190454
rect 150912 180794 150940 190426
rect 150992 189916 151044 189922
rect 150992 189858 151044 189864
rect 150636 180766 150940 180794
rect 150636 145722 150664 180766
rect 150624 145716 150676 145722
rect 150624 145658 150676 145664
rect 150532 144424 150584 144430
rect 150532 144366 150584 144372
rect 149702 142760 149758 142769
rect 149702 142695 149758 142704
rect 149716 139890 149744 142695
rect 150438 141400 150494 141409
rect 150438 141335 150494 141344
rect 150452 139890 150480 141335
rect 149716 139862 150052 139890
rect 150452 139862 150604 139890
rect 151004 139369 151032 189858
rect 151372 182174 151400 199514
rect 151464 199442 151492 199702
rect 151694 199696 151722 200124
rect 151786 199918 151814 200124
rect 151878 199918 151906 200124
rect 151970 199918 151998 200124
rect 151774 199912 151826 199918
rect 151774 199854 151826 199860
rect 151866 199912 151918 199918
rect 151866 199854 151918 199860
rect 151958 199912 152010 199918
rect 151958 199854 152010 199860
rect 151820 199776 151872 199782
rect 152062 199764 152090 200124
rect 152154 199918 152182 200124
rect 152142 199912 152194 199918
rect 152142 199854 152194 199860
rect 152246 199764 152274 200124
rect 152338 199889 152366 200124
rect 152324 199880 152380 199889
rect 152324 199815 152380 199824
rect 152062 199736 152136 199764
rect 151820 199718 151872 199724
rect 151648 199668 151722 199696
rect 151544 199640 151596 199646
rect 151544 199582 151596 199588
rect 151452 199436 151504 199442
rect 151452 199378 151504 199384
rect 151556 195945 151584 199582
rect 151542 195936 151598 195945
rect 151542 195871 151598 195880
rect 151648 189922 151676 199668
rect 151832 199560 151860 199718
rect 151912 199708 151964 199714
rect 151912 199650 151964 199656
rect 151740 199532 151860 199560
rect 151740 191146 151768 199532
rect 151820 199436 151872 199442
rect 151820 199378 151872 199384
rect 151832 191214 151860 199378
rect 151820 191208 151872 191214
rect 151820 191150 151872 191156
rect 151728 191140 151780 191146
rect 151728 191082 151780 191088
rect 151924 190874 151952 199650
rect 152004 199640 152056 199646
rect 152108 199617 152136 199736
rect 152200 199736 152274 199764
rect 152004 199582 152056 199588
rect 152094 199608 152150 199617
rect 152016 195906 152044 199582
rect 152094 199543 152150 199552
rect 152200 198734 152228 199736
rect 152430 199730 152458 200124
rect 152384 199702 152458 199730
rect 152522 199730 152550 200124
rect 152614 199889 152642 200124
rect 152600 199880 152656 199889
rect 152706 199850 152734 200124
rect 152798 199850 152826 200124
rect 152600 199815 152656 199824
rect 152694 199844 152746 199850
rect 152694 199786 152746 199792
rect 152786 199844 152838 199850
rect 152786 199786 152838 199792
rect 152890 199730 152918 200124
rect 152982 199850 153010 200124
rect 153074 199918 153102 200124
rect 153062 199912 153114 199918
rect 153062 199854 153114 199860
rect 152970 199844 153022 199850
rect 152970 199786 153022 199792
rect 153166 199730 153194 200124
rect 153258 199918 153286 200124
rect 153350 199918 153378 200124
rect 153246 199912 153298 199918
rect 153246 199854 153298 199860
rect 153338 199912 153390 199918
rect 153338 199854 153390 199860
rect 153442 199764 153470 200124
rect 153534 199918 153562 200124
rect 153522 199912 153574 199918
rect 153522 199854 153574 199860
rect 153626 199764 153654 200124
rect 153718 199918 153746 200124
rect 153810 199918 153838 200124
rect 153706 199912 153758 199918
rect 153706 199854 153758 199860
rect 153798 199912 153850 199918
rect 153798 199854 153850 199860
rect 152522 199702 152596 199730
rect 152280 199504 152332 199510
rect 152280 199446 152332 199452
rect 152108 198706 152228 198734
rect 152004 195900 152056 195906
rect 152004 195842 152056 195848
rect 152108 191593 152136 198706
rect 152292 194177 152320 199446
rect 152278 194168 152334 194177
rect 152278 194103 152334 194112
rect 152094 191584 152150 191593
rect 152094 191519 152150 191528
rect 152384 191298 152412 199702
rect 152464 199572 152516 199578
rect 152464 199514 152516 199520
rect 152476 199209 152504 199514
rect 152462 199200 152518 199209
rect 152462 199135 152518 199144
rect 152108 191270 152412 191298
rect 151912 190868 151964 190874
rect 151912 190810 151964 190816
rect 151912 190732 151964 190738
rect 151912 190674 151964 190680
rect 151636 189916 151688 189922
rect 151636 189858 151688 189864
rect 151372 182146 151768 182174
rect 151740 148442 151768 182146
rect 151728 148436 151780 148442
rect 151728 148378 151780 148384
rect 151082 144120 151138 144129
rect 151082 144055 151138 144064
rect 151096 139890 151124 144055
rect 151360 142860 151412 142866
rect 151360 142802 151412 142808
rect 151372 139890 151400 142802
rect 151924 141574 151952 190674
rect 152108 148850 152136 191270
rect 152188 191140 152240 191146
rect 152188 191082 152240 191088
rect 152096 148844 152148 148850
rect 152096 148786 152148 148792
rect 152200 148510 152228 191082
rect 152568 188873 152596 199702
rect 152844 199702 152918 199730
rect 153120 199702 153194 199730
rect 153396 199736 153470 199764
rect 153580 199736 153654 199764
rect 153902 199764 153930 200124
rect 153994 199889 154022 200124
rect 154086 199918 154114 200124
rect 154074 199912 154126 199918
rect 153980 199880 154036 199889
rect 154074 199854 154126 199860
rect 153980 199815 154036 199824
rect 154178 199764 154206 200124
rect 154270 199918 154298 200124
rect 154362 199923 154390 200124
rect 154258 199912 154310 199918
rect 154258 199854 154310 199860
rect 154348 199914 154404 199923
rect 154348 199849 154404 199858
rect 153902 199736 153976 199764
rect 152648 199572 152700 199578
rect 152648 199514 152700 199520
rect 152660 195974 152688 199514
rect 152844 199170 152872 199702
rect 152924 199640 152976 199646
rect 152924 199582 152976 199588
rect 152832 199164 152884 199170
rect 152832 199106 152884 199112
rect 152660 195946 152780 195974
rect 152648 195900 152700 195906
rect 152648 195842 152700 195848
rect 152660 190738 152688 195842
rect 152648 190732 152700 190738
rect 152648 190674 152700 190680
rect 152554 188864 152610 188873
rect 152554 188799 152610 188808
rect 152752 187377 152780 195946
rect 152738 187368 152794 187377
rect 152738 187303 152794 187312
rect 152936 180794 152964 199582
rect 153016 199436 153068 199442
rect 153016 199378 153068 199384
rect 153028 182174 153056 199378
rect 153120 195498 153148 199702
rect 153200 199572 153252 199578
rect 153200 199514 153252 199520
rect 153108 195492 153160 195498
rect 153108 195434 153160 195440
rect 153212 189378 153240 199514
rect 153292 199436 153344 199442
rect 153292 199378 153344 199384
rect 153304 197305 153332 199378
rect 153396 198150 153424 199736
rect 153476 199640 153528 199646
rect 153476 199582 153528 199588
rect 153384 198144 153436 198150
rect 153384 198086 153436 198092
rect 153290 197296 153346 197305
rect 153290 197231 153346 197240
rect 153488 197180 153516 199582
rect 153580 197305 153608 199736
rect 153752 199708 153804 199714
rect 153752 199650 153804 199656
rect 153660 199640 153712 199646
rect 153660 199582 153712 199588
rect 153566 197296 153622 197305
rect 153566 197231 153622 197240
rect 153304 197152 153516 197180
rect 153200 189372 153252 189378
rect 153200 189314 153252 189320
rect 153028 182146 153148 182174
rect 152568 180766 152964 180794
rect 152568 151814 152596 180766
rect 152476 151786 152596 151814
rect 152188 148504 152240 148510
rect 152188 148446 152240 148452
rect 151912 141568 151964 141574
rect 151912 141510 151964 141516
rect 152476 140146 152504 151786
rect 153120 145790 153148 182146
rect 153304 148578 153332 197152
rect 153672 195265 153700 199582
rect 153764 199345 153792 199650
rect 153948 199646 153976 199736
rect 154086 199736 154206 199764
rect 154304 199776 154356 199782
rect 154086 199730 154114 199736
rect 154040 199702 154114 199730
rect 154454 199764 154482 200124
rect 154546 199918 154574 200124
rect 154534 199912 154586 199918
rect 154534 199854 154586 199860
rect 154304 199718 154356 199724
rect 154408 199736 154482 199764
rect 153936 199640 153988 199646
rect 154040 199617 154068 199702
rect 153936 199582 153988 199588
rect 154026 199608 154082 199617
rect 153844 199572 153896 199578
rect 154026 199543 154082 199552
rect 153844 199514 153896 199520
rect 153750 199336 153806 199345
rect 153750 199271 153806 199280
rect 153658 195256 153714 195265
rect 153658 195191 153714 195200
rect 153384 192976 153436 192982
rect 153384 192918 153436 192924
rect 153292 148572 153344 148578
rect 153292 148514 153344 148520
rect 153396 148481 153424 192918
rect 153476 184748 153528 184754
rect 153476 184690 153528 184696
rect 153488 148918 153516 184690
rect 153476 148912 153528 148918
rect 153476 148854 153528 148860
rect 153382 148472 153438 148481
rect 153382 148407 153438 148416
rect 153108 145784 153160 145790
rect 153108 145726 153160 145732
rect 153290 145616 153346 145625
rect 153290 145551 153346 145560
rect 152648 144560 152700 144566
rect 152648 144502 152700 144508
rect 152556 144424 152608 144430
rect 152556 144366 152608 144372
rect 152464 140140 152516 140146
rect 152464 140082 152516 140088
rect 152568 139890 152596 144366
rect 151096 139862 151156 139890
rect 151372 139862 151708 139890
rect 152260 139862 152596 139890
rect 152660 139890 152688 144502
rect 153304 139890 153332 145551
rect 153856 144498 153884 199514
rect 153936 199504 153988 199510
rect 153936 199446 153988 199452
rect 154028 199504 154080 199510
rect 154028 199446 154080 199452
rect 153948 194002 153976 199446
rect 153936 193996 153988 194002
rect 153936 193938 153988 193944
rect 154040 192982 154068 199446
rect 154316 195974 154344 199718
rect 154304 195968 154356 195974
rect 154304 195910 154356 195916
rect 154408 195537 154436 199736
rect 154638 199696 154666 200124
rect 154730 199918 154758 200124
rect 154822 199923 154850 200124
rect 154718 199912 154770 199918
rect 154718 199854 154770 199860
rect 154808 199914 154864 199923
rect 154808 199849 154864 199858
rect 154914 199730 154942 200124
rect 155006 199918 155034 200124
rect 155098 199918 155126 200124
rect 155190 199918 155218 200124
rect 155282 199923 155310 200124
rect 154994 199912 155046 199918
rect 154994 199854 155046 199860
rect 155086 199912 155138 199918
rect 155086 199854 155138 199860
rect 155178 199912 155230 199918
rect 155178 199854 155230 199860
rect 155268 199914 155324 199923
rect 155374 199918 155402 200124
rect 155466 199918 155494 200124
rect 155268 199849 155324 199858
rect 155362 199912 155414 199918
rect 155362 199854 155414 199860
rect 155454 199912 155506 199918
rect 155454 199854 155506 199860
rect 155224 199776 155276 199782
rect 154592 199668 154666 199696
rect 154764 199708 154816 199714
rect 154394 195528 154450 195537
rect 154394 195463 154450 195472
rect 154302 195256 154358 195265
rect 154302 195191 154358 195200
rect 154028 192976 154080 192982
rect 154028 192918 154080 192924
rect 154316 184754 154344 195191
rect 154592 185842 154620 199668
rect 154764 199650 154816 199656
rect 154868 199702 154942 199730
rect 155144 199736 155224 199764
rect 154672 199572 154724 199578
rect 154672 199514 154724 199520
rect 154684 199481 154712 199514
rect 154670 199472 154726 199481
rect 154670 199407 154726 199416
rect 154776 198734 154804 199650
rect 154684 198706 154804 198734
rect 154684 197169 154712 198706
rect 154670 197160 154726 197169
rect 154868 197130 154896 199702
rect 155040 199504 155092 199510
rect 155040 199446 155092 199452
rect 155052 197878 155080 199446
rect 155040 197872 155092 197878
rect 155040 197814 155092 197820
rect 154670 197095 154726 197104
rect 154856 197124 154908 197130
rect 154856 197066 154908 197072
rect 155144 191162 155172 199736
rect 155408 199776 155460 199782
rect 155224 199718 155276 199724
rect 155314 199744 155370 199753
rect 155558 199764 155586 200124
rect 155512 199753 155586 199764
rect 155408 199718 155460 199724
rect 155498 199744 155586 199753
rect 155314 199679 155370 199688
rect 155328 199578 155356 199679
rect 155316 199572 155368 199578
rect 155316 199514 155368 199520
rect 155420 198734 155448 199718
rect 155554 199736 155586 199744
rect 155498 199679 155554 199688
rect 155650 199696 155678 200124
rect 155742 199764 155770 200124
rect 155834 199918 155862 200124
rect 155822 199912 155874 199918
rect 155822 199854 155874 199860
rect 155926 199764 155954 200124
rect 156018 199889 156046 200124
rect 156110 199918 156138 200124
rect 156098 199912 156150 199918
rect 156004 199880 156060 199889
rect 156098 199854 156150 199860
rect 156004 199815 156060 199824
rect 156202 199764 156230 200124
rect 156294 199850 156322 200124
rect 156386 199889 156414 200124
rect 156478 199918 156506 200124
rect 156466 199912 156518 199918
rect 156372 199880 156428 199889
rect 156282 199844 156334 199850
rect 156466 199854 156518 199860
rect 156372 199815 156428 199824
rect 156282 199786 156334 199792
rect 156570 199764 156598 200124
rect 156662 199918 156690 200124
rect 156754 199918 156782 200124
rect 156846 199923 156874 200124
rect 156650 199912 156702 199918
rect 156650 199854 156702 199860
rect 156742 199912 156794 199918
rect 156742 199854 156794 199860
rect 156832 199914 156888 199923
rect 156938 199918 156966 200124
rect 156832 199849 156888 199858
rect 156926 199912 156978 199918
rect 156926 199854 156978 199860
rect 155742 199753 155816 199764
rect 155742 199744 155830 199753
rect 155742 199736 155774 199744
rect 155650 199668 155724 199696
rect 155926 199736 156092 199764
rect 155774 199679 155830 199688
rect 155592 199504 155644 199510
rect 155696 199481 155724 199668
rect 155776 199640 155828 199646
rect 155776 199582 155828 199588
rect 155960 199640 156012 199646
rect 155960 199582 156012 199588
rect 155592 199446 155644 199452
rect 155682 199472 155738 199481
rect 155420 198706 155540 198734
rect 154868 191134 155172 191162
rect 154764 188828 154816 188834
rect 154764 188770 154816 188776
rect 154580 185836 154632 185842
rect 154580 185778 154632 185784
rect 154304 184748 154356 184754
rect 154304 184690 154356 184696
rect 154776 147257 154804 188770
rect 154868 149054 154896 191134
rect 154946 189952 155002 189961
rect 154946 189887 155002 189896
rect 154960 149841 154988 189887
rect 155512 188834 155540 198706
rect 155500 188828 155552 188834
rect 155500 188770 155552 188776
rect 155604 182174 155632 199446
rect 155682 199407 155738 199416
rect 155604 182146 155724 182174
rect 155696 151814 155724 182146
rect 155236 151786 155724 151814
rect 154946 149832 155002 149841
rect 154946 149767 155002 149776
rect 154856 149048 154908 149054
rect 154856 148990 154908 148996
rect 154762 147248 154818 147257
rect 154762 147183 154818 147192
rect 153844 144492 153896 144498
rect 153844 144434 153896 144440
rect 154486 144392 154542 144401
rect 154486 144327 154542 144336
rect 153568 141432 153620 141438
rect 153568 141374 153620 141380
rect 153580 139890 153608 141374
rect 154500 140162 154528 144327
rect 155130 142896 155186 142905
rect 155130 142831 155186 142840
rect 154454 140134 154528 140162
rect 152660 139862 152812 139890
rect 153304 139862 153364 139890
rect 153580 139862 153916 139890
rect 154454 139876 154482 140134
rect 155144 139890 155172 142831
rect 155020 139862 155172 139890
rect 155236 139369 155264 151786
rect 155684 142248 155736 142254
rect 155684 142190 155736 142196
rect 155696 139890 155724 142190
rect 155572 139862 155724 139890
rect 155788 139369 155816 199582
rect 155868 199572 155920 199578
rect 155868 199514 155920 199520
rect 155880 195945 155908 199514
rect 155972 199374 156000 199582
rect 155960 199368 156012 199374
rect 155960 199310 156012 199316
rect 156064 198812 156092 199736
rect 156156 199736 156230 199764
rect 156326 199744 156382 199753
rect 156156 199646 156184 199736
rect 156524 199736 156598 199764
rect 156880 199776 156932 199782
rect 156326 199679 156382 199688
rect 156420 199708 156472 199714
rect 156144 199640 156196 199646
rect 156144 199582 156196 199588
rect 156236 199640 156288 199646
rect 156236 199582 156288 199588
rect 156144 199436 156196 199442
rect 156144 199378 156196 199384
rect 156156 199238 156184 199378
rect 156144 199232 156196 199238
rect 156144 199174 156196 199180
rect 156064 198801 156184 198812
rect 155958 198792 156014 198801
rect 156064 198792 156198 198801
rect 156064 198784 156142 198792
rect 155958 198734 156014 198736
rect 155958 198727 156092 198734
rect 156142 198727 156198 198736
rect 155972 198706 156092 198727
rect 155866 195936 155922 195945
rect 155866 195871 155922 195880
rect 156064 147393 156092 198706
rect 156248 192438 156276 199582
rect 156340 193186 156368 199679
rect 156420 199650 156472 199656
rect 156432 198218 156460 199650
rect 156420 198212 156472 198218
rect 156420 198154 156472 198160
rect 156328 193180 156380 193186
rect 156328 193122 156380 193128
rect 156236 192432 156288 192438
rect 156236 192374 156288 192380
rect 156524 185026 156552 199736
rect 156880 199718 156932 199724
rect 156604 199640 156656 199646
rect 156604 199582 156656 199588
rect 156616 197441 156644 199582
rect 156696 199572 156748 199578
rect 156696 199514 156748 199520
rect 156708 198490 156736 199514
rect 156892 199424 156920 199718
rect 157030 199696 157058 200124
rect 157122 199918 157150 200124
rect 157110 199912 157162 199918
rect 157110 199854 157162 199860
rect 157214 199764 157242 200124
rect 157306 199918 157334 200124
rect 157398 199918 157426 200124
rect 157294 199912 157346 199918
rect 157294 199854 157346 199860
rect 157386 199912 157438 199918
rect 157386 199854 157438 199860
rect 157490 199764 157518 200124
rect 156800 199396 156920 199424
rect 156984 199668 157058 199696
rect 157168 199736 157242 199764
rect 157444 199736 157518 199764
rect 156696 198484 156748 198490
rect 156696 198426 156748 198432
rect 156800 198393 156828 199396
rect 156878 199336 156934 199345
rect 156878 199271 156934 199280
rect 156786 198384 156842 198393
rect 156786 198319 156842 198328
rect 156892 198200 156920 199271
rect 156800 198172 156920 198200
rect 156602 197432 156658 197441
rect 156602 197367 156658 197376
rect 156512 185020 156564 185026
rect 156512 184962 156564 184968
rect 156800 180794 156828 198172
rect 156984 195838 157012 199668
rect 157064 199572 157116 199578
rect 157064 199514 157116 199520
rect 156972 195832 157024 195838
rect 156972 195774 157024 195780
rect 157076 180794 157104 199514
rect 157168 199481 157196 199736
rect 157340 199708 157392 199714
rect 157340 199650 157392 199656
rect 157248 199640 157300 199646
rect 157248 199582 157300 199588
rect 157154 199472 157210 199481
rect 157154 199407 157210 199416
rect 157154 199336 157210 199345
rect 157154 199271 157156 199280
rect 157208 199271 157210 199280
rect 157156 199242 157208 199248
rect 157260 195294 157288 199582
rect 157352 195430 157380 199650
rect 157444 198914 157472 199736
rect 157582 199696 157610 200124
rect 157674 199918 157702 200124
rect 157662 199912 157714 199918
rect 157766 199889 157794 200124
rect 157662 199854 157714 199860
rect 157752 199880 157808 199889
rect 157752 199815 157808 199824
rect 157858 199764 157886 200124
rect 157950 199918 157978 200124
rect 157938 199912 157990 199918
rect 157938 199854 157990 199860
rect 158042 199764 158070 200124
rect 157858 199736 157932 199764
rect 157582 199668 157656 199696
rect 157444 198886 157564 198914
rect 157432 198824 157484 198830
rect 157432 198766 157484 198772
rect 157444 198121 157472 198766
rect 157430 198112 157486 198121
rect 157430 198047 157486 198056
rect 157340 195424 157392 195430
rect 157340 195366 157392 195372
rect 157248 195288 157300 195294
rect 157248 195230 157300 195236
rect 157536 192370 157564 198886
rect 157628 198014 157656 199668
rect 157904 198558 157932 199736
rect 157996 199736 158070 199764
rect 157892 198552 157944 198558
rect 157892 198494 157944 198500
rect 157616 198008 157668 198014
rect 157616 197950 157668 197956
rect 157892 196240 157944 196246
rect 157892 196182 157944 196188
rect 157800 195288 157852 195294
rect 157800 195230 157852 195236
rect 157524 192364 157576 192370
rect 157524 192306 157576 192312
rect 157432 192296 157484 192302
rect 157432 192238 157484 192244
rect 157248 190256 157300 190262
rect 157248 190198 157300 190204
rect 156156 180766 156828 180794
rect 156984 180766 157104 180794
rect 156156 148714 156184 180766
rect 156984 151814 157012 180766
rect 156984 151786 157104 151814
rect 156144 148708 156196 148714
rect 156144 148650 156196 148656
rect 156050 147384 156106 147393
rect 156050 147319 156106 147328
rect 156420 144356 156472 144362
rect 156420 144298 156472 144304
rect 156432 139890 156460 144298
rect 156970 142760 157026 142769
rect 156970 142695 157026 142704
rect 156984 139890 157012 142695
rect 157076 140185 157104 151786
rect 157260 149977 157288 190198
rect 157444 150249 157472 192238
rect 157616 191140 157668 191146
rect 157616 191082 157668 191088
rect 157628 150385 157656 191082
rect 157614 150376 157670 150385
rect 157614 150311 157670 150320
rect 157430 150240 157486 150249
rect 157430 150175 157486 150184
rect 157246 149968 157302 149977
rect 157246 149903 157302 149912
rect 157812 149569 157840 195230
rect 157904 190454 157932 196182
rect 157996 194041 158024 199736
rect 158134 199696 158162 200124
rect 158226 199918 158254 200124
rect 158318 199923 158346 200124
rect 158214 199912 158266 199918
rect 158214 199854 158266 199860
rect 158304 199914 158360 199923
rect 158304 199849 158360 199858
rect 158088 199668 158162 199696
rect 158258 199744 158314 199753
rect 158410 199730 158438 200124
rect 158502 199918 158530 200124
rect 158490 199912 158542 199918
rect 158490 199854 158542 199860
rect 158314 199702 158438 199730
rect 158594 199696 158622 200124
rect 158258 199679 158314 199688
rect 158548 199668 158622 199696
rect 158686 199696 158714 200124
rect 158778 199918 158806 200124
rect 158766 199912 158818 199918
rect 158766 199854 158818 199860
rect 158870 199730 158898 200124
rect 158962 199918 158990 200124
rect 158950 199912 159002 199918
rect 159054 199889 159082 200124
rect 158950 199854 159002 199860
rect 159040 199880 159096 199889
rect 159040 199815 159096 199824
rect 158996 199776 159048 199782
rect 158870 199702 158944 199730
rect 159146 199764 159174 200124
rect 159238 199918 159266 200124
rect 159330 199918 159358 200124
rect 159226 199912 159278 199918
rect 159226 199854 159278 199860
rect 159318 199912 159370 199918
rect 159318 199854 159370 199860
rect 158996 199718 159048 199724
rect 159100 199736 159174 199764
rect 159272 199776 159324 199782
rect 158686 199668 158760 199696
rect 158088 195770 158116 199668
rect 158260 199640 158312 199646
rect 158260 199582 158312 199588
rect 158444 199640 158496 199646
rect 158444 199582 158496 199588
rect 158076 195764 158128 195770
rect 158076 195706 158128 195712
rect 157982 194032 158038 194041
rect 157982 193967 158038 193976
rect 158272 192302 158300 199582
rect 158260 192296 158312 192302
rect 158260 192238 158312 192244
rect 158456 191146 158484 199582
rect 158548 191185 158576 199668
rect 158628 199572 158680 199578
rect 158628 199514 158680 199520
rect 158534 191176 158590 191185
rect 158444 191140 158496 191146
rect 158534 191111 158590 191120
rect 158444 191082 158496 191088
rect 157904 190426 158208 190454
rect 157798 149560 157854 149569
rect 157798 149495 157854 149504
rect 158180 144498 158208 190426
rect 158640 151814 158668 199514
rect 158732 195362 158760 199668
rect 158812 199504 158864 199510
rect 158812 199446 158864 199452
rect 158720 195356 158772 195362
rect 158720 195298 158772 195304
rect 158824 190262 158852 199446
rect 158812 190256 158864 190262
rect 158812 190198 158864 190204
rect 158916 189281 158944 199702
rect 159008 198830 159036 199718
rect 158996 198824 159048 198830
rect 158996 198766 159048 198772
rect 158994 198520 159050 198529
rect 158994 198455 159050 198464
rect 159008 196790 159036 198455
rect 158996 196784 159048 196790
rect 158996 196726 159048 196732
rect 158996 191276 159048 191282
rect 158996 191218 159048 191224
rect 158902 189272 158958 189281
rect 158902 189207 158958 189216
rect 159008 152862 159036 191218
rect 159100 191049 159128 199736
rect 159272 199718 159324 199724
rect 159180 199640 159232 199646
rect 159180 199582 159232 199588
rect 159192 198898 159220 199582
rect 159180 198892 159232 198898
rect 159180 198834 159232 198840
rect 159086 191040 159142 191049
rect 159086 190975 159142 190984
rect 159284 184074 159312 199718
rect 159422 199696 159450 200124
rect 159514 199918 159542 200124
rect 159502 199912 159554 199918
rect 159502 199854 159554 199860
rect 159606 199764 159634 200124
rect 159698 199889 159726 200124
rect 159684 199880 159740 199889
rect 159684 199815 159740 199824
rect 159790 199764 159818 200124
rect 159882 199918 159910 200124
rect 159870 199912 159922 199918
rect 159870 199854 159922 199860
rect 159606 199736 159680 199764
rect 159376 199668 159450 199696
rect 159376 199481 159404 199668
rect 159548 199640 159600 199646
rect 159548 199582 159600 199588
rect 159362 199472 159418 199481
rect 159362 199407 159418 199416
rect 159364 199368 159416 199374
rect 159364 199310 159416 199316
rect 159376 184113 159404 199310
rect 159456 199096 159508 199102
rect 159456 199038 159508 199044
rect 159362 184104 159418 184113
rect 159272 184068 159324 184074
rect 159362 184039 159418 184048
rect 159272 184010 159324 184016
rect 159468 182174 159496 199038
rect 159560 196654 159588 199582
rect 159652 198966 159680 199736
rect 159744 199736 159818 199764
rect 159744 199238 159772 199736
rect 159974 199696 160002 200124
rect 160066 199764 160094 200124
rect 160158 199918 160186 200124
rect 160146 199912 160198 199918
rect 160146 199854 160198 199860
rect 160250 199764 160278 200124
rect 160342 199918 160370 200124
rect 160330 199912 160382 199918
rect 160330 199854 160382 199860
rect 160434 199764 160462 200124
rect 160526 199918 160554 200124
rect 160514 199912 160566 199918
rect 160514 199854 160566 199860
rect 160618 199764 160646 200124
rect 160710 199918 160738 200124
rect 160802 199918 160830 200124
rect 160698 199912 160750 199918
rect 160698 199854 160750 199860
rect 160790 199912 160842 199918
rect 160790 199854 160842 199860
rect 160894 199764 160922 200124
rect 160066 199753 160140 199764
rect 160066 199744 160154 199753
rect 160066 199736 160098 199744
rect 159974 199668 160048 199696
rect 160250 199736 160324 199764
rect 160388 199753 160462 199764
rect 160098 199679 160154 199688
rect 159824 199640 159876 199646
rect 159824 199582 159876 199588
rect 159732 199232 159784 199238
rect 159732 199174 159784 199180
rect 159836 199034 159864 199582
rect 159916 199504 159968 199510
rect 159916 199446 159968 199452
rect 159824 199028 159876 199034
rect 159824 198970 159876 198976
rect 159640 198960 159692 198966
rect 159640 198902 159692 198908
rect 159824 198416 159876 198422
rect 159824 198358 159876 198364
rect 159548 196648 159600 196654
rect 159548 196590 159600 196596
rect 159836 194594 159864 198358
rect 159652 194566 159864 194594
rect 159652 190454 159680 194566
rect 159928 191282 159956 199446
rect 160020 199102 160048 199668
rect 160192 199640 160244 199646
rect 160192 199582 160244 199588
rect 160008 199096 160060 199102
rect 160008 199038 160060 199044
rect 160008 198960 160060 198966
rect 160008 198902 160060 198908
rect 159916 191276 159968 191282
rect 159916 191218 159968 191224
rect 160020 191162 160048 198902
rect 160204 196194 160232 199582
rect 159928 191134 160048 191162
rect 160112 196166 160232 196194
rect 160112 191162 160140 196166
rect 160296 196058 160324 199736
rect 160374 199744 160462 199753
rect 160430 199736 160462 199744
rect 160572 199736 160646 199764
rect 160848 199736 160922 199764
rect 160374 199679 160430 199688
rect 160376 199640 160428 199646
rect 160376 199582 160428 199588
rect 160468 199640 160520 199646
rect 160468 199582 160520 199588
rect 160388 196926 160416 199582
rect 160376 196920 160428 196926
rect 160376 196862 160428 196868
rect 160204 196030 160324 196058
rect 160204 191321 160232 196030
rect 160282 195936 160338 195945
rect 160282 195871 160338 195880
rect 160190 191312 160246 191321
rect 160296 191298 160324 195871
rect 160480 191457 160508 199582
rect 160572 199306 160600 199736
rect 160744 199708 160796 199714
rect 160744 199650 160796 199656
rect 160652 199572 160704 199578
rect 160652 199514 160704 199520
rect 160560 199300 160612 199306
rect 160560 199242 160612 199248
rect 160664 194993 160692 199514
rect 160650 194984 160706 194993
rect 160650 194919 160706 194928
rect 160466 191448 160522 191457
rect 160466 191383 160522 191392
rect 160296 191270 160508 191298
rect 160190 191247 160246 191256
rect 160112 191134 160324 191162
rect 159652 190426 159864 190454
rect 159468 182146 159588 182174
rect 158996 152856 159048 152862
rect 158996 152798 159048 152804
rect 158548 151786 158668 151814
rect 158168 144492 158220 144498
rect 158168 144434 158220 144440
rect 158074 144120 158130 144129
rect 158074 144055 158130 144064
rect 157340 142248 157392 142254
rect 157340 142190 157392 142196
rect 157352 142089 157380 142190
rect 157338 142080 157394 142089
rect 157338 142015 157394 142024
rect 157154 141400 157210 141409
rect 157154 141335 157210 141344
rect 157062 140176 157118 140185
rect 157062 140111 157118 140120
rect 156124 139862 156460 139890
rect 156676 139862 157012 139890
rect 157168 139754 157196 141335
rect 158088 139890 158116 144055
rect 158548 140049 158576 151786
rect 159454 144256 159510 144265
rect 159454 144191 159510 144200
rect 158628 142860 158680 142866
rect 158628 142802 158680 142808
rect 158534 140040 158590 140049
rect 158534 139975 158590 139984
rect 158640 139890 158668 142802
rect 159180 142248 159232 142254
rect 159180 142190 159232 142196
rect 159192 139890 159220 142190
rect 159468 140162 159496 144191
rect 157780 139862 158116 139890
rect 158332 139862 158668 139890
rect 158884 139862 159220 139890
rect 159422 140134 159496 140162
rect 159422 139876 159450 140134
rect 157168 139726 157228 139754
rect 159560 139369 159588 182146
rect 159836 139369 159864 190426
rect 159928 145722 159956 191134
rect 160192 191072 160244 191078
rect 160192 191014 160244 191020
rect 160100 191004 160152 191010
rect 160100 190946 160152 190952
rect 160008 184068 160060 184074
rect 160008 184010 160060 184016
rect 160020 152726 160048 184010
rect 160008 152720 160060 152726
rect 160008 152662 160060 152668
rect 160112 145790 160140 190946
rect 160204 148646 160232 191014
rect 160296 153066 160324 191134
rect 160376 191140 160428 191146
rect 160376 191082 160428 191088
rect 160284 153060 160336 153066
rect 160284 153002 160336 153008
rect 160388 152794 160416 191082
rect 160480 152930 160508 191270
rect 160756 191185 160784 199650
rect 160848 197062 160876 199736
rect 160986 199730 161014 200124
rect 161078 199889 161106 200124
rect 161170 199918 161198 200124
rect 161158 199912 161210 199918
rect 161064 199880 161120 199889
rect 161158 199854 161210 199860
rect 161064 199815 161120 199824
rect 160986 199702 161060 199730
rect 160928 199640 160980 199646
rect 160928 199582 160980 199588
rect 160836 197056 160888 197062
rect 160836 196998 160888 197004
rect 160742 191176 160798 191185
rect 160742 191111 160798 191120
rect 160940 191078 160968 199582
rect 160928 191072 160980 191078
rect 160928 191014 160980 191020
rect 161032 191010 161060 199702
rect 161262 199696 161290 200124
rect 161354 199764 161382 200124
rect 161446 199918 161474 200124
rect 161434 199912 161486 199918
rect 161434 199854 161486 199860
rect 161538 199764 161566 200124
rect 161354 199736 161428 199764
rect 161262 199668 161336 199696
rect 161202 199472 161258 199481
rect 161202 199407 161204 199416
rect 161256 199407 161258 199416
rect 161204 199378 161256 199384
rect 161308 191146 161336 199668
rect 161296 191140 161348 191146
rect 161296 191082 161348 191088
rect 161400 191049 161428 199736
rect 161492 199736 161566 199764
rect 161630 199764 161658 200124
rect 161722 199918 161750 200124
rect 161710 199912 161762 199918
rect 161710 199854 161762 199860
rect 161814 199764 161842 200124
rect 161906 199918 161934 200124
rect 161894 199912 161946 199918
rect 161894 199854 161946 199860
rect 161998 199764 162026 200124
rect 162090 199782 162118 200124
rect 162182 199918 162210 200124
rect 162274 199918 162302 200124
rect 162366 199918 162394 200124
rect 162458 199918 162486 200124
rect 162170 199912 162222 199918
rect 162170 199854 162222 199860
rect 162262 199912 162314 199918
rect 162262 199854 162314 199860
rect 162354 199912 162406 199918
rect 162354 199854 162406 199860
rect 162446 199912 162498 199918
rect 162446 199854 162498 199860
rect 161630 199736 161704 199764
rect 161814 199736 161888 199764
rect 161492 194274 161520 199736
rect 161572 199640 161624 199646
rect 161572 199582 161624 199588
rect 161584 195634 161612 199582
rect 161676 199578 161704 199736
rect 161664 199572 161716 199578
rect 161664 199514 161716 199520
rect 161860 199424 161888 199736
rect 161676 199396 161888 199424
rect 161952 199736 162026 199764
rect 162078 199776 162130 199782
rect 161572 195628 161624 195634
rect 161572 195570 161624 195576
rect 161676 195276 161704 199396
rect 161848 199300 161900 199306
rect 161848 199242 161900 199248
rect 161860 195294 161888 199242
rect 161584 195248 161704 195276
rect 161848 195288 161900 195294
rect 161480 194268 161532 194274
rect 161480 194210 161532 194216
rect 161386 191040 161442 191049
rect 161020 191004 161072 191010
rect 161386 190975 161442 190984
rect 161020 190946 161072 190952
rect 161480 185156 161532 185162
rect 161480 185098 161532 185104
rect 160468 152924 160520 152930
rect 160468 152866 160520 152872
rect 160376 152788 160428 152794
rect 160376 152730 160428 152736
rect 160192 148640 160244 148646
rect 160192 148582 160244 148588
rect 161492 145926 161520 185098
rect 161584 146062 161612 195248
rect 161848 195230 161900 195236
rect 161846 195120 161902 195129
rect 161846 195055 161902 195064
rect 161756 194268 161808 194274
rect 161756 194210 161808 194216
rect 161664 191140 161716 191146
rect 161664 191082 161716 191088
rect 161572 146056 161624 146062
rect 161572 145998 161624 146004
rect 161480 145920 161532 145926
rect 161480 145862 161532 145868
rect 160100 145784 160152 145790
rect 160100 145726 160152 145732
rect 160650 145752 160706 145761
rect 159916 145716 159968 145722
rect 160650 145687 160706 145696
rect 159916 145658 159968 145664
rect 160100 145648 160152 145654
rect 160100 145590 160152 145596
rect 160006 143032 160062 143041
rect 160006 142967 160062 142976
rect 160020 140162 160048 142967
rect 159974 140134 160048 140162
rect 159974 139876 160002 140134
rect 160112 139890 160140 145590
rect 160664 139890 160692 145687
rect 161676 145654 161704 191082
rect 161768 153134 161796 194210
rect 161860 193934 161888 195055
rect 161848 193928 161900 193934
rect 161848 193870 161900 193876
rect 161952 187105 161980 199736
rect 162078 199718 162130 199724
rect 162308 199776 162360 199782
rect 162550 199730 162578 200124
rect 162642 199918 162670 200124
rect 162630 199912 162682 199918
rect 162630 199854 162682 199860
rect 162734 199764 162762 200124
rect 162308 199718 162360 199724
rect 162320 199594 162348 199718
rect 162504 199702 162578 199730
rect 162688 199736 162762 199764
rect 162504 199696 162532 199702
rect 162032 199572 162084 199578
rect 162032 199514 162084 199520
rect 162136 199566 162348 199594
rect 162412 199668 162532 199696
rect 161938 187096 161994 187105
rect 161938 187031 161994 187040
rect 162044 180794 162072 199514
rect 162136 185162 162164 199566
rect 162216 199504 162268 199510
rect 162216 199446 162268 199452
rect 162228 195498 162256 199446
rect 162412 199170 162440 199668
rect 162584 199640 162636 199646
rect 162584 199582 162636 199588
rect 162492 199572 162544 199578
rect 162492 199514 162544 199520
rect 162400 199164 162452 199170
rect 162400 199106 162452 199112
rect 162306 198384 162362 198393
rect 162306 198319 162362 198328
rect 162320 196518 162348 198319
rect 162308 196512 162360 196518
rect 162308 196454 162360 196460
rect 162216 195492 162268 195498
rect 162216 195434 162268 195440
rect 162504 187513 162532 199514
rect 162596 191146 162624 199582
rect 162688 191185 162716 199736
rect 162826 199696 162854 200124
rect 162780 199668 162854 199696
rect 162780 199510 162808 199668
rect 162918 199628 162946 200124
rect 163010 199764 163038 200124
rect 163102 199889 163130 200124
rect 163088 199880 163144 199889
rect 163088 199815 163144 199824
rect 163194 199764 163222 200124
rect 163010 199753 163084 199764
rect 163010 199744 163098 199753
rect 163010 199736 163042 199744
rect 163042 199679 163098 199688
rect 163148 199736 163222 199764
rect 163286 199753 163314 200124
rect 163272 199744 163328 199753
rect 162872 199600 162946 199628
rect 163044 199640 163096 199646
rect 162768 199504 162820 199510
rect 162768 199446 162820 199452
rect 162768 199368 162820 199374
rect 162768 199310 162820 199316
rect 162780 198898 162808 199310
rect 162768 198892 162820 198898
rect 162768 198834 162820 198840
rect 162674 191176 162730 191185
rect 162584 191140 162636 191146
rect 162674 191111 162730 191120
rect 162584 191082 162636 191088
rect 162872 189718 162900 199600
rect 163044 199582 163096 199588
rect 162950 199472 163006 199481
rect 162950 199407 163006 199416
rect 162964 195401 162992 199407
rect 163056 195945 163084 199582
rect 163042 195936 163098 195945
rect 163042 195871 163098 195880
rect 162950 195392 163006 195401
rect 162950 195327 163006 195336
rect 163148 195242 163176 199736
rect 163272 199679 163328 199688
rect 163378 199628 163406 200124
rect 163332 199600 163406 199628
rect 163226 199472 163282 199481
rect 163226 199407 163282 199416
rect 162964 195214 163176 195242
rect 162860 189712 162912 189718
rect 162860 189654 162912 189660
rect 162860 189372 162912 189378
rect 162860 189314 162912 189320
rect 162490 187504 162546 187513
rect 162490 187439 162546 187448
rect 162124 185156 162176 185162
rect 162124 185098 162176 185104
rect 161860 180766 162072 180794
rect 161756 153128 161808 153134
rect 161756 153070 161808 153076
rect 161860 152998 161888 180766
rect 161848 152992 161900 152998
rect 161848 152934 161900 152940
rect 162306 145888 162362 145897
rect 162306 145823 162362 145832
rect 161664 145648 161716 145654
rect 161664 145590 161716 145596
rect 162214 144528 162270 144537
rect 162214 144463 162270 144472
rect 161938 143168 161994 143177
rect 161938 143103 161994 143112
rect 161480 142248 161532 142254
rect 161480 142190 161532 142196
rect 161492 142118 161520 142190
rect 161480 142112 161532 142118
rect 161480 142054 161532 142060
rect 161952 139890 161980 143103
rect 162228 140162 162256 144463
rect 160112 139862 160540 139890
rect 160664 139862 161092 139890
rect 161644 139862 161980 139890
rect 162182 140134 162256 140162
rect 162182 139876 162210 140134
rect 162320 139890 162348 145823
rect 162872 141438 162900 189314
rect 162964 145858 162992 195214
rect 163044 192840 163096 192846
rect 163044 192782 163096 192788
rect 163056 148510 163084 192782
rect 163240 190482 163268 199407
rect 163332 197946 163360 199600
rect 163470 199560 163498 200124
rect 163562 199628 163590 200124
rect 163654 199764 163682 200124
rect 163746 199889 163774 200124
rect 163732 199880 163788 199889
rect 163732 199815 163788 199824
rect 163654 199736 163728 199764
rect 163562 199600 163636 199628
rect 163424 199532 163498 199560
rect 163320 197940 163372 197946
rect 163320 197882 163372 197888
rect 163424 192846 163452 199532
rect 163608 198257 163636 199600
rect 163594 198248 163650 198257
rect 163594 198183 163650 198192
rect 163504 197940 163556 197946
rect 163504 197882 163556 197888
rect 163516 197130 163544 197882
rect 163504 197124 163556 197130
rect 163504 197066 163556 197072
rect 163700 196994 163728 199736
rect 163838 199730 163866 200124
rect 163930 199918 163958 200124
rect 163918 199912 163970 199918
rect 164022 199889 164050 200124
rect 163918 199854 163970 199860
rect 164008 199880 164064 199889
rect 164008 199815 164064 199824
rect 164114 199764 164142 200124
rect 163962 199744 164018 199753
rect 163838 199702 163912 199730
rect 163780 199640 163832 199646
rect 163780 199582 163832 199588
rect 163792 197742 163820 199582
rect 163780 197736 163832 197742
rect 163780 197678 163832 197684
rect 163688 196988 163740 196994
rect 163688 196930 163740 196936
rect 163412 192840 163464 192846
rect 163412 192782 163464 192788
rect 163148 190454 163268 190482
rect 163148 153202 163176 190454
rect 163228 189712 163280 189718
rect 163228 189654 163280 189660
rect 163136 153196 163188 153202
rect 163136 153138 163188 153144
rect 163240 152454 163268 189654
rect 163884 187377 163912 199702
rect 163962 199679 164018 199688
rect 164068 199736 164142 199764
rect 163976 189378 164004 199679
rect 164068 195265 164096 199736
rect 164206 199594 164234 200124
rect 164298 199628 164326 200124
rect 164390 199889 164418 200124
rect 164376 199880 164432 199889
rect 164376 199815 164432 199824
rect 164482 199764 164510 200124
rect 164574 199918 164602 200124
rect 164666 199918 164694 200124
rect 164758 199918 164786 200124
rect 164562 199912 164614 199918
rect 164562 199854 164614 199860
rect 164654 199912 164706 199918
rect 164654 199854 164706 199860
rect 164746 199912 164798 199918
rect 164850 199889 164878 200124
rect 164942 199918 164970 200124
rect 165034 199918 165062 200124
rect 165126 199918 165154 200124
rect 164930 199912 164982 199918
rect 164746 199854 164798 199860
rect 164836 199880 164892 199889
rect 164930 199854 164982 199860
rect 165022 199912 165074 199918
rect 165022 199854 165074 199860
rect 165114 199912 165166 199918
rect 165218 199889 165246 200124
rect 165310 199918 165338 200124
rect 165402 199918 165430 200124
rect 165494 199918 165522 200124
rect 165586 199918 165614 200124
rect 165678 199918 165706 200124
rect 165770 199918 165798 200124
rect 165862 199923 165890 200124
rect 165298 199912 165350 199918
rect 165114 199854 165166 199860
rect 165204 199880 165260 199889
rect 164836 199815 164892 199824
rect 165298 199854 165350 199860
rect 165390 199912 165442 199918
rect 165390 199854 165442 199860
rect 165482 199912 165534 199918
rect 165482 199854 165534 199860
rect 165574 199912 165626 199918
rect 165574 199854 165626 199860
rect 165666 199912 165718 199918
rect 165666 199854 165718 199860
rect 165758 199912 165810 199918
rect 165758 199854 165810 199860
rect 165848 199914 165904 199923
rect 165848 199849 165904 199858
rect 165204 199815 165260 199824
rect 164436 199736 164510 199764
rect 165436 199776 165488 199782
rect 164298 199600 164372 199628
rect 164160 199566 164234 199594
rect 164160 197266 164188 199566
rect 164240 199504 164292 199510
rect 164240 199446 164292 199452
rect 164148 197260 164200 197266
rect 164148 197202 164200 197208
rect 164054 195256 164110 195265
rect 164054 195191 164110 195200
rect 164252 192778 164280 199446
rect 164240 192772 164292 192778
rect 164240 192714 164292 192720
rect 164344 191282 164372 199600
rect 164436 197198 164464 199736
rect 165436 199718 165488 199724
rect 165618 199744 165674 199753
rect 164792 199708 164844 199714
rect 164792 199650 164844 199656
rect 164976 199708 165028 199714
rect 164976 199650 165028 199656
rect 165068 199708 165120 199714
rect 165068 199650 165120 199656
rect 165344 199708 165396 199714
rect 165344 199650 165396 199656
rect 164516 199640 164568 199646
rect 164516 199582 164568 199588
rect 164700 199640 164752 199646
rect 164700 199582 164752 199588
rect 164424 197192 164476 197198
rect 164424 197134 164476 197140
rect 164528 195242 164556 199582
rect 164712 195265 164740 199582
rect 164804 197334 164832 199650
rect 164884 199300 164936 199306
rect 164884 199242 164936 199248
rect 164896 199102 164924 199242
rect 164884 199096 164936 199102
rect 164884 199038 164936 199044
rect 164792 197328 164844 197334
rect 164792 197270 164844 197276
rect 164988 196625 165016 199650
rect 164974 196616 165030 196625
rect 164974 196551 165030 196560
rect 164436 195214 164556 195242
rect 164698 195256 164754 195265
rect 164332 191276 164384 191282
rect 164332 191218 164384 191224
rect 163964 189372 164016 189378
rect 163964 189314 164016 189320
rect 163870 187368 163926 187377
rect 163870 187303 163926 187312
rect 164332 183388 164384 183394
rect 164332 183330 164384 183336
rect 163228 152448 163280 152454
rect 163228 152390 163280 152396
rect 163044 148504 163096 148510
rect 163044 148446 163096 148452
rect 162952 145852 163004 145858
rect 162952 145794 163004 145800
rect 163594 143304 163650 143313
rect 163594 143239 163650 143248
rect 162860 141432 162912 141438
rect 162860 141374 162912 141380
rect 163608 139890 163636 143239
rect 164146 141536 164202 141545
rect 164344 141506 164372 183330
rect 164436 148714 164464 195214
rect 164698 195191 164754 195200
rect 164976 195220 165028 195226
rect 164976 195162 165028 195168
rect 164514 194984 164570 194993
rect 164514 194919 164570 194928
rect 164424 148708 164476 148714
rect 164424 148650 164476 148656
rect 164528 148442 164556 194919
rect 164608 191276 164660 191282
rect 164608 191218 164660 191224
rect 164620 152590 164648 191218
rect 164988 188601 165016 195162
rect 165080 190454 165108 199650
rect 165160 199640 165212 199646
rect 165160 199582 165212 199588
rect 165172 195226 165200 199582
rect 165252 199436 165304 199442
rect 165252 199378 165304 199384
rect 165160 195220 165212 195226
rect 165160 195162 165212 195168
rect 165080 190426 165200 190454
rect 164974 188592 165030 188601
rect 164974 188527 165030 188536
rect 164608 152584 164660 152590
rect 164608 152526 164660 152532
rect 165172 151814 165200 190426
rect 165264 182617 165292 199378
rect 165356 183394 165384 199650
rect 165448 185881 165476 199718
rect 165528 199708 165580 199714
rect 165954 199730 165982 200124
rect 166046 199850 166074 200124
rect 166034 199844 166086 199850
rect 166034 199786 166086 199792
rect 165618 199679 165674 199688
rect 165712 199708 165764 199714
rect 165528 199650 165580 199656
rect 165540 193050 165568 199650
rect 165632 199442 165660 199679
rect 165712 199650 165764 199656
rect 165908 199702 165982 199730
rect 165620 199436 165672 199442
rect 165620 199378 165672 199384
rect 165724 199288 165752 199650
rect 165632 199260 165752 199288
rect 165632 197606 165660 199260
rect 165712 199164 165764 199170
rect 165712 199106 165764 199112
rect 165620 197600 165672 197606
rect 165620 197542 165672 197548
rect 165620 196240 165672 196246
rect 165620 196182 165672 196188
rect 165528 193044 165580 193050
rect 165528 192986 165580 192992
rect 165434 185872 165490 185881
rect 165434 185807 165490 185816
rect 165344 183388 165396 183394
rect 165344 183330 165396 183336
rect 165250 182608 165306 182617
rect 165250 182543 165306 182552
rect 165172 151786 165384 151814
rect 164516 148436 164568 148442
rect 164516 148378 164568 148384
rect 164422 146024 164478 146033
rect 164422 145959 164478 145968
rect 164146 141471 164202 141480
rect 164332 141500 164384 141506
rect 164160 139890 164188 141471
rect 164332 141442 164384 141448
rect 164436 140162 164464 145959
rect 165250 143440 165306 143449
rect 165250 143375 165306 143384
rect 162320 139862 162748 139890
rect 163300 139862 163636 139890
rect 163852 139862 164188 139890
rect 164390 140134 164464 140162
rect 164390 139876 164418 140134
rect 165264 139890 165292 143375
rect 164956 139862 165292 139890
rect 165356 139369 165384 151786
rect 165632 145994 165660 196182
rect 165724 195702 165752 199106
rect 165712 195696 165764 195702
rect 165712 195638 165764 195644
rect 165908 194594 165936 199702
rect 165988 199640 166040 199646
rect 166138 199594 166166 200124
rect 166230 199918 166258 200124
rect 166218 199912 166270 199918
rect 166218 199854 166270 199860
rect 166322 199850 166350 200124
rect 166414 199923 166442 200124
rect 166400 199914 166456 199923
rect 166310 199844 166362 199850
rect 166400 199849 166456 199858
rect 166310 199786 166362 199792
rect 166506 199764 166534 200124
rect 166354 199744 166410 199753
rect 166354 199679 166410 199688
rect 166460 199736 166534 199764
rect 165988 199582 166040 199588
rect 165724 194566 165936 194594
rect 165724 152522 165752 194566
rect 165804 192296 165856 192302
rect 165804 192238 165856 192244
rect 165712 152516 165764 152522
rect 165712 152458 165764 152464
rect 165816 152386 165844 192238
rect 166000 190097 166028 199582
rect 166092 199566 166166 199594
rect 166092 194410 166120 199566
rect 166172 199504 166224 199510
rect 166172 199446 166224 199452
rect 166184 196246 166212 199446
rect 166368 199034 166396 199679
rect 166356 199028 166408 199034
rect 166356 198970 166408 198976
rect 166172 196240 166224 196246
rect 166172 196182 166224 196188
rect 166264 195832 166316 195838
rect 166264 195774 166316 195780
rect 166276 195566 166304 195774
rect 166264 195560 166316 195566
rect 166264 195502 166316 195508
rect 166460 194594 166488 199736
rect 166598 199696 166626 200124
rect 166690 199923 166718 200124
rect 166676 199914 166732 199923
rect 166782 199918 166810 200124
rect 166874 199918 166902 200124
rect 166676 199849 166732 199858
rect 166770 199912 166822 199918
rect 166770 199854 166822 199860
rect 166862 199912 166914 199918
rect 166966 199889 166994 200124
rect 167058 199918 167086 200124
rect 167150 199918 167178 200124
rect 167242 199918 167270 200124
rect 167046 199912 167098 199918
rect 166862 199854 166914 199860
rect 166952 199880 167008 199889
rect 167046 199854 167098 199860
rect 167138 199912 167190 199918
rect 167138 199854 167190 199860
rect 167230 199912 167282 199918
rect 167230 199854 167282 199860
rect 166952 199815 167008 199824
rect 166724 199776 166776 199782
rect 166908 199776 166960 199782
rect 166724 199718 166776 199724
rect 166814 199744 166870 199753
rect 166552 199668 166626 199696
rect 166552 197305 166580 199668
rect 166538 197296 166594 197305
rect 166538 197231 166594 197240
rect 166460 194566 166580 194594
rect 166080 194404 166132 194410
rect 166080 194346 166132 194352
rect 166552 190454 166580 194566
rect 166736 192302 166764 199718
rect 167334 199764 167362 200124
rect 167426 199918 167454 200124
rect 167414 199912 167466 199918
rect 167414 199854 167466 199860
rect 167518 199764 167546 200124
rect 166908 199718 166960 199724
rect 167090 199744 167146 199753
rect 166814 199679 166816 199688
rect 166868 199679 166870 199688
rect 166816 199650 166868 199656
rect 166816 199572 166868 199578
rect 166816 199514 166868 199520
rect 166828 192506 166856 199514
rect 166816 192500 166868 192506
rect 166816 192442 166868 192448
rect 166724 192296 166776 192302
rect 166724 192238 166776 192244
rect 166920 191185 166948 199718
rect 167288 199736 167362 199764
rect 167472 199736 167546 199764
rect 167090 199679 167146 199688
rect 167184 199708 167236 199714
rect 167000 199572 167052 199578
rect 167000 199514 167052 199520
rect 167012 194682 167040 199514
rect 167104 198626 167132 199679
rect 167184 199650 167236 199656
rect 167092 198620 167144 198626
rect 167092 198562 167144 198568
rect 167090 198112 167146 198121
rect 167090 198047 167146 198056
rect 167104 197713 167132 198047
rect 167090 197704 167146 197713
rect 167090 197639 167146 197648
rect 167000 194676 167052 194682
rect 167000 194618 167052 194624
rect 167000 194540 167052 194546
rect 167000 194482 167052 194488
rect 166906 191176 166962 191185
rect 166906 191111 166962 191120
rect 166460 190426 166580 190454
rect 165986 190088 166042 190097
rect 165986 190023 166042 190032
rect 166460 180794 166488 190426
rect 165908 180766 166488 180794
rect 165908 152561 165936 180766
rect 165894 152552 165950 152561
rect 165894 152487 165950 152496
rect 165804 152380 165856 152386
rect 165804 152322 165856 152328
rect 167012 148578 167040 194482
rect 167196 194070 167224 199650
rect 167184 194064 167236 194070
rect 167184 194006 167236 194012
rect 167288 192914 167316 199736
rect 167368 199640 167420 199646
rect 167368 199582 167420 199588
rect 167380 195537 167408 199582
rect 167472 198898 167500 199736
rect 167610 199696 167638 200124
rect 167564 199668 167638 199696
rect 167460 198892 167512 198898
rect 167460 198834 167512 198840
rect 167366 195528 167422 195537
rect 167366 195463 167422 195472
rect 167276 192908 167328 192914
rect 167276 192850 167328 192856
rect 167092 191276 167144 191282
rect 167092 191218 167144 191224
rect 167104 152658 167132 191218
rect 167564 176654 167592 199668
rect 167702 199628 167730 200124
rect 167794 199764 167822 200124
rect 167886 199918 167914 200124
rect 167978 199918 168006 200124
rect 168070 199918 168098 200124
rect 167874 199912 167926 199918
rect 167874 199854 167926 199860
rect 167966 199912 168018 199918
rect 167966 199854 168018 199860
rect 168058 199912 168110 199918
rect 168058 199854 168110 199860
rect 167920 199776 167972 199782
rect 167794 199736 167868 199764
rect 167656 199600 167730 199628
rect 167656 198665 167684 199600
rect 167736 199368 167788 199374
rect 167736 199310 167788 199316
rect 167748 198830 167776 199310
rect 167840 198830 167868 199736
rect 168162 199764 168190 200124
rect 168254 199889 168282 200124
rect 168240 199880 168296 199889
rect 168240 199815 168296 199824
rect 167920 199718 167972 199724
rect 168116 199736 168190 199764
rect 167736 198824 167788 198830
rect 167736 198766 167788 198772
rect 167828 198824 167880 198830
rect 167828 198766 167880 198772
rect 167642 198656 167698 198665
rect 167642 198591 167698 198600
rect 167932 195401 167960 199718
rect 168012 199708 168064 199714
rect 168012 199650 168064 199656
rect 167918 195392 167974 195401
rect 167918 195327 167974 195336
rect 168024 194274 168052 199650
rect 168012 194268 168064 194274
rect 168012 194210 168064 194216
rect 168116 191282 168144 199736
rect 168346 199696 168374 200124
rect 168438 199918 168466 200124
rect 168426 199912 168478 199918
rect 168426 199854 168478 199860
rect 168530 199764 168558 200124
rect 168622 199889 168650 200124
rect 168608 199880 168664 199889
rect 168608 199815 168664 199824
rect 168530 199736 168604 199764
rect 168346 199668 168420 199696
rect 168392 199050 168420 199668
rect 168472 199640 168524 199646
rect 168472 199582 168524 199588
rect 168208 199022 168420 199050
rect 168208 192642 168236 199022
rect 168378 195528 168434 195537
rect 168378 195463 168434 195472
rect 168288 192908 168340 192914
rect 168288 192850 168340 192856
rect 168196 192636 168248 192642
rect 168196 192578 168248 192584
rect 168104 191276 168156 191282
rect 168104 191218 168156 191224
rect 167288 176626 167592 176654
rect 167288 155242 167316 176626
rect 167276 155236 167328 155242
rect 167276 155178 167328 155184
rect 167092 152652 167144 152658
rect 167092 152594 167144 152600
rect 168300 152425 168328 192850
rect 168286 152416 168342 152425
rect 168286 152351 168342 152360
rect 168392 152318 168420 195463
rect 168484 154465 168512 199582
rect 168576 194206 168604 199736
rect 168714 199730 168742 200124
rect 168806 199918 168834 200124
rect 168898 199918 168926 200124
rect 168990 199918 169018 200124
rect 169082 199923 169110 200124
rect 168794 199912 168846 199918
rect 168794 199854 168846 199860
rect 168886 199912 168938 199918
rect 168886 199854 168938 199860
rect 168978 199912 169030 199918
rect 168978 199854 169030 199860
rect 169068 199914 169124 199923
rect 169068 199849 169124 199858
rect 169174 199730 169202 200124
rect 169266 199918 169294 200124
rect 169254 199912 169306 199918
rect 169254 199854 169306 199860
rect 169358 199764 169386 200124
rect 168714 199702 168788 199730
rect 168656 199504 168708 199510
rect 168656 199446 168708 199452
rect 168668 194546 168696 199446
rect 168760 195401 168788 199702
rect 168840 199708 168892 199714
rect 168840 199650 168892 199656
rect 168932 199708 168984 199714
rect 168932 199650 168984 199656
rect 169128 199702 169202 199730
rect 169312 199736 169386 199764
rect 169450 199764 169478 200124
rect 169542 199889 169570 200124
rect 169634 199918 169662 200124
rect 169726 199918 169754 200124
rect 169818 199918 169846 200124
rect 169910 199918 169938 200124
rect 169622 199912 169674 199918
rect 169528 199880 169584 199889
rect 169622 199854 169674 199860
rect 169714 199912 169766 199918
rect 169714 199854 169766 199860
rect 169806 199912 169858 199918
rect 169806 199854 169858 199860
rect 169898 199912 169950 199918
rect 170002 199889 170030 200124
rect 170094 199918 170122 200124
rect 170186 199918 170214 200124
rect 170082 199912 170134 199918
rect 169898 199854 169950 199860
rect 169988 199880 170044 199889
rect 169528 199815 169584 199824
rect 170082 199854 170134 199860
rect 170174 199912 170226 199918
rect 170174 199854 170226 199860
rect 169988 199815 170044 199824
rect 170036 199776 170088 199782
rect 169450 199736 169524 199764
rect 168746 195392 168802 195401
rect 168746 195327 168802 195336
rect 168748 195152 168800 195158
rect 168748 195094 168800 195100
rect 168656 194540 168708 194546
rect 168656 194482 168708 194488
rect 168564 194200 168616 194206
rect 168564 194142 168616 194148
rect 168760 185881 168788 195094
rect 168852 190454 168880 199650
rect 168944 198812 168972 199650
rect 168944 198784 169064 198812
rect 169036 195226 169064 198784
rect 169024 195220 169076 195226
rect 169024 195162 169076 195168
rect 169128 194138 169156 199702
rect 169208 199572 169260 199578
rect 169208 199514 169260 199520
rect 169220 195158 169248 199514
rect 169208 195152 169260 195158
rect 169208 195094 169260 195100
rect 169116 194132 169168 194138
rect 169116 194074 169168 194080
rect 169312 191185 169340 199736
rect 169392 199640 169444 199646
rect 169392 199582 169444 199588
rect 169404 199238 169432 199582
rect 169392 199232 169444 199238
rect 169392 199174 169444 199180
rect 169392 199096 169444 199102
rect 169392 199038 169444 199044
rect 169404 198966 169432 199038
rect 169392 198960 169444 198966
rect 169392 198902 169444 198908
rect 169496 192710 169524 199736
rect 170278 199764 170306 200124
rect 170036 199718 170088 199724
rect 170232 199736 170306 199764
rect 169576 199708 169628 199714
rect 169576 199650 169628 199656
rect 169668 199708 169720 199714
rect 169668 199650 169720 199656
rect 169852 199708 169904 199714
rect 169852 199650 169904 199656
rect 169588 199578 169616 199650
rect 169576 199572 169628 199578
rect 169576 199514 169628 199520
rect 169574 199472 169630 199481
rect 169574 199407 169630 199416
rect 169588 196761 169616 199407
rect 169680 198529 169708 199650
rect 169760 199504 169812 199510
rect 169758 199472 169760 199481
rect 169812 199472 169814 199481
rect 169758 199407 169814 199416
rect 169760 199368 169812 199374
rect 169760 199310 169812 199316
rect 169666 198520 169722 198529
rect 169666 198455 169722 198464
rect 169772 198121 169800 199310
rect 169758 198112 169814 198121
rect 169758 198047 169814 198056
rect 169760 198008 169812 198014
rect 169760 197950 169812 197956
rect 169574 196752 169630 196761
rect 169574 196687 169630 196696
rect 169772 195838 169800 197950
rect 169864 197033 169892 199650
rect 169944 199096 169996 199102
rect 169944 199038 169996 199044
rect 169956 198354 169984 199038
rect 169944 198348 169996 198354
rect 169944 198290 169996 198296
rect 169850 197024 169906 197033
rect 169850 196959 169906 196968
rect 169760 195832 169812 195838
rect 169760 195774 169812 195780
rect 169576 195220 169628 195226
rect 169576 195162 169628 195168
rect 169484 192704 169536 192710
rect 169484 192646 169536 192652
rect 169298 191176 169354 191185
rect 169298 191111 169354 191120
rect 168852 190426 168972 190454
rect 168746 185872 168802 185881
rect 168746 185807 168802 185816
rect 168944 182174 168972 190426
rect 168944 182146 169248 182174
rect 169220 176654 169248 182146
rect 168668 176626 169248 176654
rect 168668 155378 168696 176626
rect 168656 155372 168708 155378
rect 168656 155314 168708 155320
rect 169588 155310 169616 195162
rect 170048 191162 170076 199718
rect 170128 199640 170180 199646
rect 170128 199582 170180 199588
rect 170140 199481 170168 199582
rect 170126 199472 170182 199481
rect 170126 199407 170182 199416
rect 170128 198824 170180 198830
rect 170128 198766 170180 198772
rect 170140 192982 170168 198766
rect 170232 197810 170260 199736
rect 170370 199628 170398 200124
rect 170462 199889 170490 200124
rect 170554 199918 170582 200124
rect 170646 199918 170674 200124
rect 170738 199918 170766 200124
rect 170830 199918 170858 200124
rect 170542 199912 170594 199918
rect 170448 199880 170504 199889
rect 170542 199854 170594 199860
rect 170634 199912 170686 199918
rect 170634 199854 170686 199860
rect 170726 199912 170778 199918
rect 170726 199854 170778 199860
rect 170818 199912 170870 199918
rect 170818 199854 170870 199860
rect 170448 199815 170504 199824
rect 170496 199776 170548 199782
rect 170922 199764 170950 200124
rect 171014 199889 171042 200124
rect 171106 199918 171134 200124
rect 171094 199912 171146 199918
rect 171000 199880 171056 199889
rect 171094 199854 171146 199860
rect 171000 199815 171056 199824
rect 171048 199776 171100 199782
rect 170770 199744 170826 199753
rect 170496 199718 170548 199724
rect 170324 199600 170398 199628
rect 170220 197804 170272 197810
rect 170220 197746 170272 197752
rect 170128 192976 170180 192982
rect 170128 192918 170180 192924
rect 169864 191134 170076 191162
rect 169760 189032 169812 189038
rect 169760 188974 169812 188980
rect 169576 155304 169628 155310
rect 169576 155246 169628 155252
rect 168470 154456 168526 154465
rect 168470 154391 168526 154400
rect 168380 152312 168432 152318
rect 168380 152254 168432 152260
rect 167000 148572 167052 148578
rect 167000 148514 167052 148520
rect 165620 145988 165672 145994
rect 165620 145930 165672 145936
rect 168010 144800 168066 144809
rect 168010 144735 168066 144744
rect 166354 144664 166410 144673
rect 166354 144599 166410 144608
rect 165526 143984 165582 143993
rect 165526 143919 165582 143928
rect 165540 140162 165568 143919
rect 165494 140134 165568 140162
rect 165494 139876 165522 140134
rect 166368 139890 166396 144599
rect 166908 142928 166960 142934
rect 166908 142870 166960 142876
rect 166920 139890 166948 142870
rect 167460 141568 167512 141574
rect 167460 141510 167512 141516
rect 167472 139890 167500 141510
rect 168024 139890 168052 144735
rect 169116 144560 169168 144566
rect 169116 144502 169168 144508
rect 168288 142996 168340 143002
rect 168288 142938 168340 142944
rect 168300 140162 168328 142938
rect 166060 139862 166396 139890
rect 166612 139862 166948 139890
rect 167164 139862 167500 139890
rect 167716 139862 168052 139890
rect 168254 140134 168328 140162
rect 168254 139876 168282 140134
rect 169128 139890 169156 144502
rect 169668 143200 169720 143206
rect 169668 143142 169720 143148
rect 169680 139890 169708 143142
rect 169772 140457 169800 188974
rect 169758 140448 169814 140457
rect 169758 140383 169814 140392
rect 169864 140146 169892 191134
rect 169944 188692 169996 188698
rect 169944 188634 169996 188640
rect 169956 140321 169984 188634
rect 170324 176654 170352 199600
rect 170402 199472 170458 199481
rect 170402 199407 170458 199416
rect 170416 189281 170444 199407
rect 170508 197878 170536 199718
rect 170588 199708 170640 199714
rect 170588 199650 170640 199656
rect 170692 199702 170770 199730
rect 170496 197872 170548 197878
rect 170496 197814 170548 197820
rect 170402 189272 170458 189281
rect 170402 189207 170458 189216
rect 170600 188698 170628 199650
rect 170692 199322 170720 199702
rect 170922 199736 170996 199764
rect 170770 199679 170826 199688
rect 170864 199572 170916 199578
rect 170864 199514 170916 199520
rect 170772 199504 170824 199510
rect 170770 199472 170772 199481
rect 170824 199472 170826 199481
rect 170770 199407 170826 199416
rect 170692 199294 170812 199322
rect 170784 199102 170812 199294
rect 170772 199096 170824 199102
rect 170772 199038 170824 199044
rect 170772 198960 170824 198966
rect 170772 198902 170824 198908
rect 170784 198762 170812 198902
rect 170772 198756 170824 198762
rect 170772 198698 170824 198704
rect 170876 198393 170904 199514
rect 170862 198384 170918 198393
rect 170862 198319 170918 198328
rect 170678 195528 170734 195537
rect 170678 195463 170734 195472
rect 170692 191146 170720 195463
rect 170680 191140 170732 191146
rect 170680 191082 170732 191088
rect 170968 189038 170996 199736
rect 171046 199744 171048 199753
rect 171198 199764 171226 200124
rect 171290 199918 171318 200124
rect 171382 199923 171410 200124
rect 171278 199912 171330 199918
rect 171278 199854 171330 199860
rect 171368 199914 171424 199923
rect 171368 199849 171424 199858
rect 171474 199764 171502 200124
rect 171100 199744 171102 199753
rect 171046 199679 171102 199688
rect 171152 199736 171226 199764
rect 171428 199736 171502 199764
rect 171152 199288 171180 199736
rect 171324 199640 171376 199646
rect 171324 199582 171376 199588
rect 171060 199260 171180 199288
rect 171060 198734 171088 199260
rect 171140 199164 171192 199170
rect 171140 199106 171192 199112
rect 171152 198830 171180 199106
rect 171140 198824 171192 198830
rect 171140 198766 171192 198772
rect 171060 198706 171272 198734
rect 171140 198144 171192 198150
rect 171140 198086 171192 198092
rect 171152 194886 171180 198086
rect 171140 194880 171192 194886
rect 171140 194822 171192 194828
rect 171244 191298 171272 198706
rect 171336 198422 171364 199582
rect 171324 198416 171376 198422
rect 171324 198358 171376 198364
rect 171324 198212 171376 198218
rect 171324 198154 171376 198160
rect 171336 197538 171364 198154
rect 171324 197532 171376 197538
rect 171324 197474 171376 197480
rect 171152 191270 171272 191298
rect 170956 189032 171008 189038
rect 170956 188974 171008 188980
rect 170588 188692 170640 188698
rect 170588 188634 170640 188640
rect 171152 181490 171180 191270
rect 171428 191162 171456 199736
rect 171566 199696 171594 200124
rect 171658 199889 171686 200124
rect 171644 199880 171700 199889
rect 171644 199815 171700 199824
rect 171750 199764 171778 200124
rect 171842 199918 171870 200124
rect 171934 199918 171962 200124
rect 171830 199912 171882 199918
rect 171830 199854 171882 199860
rect 171922 199912 171974 199918
rect 171922 199854 171974 199860
rect 171520 199668 171594 199696
rect 171704 199736 171778 199764
rect 171520 198665 171548 199668
rect 171600 199504 171652 199510
rect 171600 199446 171652 199452
rect 171506 198656 171562 198665
rect 171506 198591 171562 198600
rect 171508 198484 171560 198490
rect 171508 198426 171560 198432
rect 171520 197470 171548 198426
rect 171508 197464 171560 197470
rect 171508 197406 171560 197412
rect 171244 191134 171456 191162
rect 171508 191140 171560 191146
rect 171140 181484 171192 181490
rect 171140 181426 171192 181432
rect 170048 176626 170352 176654
rect 170048 147286 170076 176626
rect 171244 147490 171272 191134
rect 171508 191082 171560 191088
rect 171416 188964 171468 188970
rect 171416 188906 171468 188912
rect 171324 181484 171376 181490
rect 171324 181426 171376 181432
rect 171232 147484 171284 147490
rect 171232 147426 171284 147432
rect 170036 147280 170088 147286
rect 170036 147222 170088 147228
rect 171336 147218 171364 181426
rect 171324 147212 171376 147218
rect 171324 147154 171376 147160
rect 171428 147082 171456 188906
rect 171416 147076 171468 147082
rect 171416 147018 171468 147024
rect 171520 147014 171548 191082
rect 171612 188970 171640 199446
rect 171600 188964 171652 188970
rect 171600 188906 171652 188912
rect 171508 147008 171560 147014
rect 171508 146950 171560 146956
rect 170772 144696 170824 144702
rect 170772 144638 170824 144644
rect 170220 143064 170272 143070
rect 170220 143006 170272 143012
rect 169942 140312 169998 140321
rect 169942 140247 169998 140256
rect 169852 140140 169904 140146
rect 169852 140082 169904 140088
rect 170232 139890 170260 143006
rect 170784 139890 170812 144638
rect 171704 140622 171732 199736
rect 172026 199730 172054 200124
rect 172118 199764 172146 200124
rect 172210 199918 172238 200124
rect 172198 199912 172250 199918
rect 172302 199889 172330 200124
rect 172198 199854 172250 199860
rect 172288 199880 172344 199889
rect 172288 199815 172344 199824
rect 172394 199764 172422 200124
rect 172118 199736 172284 199764
rect 172348 199753 172422 199764
rect 171876 199708 171928 199714
rect 171876 199650 171928 199656
rect 171980 199702 172054 199730
rect 171784 198552 171836 198558
rect 171784 198494 171836 198500
rect 171796 197674 171824 198494
rect 171888 198121 171916 199650
rect 171980 199510 172008 199702
rect 172256 199646 172284 199736
rect 172334 199744 172422 199753
rect 172390 199736 172422 199744
rect 172486 199764 172514 200124
rect 172578 199918 172606 200124
rect 172566 199912 172618 199918
rect 172566 199854 172618 199860
rect 172486 199736 172560 199764
rect 172334 199679 172390 199688
rect 172060 199640 172112 199646
rect 172060 199582 172112 199588
rect 172244 199640 172296 199646
rect 172244 199582 172296 199588
rect 171968 199504 172020 199510
rect 171968 199446 172020 199452
rect 171968 199368 172020 199374
rect 171968 199310 172020 199316
rect 171874 198112 171930 198121
rect 171874 198047 171930 198056
rect 171876 197940 171928 197946
rect 171876 197882 171928 197888
rect 171784 197668 171836 197674
rect 171784 197610 171836 197616
rect 171782 196888 171838 196897
rect 171782 196823 171838 196832
rect 171796 196722 171824 196823
rect 171784 196716 171836 196722
rect 171784 196658 171836 196664
rect 171888 194954 171916 197882
rect 171876 194948 171928 194954
rect 171876 194890 171928 194896
rect 171980 191078 172008 199310
rect 172072 191185 172100 199582
rect 172152 199572 172204 199578
rect 172152 199514 172204 199520
rect 172336 199572 172388 199578
rect 172336 199514 172388 199520
rect 172428 199572 172480 199578
rect 172428 199514 172480 199520
rect 172164 198218 172192 199514
rect 172242 199472 172298 199481
rect 172242 199407 172298 199416
rect 172152 198212 172204 198218
rect 172152 198154 172204 198160
rect 172256 198014 172284 199407
rect 172348 199322 172376 199514
rect 172440 199481 172468 199514
rect 172426 199472 172482 199481
rect 172426 199407 172482 199416
rect 172348 199294 172468 199322
rect 172336 199232 172388 199238
rect 172336 199174 172388 199180
rect 172244 198008 172296 198014
rect 172244 197950 172296 197956
rect 172152 197464 172204 197470
rect 172152 197406 172204 197412
rect 172164 195974 172192 197406
rect 172152 195968 172204 195974
rect 172152 195910 172204 195916
rect 172348 193032 172376 199174
rect 172440 197656 172468 199294
rect 172532 198286 172560 199736
rect 172670 199458 172698 200124
rect 172762 199918 172790 200124
rect 172750 199912 172802 199918
rect 172750 199854 172802 199860
rect 172854 199764 172882 200124
rect 172808 199736 172882 199764
rect 172808 199578 172836 199736
rect 172946 199628 172974 200124
rect 173038 199730 173066 200124
rect 173130 199918 173158 200124
rect 173118 199912 173170 199918
rect 173118 199854 173170 199860
rect 173222 199730 173250 200124
rect 173038 199702 173112 199730
rect 172946 199600 173020 199628
rect 172796 199572 172848 199578
rect 172796 199514 172848 199520
rect 172794 199472 172850 199481
rect 172670 199430 172744 199458
rect 172520 198280 172572 198286
rect 172520 198222 172572 198228
rect 172440 197628 172652 197656
rect 172428 197532 172480 197538
rect 172428 197474 172480 197480
rect 172440 195906 172468 197474
rect 172428 195900 172480 195906
rect 172428 195842 172480 195848
rect 172348 193004 172560 193032
rect 172058 191176 172114 191185
rect 172058 191111 172114 191120
rect 171968 191072 172020 191078
rect 171968 191014 172020 191020
rect 172428 144628 172480 144634
rect 172428 144570 172480 144576
rect 171876 141636 171928 141642
rect 171876 141578 171928 141584
rect 171692 140616 171744 140622
rect 171692 140558 171744 140564
rect 171888 139890 171916 141578
rect 172440 139890 172468 144570
rect 172532 140690 172560 193004
rect 172624 191162 172652 197628
rect 172716 192846 172744 199430
rect 172794 199407 172850 199416
rect 172704 192840 172756 192846
rect 172704 192782 172756 192788
rect 172808 191298 172836 199407
rect 172808 191270 172928 191298
rect 172624 191134 172836 191162
rect 172704 191072 172756 191078
rect 172704 191014 172756 191020
rect 172612 183524 172664 183530
rect 172612 183466 172664 183472
rect 172624 147121 172652 183466
rect 172716 147150 172744 191014
rect 172808 147422 172836 191134
rect 172900 183530 172928 191270
rect 172992 191185 173020 199600
rect 173084 198694 173112 199702
rect 173176 199702 173250 199730
rect 173072 198688 173124 198694
rect 173072 198630 173124 198636
rect 173176 191321 173204 199702
rect 173314 199628 173342 200124
rect 173406 199696 173434 200124
rect 173498 199764 173526 200124
rect 173590 199918 173618 200124
rect 173578 199912 173630 199918
rect 173578 199854 173630 199860
rect 173682 199764 173710 200124
rect 173774 199889 173802 200124
rect 173760 199880 173816 199889
rect 173760 199815 173816 199824
rect 173498 199736 173572 199764
rect 173682 199736 173756 199764
rect 173544 199696 173572 199736
rect 173406 199668 173480 199696
rect 173544 199668 173664 199696
rect 173268 199600 173342 199628
rect 173268 198490 173296 199600
rect 173348 199504 173400 199510
rect 173348 199446 173400 199452
rect 173256 198484 173308 198490
rect 173256 198426 173308 198432
rect 173360 198082 173388 199446
rect 173348 198076 173400 198082
rect 173348 198018 173400 198024
rect 173162 191312 173218 191321
rect 173162 191247 173218 191256
rect 172978 191176 173034 191185
rect 172978 191111 173034 191120
rect 172888 183524 172940 183530
rect 172888 183466 172940 183472
rect 173452 182174 173480 199668
rect 173532 199572 173584 199578
rect 173532 199514 173584 199520
rect 173544 197946 173572 199514
rect 173636 198734 173664 199668
rect 173728 199238 173756 199736
rect 173866 199696 173894 200124
rect 173958 199764 173986 200124
rect 174050 199918 174078 200124
rect 174142 199918 174170 200124
rect 174234 199918 174262 200124
rect 174326 199923 174354 200124
rect 174038 199912 174090 199918
rect 174038 199854 174090 199860
rect 174130 199912 174182 199918
rect 174130 199854 174182 199860
rect 174222 199912 174274 199918
rect 174222 199854 174274 199860
rect 174312 199914 174368 199923
rect 174418 199918 174446 200124
rect 174510 199918 174538 200124
rect 174312 199849 174368 199858
rect 174406 199912 174458 199918
rect 174406 199854 174458 199860
rect 174498 199912 174550 199918
rect 174498 199854 174550 199860
rect 174084 199776 174136 199782
rect 173958 199736 174032 199764
rect 173866 199668 173940 199696
rect 173806 199472 173862 199481
rect 173806 199407 173808 199416
rect 173860 199407 173862 199416
rect 173808 199378 173860 199384
rect 173716 199232 173768 199238
rect 173716 199174 173768 199180
rect 173636 198706 173756 198734
rect 173532 197940 173584 197946
rect 173532 197882 173584 197888
rect 173728 191049 173756 198706
rect 173912 198150 173940 199668
rect 173900 198144 173952 198150
rect 173900 198086 173952 198092
rect 174004 191298 174032 199736
rect 174602 199764 174630 200124
rect 174694 199918 174722 200124
rect 174786 199918 174814 200124
rect 174682 199912 174734 199918
rect 174682 199854 174734 199860
rect 174774 199912 174826 199918
rect 174774 199854 174826 199860
rect 174878 199764 174906 200124
rect 174970 199918 174998 200124
rect 174958 199912 175010 199918
rect 174958 199854 175010 199860
rect 175062 199764 175090 200124
rect 175154 199889 175182 200124
rect 175140 199880 175196 199889
rect 175140 199815 175196 199824
rect 174602 199736 174676 199764
rect 174878 199736 174952 199764
rect 175062 199736 175136 199764
rect 174084 199718 174136 199724
rect 174096 197402 174124 199718
rect 174452 199708 174504 199714
rect 174452 199650 174504 199656
rect 174268 199572 174320 199578
rect 174320 199532 174400 199560
rect 174268 199514 174320 199520
rect 174176 199504 174228 199510
rect 174176 199446 174228 199452
rect 174084 197396 174136 197402
rect 174084 197338 174136 197344
rect 174004 191270 174124 191298
rect 173992 191208 174044 191214
rect 173992 191150 174044 191156
rect 173714 191040 173770 191049
rect 173714 190975 173770 190984
rect 173900 190596 173952 190602
rect 173900 190538 173952 190544
rect 173360 182146 173480 182174
rect 173360 176654 173388 182146
rect 172900 176626 173388 176654
rect 172796 147416 172848 147422
rect 172796 147358 172848 147364
rect 172900 147354 172928 176626
rect 172888 147348 172940 147354
rect 172888 147290 172940 147296
rect 172704 147144 172756 147150
rect 172610 147112 172666 147121
rect 172704 147086 172756 147092
rect 172610 147047 172666 147056
rect 173912 146169 173940 190538
rect 174004 146946 174032 191150
rect 173992 146940 174044 146946
rect 173992 146882 174044 146888
rect 174096 146305 174124 191270
rect 174188 190602 174216 199446
rect 174268 198960 174320 198966
rect 174268 198902 174320 198908
rect 174280 198830 174308 198902
rect 174268 198824 174320 198830
rect 174268 198766 174320 198772
rect 174268 191140 174320 191146
rect 174268 191082 174320 191088
rect 174176 190596 174228 190602
rect 174176 190538 174228 190544
rect 174176 190460 174228 190466
rect 174176 190402 174228 190408
rect 174188 150006 174216 190402
rect 174280 150113 174308 191082
rect 174266 150104 174322 150113
rect 174372 150074 174400 199532
rect 174464 198734 174492 199650
rect 174464 198706 174584 198734
rect 174452 197396 174504 197402
rect 174452 197338 174504 197344
rect 174464 192914 174492 197338
rect 174452 192908 174504 192914
rect 174452 192850 174504 192856
rect 174556 190466 174584 198706
rect 174648 196489 174676 199736
rect 174820 199640 174872 199646
rect 174820 199582 174872 199588
rect 174728 199572 174780 199578
rect 174728 199514 174780 199520
rect 174634 196480 174690 196489
rect 174634 196415 174690 196424
rect 174740 191146 174768 199514
rect 174832 198762 174860 199582
rect 174820 198756 174872 198762
rect 174820 198698 174872 198704
rect 174924 198121 174952 199736
rect 175004 199640 175056 199646
rect 175004 199582 175056 199588
rect 174910 198112 174966 198121
rect 174910 198047 174966 198056
rect 175016 195537 175044 199582
rect 175108 198734 175136 199736
rect 175246 199628 175274 200124
rect 175338 199696 175366 200124
rect 175430 199889 175458 200124
rect 175522 199918 175550 200124
rect 175614 199918 175642 200124
rect 175510 199912 175562 199918
rect 175416 199880 175472 199889
rect 175510 199854 175562 199860
rect 175602 199912 175654 199918
rect 175602 199854 175654 199860
rect 175416 199815 175472 199824
rect 175706 199764 175734 200124
rect 175462 199744 175518 199753
rect 175338 199668 175412 199696
rect 175660 199736 175734 199764
rect 175462 199679 175518 199688
rect 175556 199708 175608 199714
rect 175246 199600 175320 199628
rect 175188 199504 175240 199510
rect 175188 199446 175240 199452
rect 175200 199170 175228 199446
rect 175188 199164 175240 199170
rect 175188 199106 175240 199112
rect 175108 198706 175228 198734
rect 175002 195528 175058 195537
rect 175002 195463 175058 195472
rect 175200 194594 175228 198706
rect 175292 195673 175320 199600
rect 175278 195664 175334 195673
rect 175278 195599 175334 195608
rect 175200 194566 175320 194594
rect 175292 193214 175320 194566
rect 175016 193186 175320 193214
rect 175016 191214 175044 193186
rect 175004 191208 175056 191214
rect 175004 191150 175056 191156
rect 174728 191140 174780 191146
rect 174728 191082 174780 191088
rect 174544 190460 174596 190466
rect 174544 190402 174596 190408
rect 175280 185020 175332 185026
rect 175280 184962 175332 184968
rect 174266 150039 174322 150048
rect 174360 150068 174412 150074
rect 174360 150010 174412 150016
rect 174176 150000 174228 150006
rect 174176 149942 174228 149948
rect 175292 149870 175320 184962
rect 175280 149864 175332 149870
rect 175280 149806 175332 149812
rect 175384 149802 175412 199668
rect 175476 192545 175504 199679
rect 175556 199650 175608 199656
rect 175462 192536 175518 192545
rect 175462 192471 175518 192480
rect 175568 190454 175596 199650
rect 175660 194857 175688 199736
rect 175798 199696 175826 200124
rect 175890 199889 175918 200124
rect 175982 199918 176010 200124
rect 176074 199918 176102 200124
rect 176166 199918 176194 200124
rect 176258 199918 176286 200124
rect 175970 199912 176022 199918
rect 175876 199880 175932 199889
rect 175970 199854 176022 199860
rect 176062 199912 176114 199918
rect 176062 199854 176114 199860
rect 176154 199912 176206 199918
rect 176154 199854 176206 199860
rect 176246 199912 176298 199918
rect 176350 199889 176378 200124
rect 176246 199854 176298 199860
rect 176336 199880 176392 199889
rect 175876 199815 175932 199824
rect 176336 199815 176392 199824
rect 175924 199776 175976 199782
rect 175752 199668 175826 199696
rect 175922 199744 175924 199753
rect 176108 199776 176160 199782
rect 175976 199744 175978 199753
rect 176108 199718 176160 199724
rect 176290 199744 176346 199753
rect 175922 199679 175978 199688
rect 175752 199102 175780 199668
rect 176016 199640 176068 199646
rect 176016 199582 176068 199588
rect 175924 199504 175976 199510
rect 175924 199446 175976 199452
rect 175740 199096 175792 199102
rect 175740 199038 175792 199044
rect 175646 194848 175702 194857
rect 175646 194783 175702 194792
rect 175568 190426 175688 190454
rect 175462 187776 175518 187785
rect 175462 187711 175518 187720
rect 175476 150142 175504 187711
rect 175556 184748 175608 184754
rect 175556 184690 175608 184696
rect 175568 150210 175596 184690
rect 175556 150204 175608 150210
rect 175556 150146 175608 150152
rect 175464 150136 175516 150142
rect 175464 150078 175516 150084
rect 175660 149938 175688 190426
rect 175936 184754 175964 199446
rect 176028 193594 176056 199582
rect 176016 193588 176068 193594
rect 176016 193530 176068 193536
rect 176120 185026 176148 199718
rect 176290 199679 176346 199688
rect 176200 199640 176252 199646
rect 176200 199582 176252 199588
rect 176212 188465 176240 199582
rect 176304 197033 176332 199679
rect 176442 199628 176470 200124
rect 176396 199600 176470 199628
rect 176396 199510 176424 199600
rect 176534 199560 176562 200124
rect 176626 199764 176654 200124
rect 176718 199918 176746 200124
rect 176810 199918 176838 200124
rect 176706 199912 176758 199918
rect 176706 199854 176758 199860
rect 176798 199912 176850 199918
rect 176902 199889 176930 200124
rect 176994 199918 177022 200124
rect 176982 199912 177034 199918
rect 176798 199854 176850 199860
rect 176888 199880 176944 199889
rect 177086 199889 177114 200124
rect 176982 199854 177034 199860
rect 177072 199880 177128 199889
rect 176888 199815 176944 199824
rect 177072 199815 177128 199824
rect 177178 199782 177206 200124
rect 177270 199918 177298 200124
rect 177258 199912 177310 199918
rect 177258 199854 177310 199860
rect 176844 199776 176896 199782
rect 176626 199736 176700 199764
rect 176488 199532 176562 199560
rect 176384 199504 176436 199510
rect 176384 199446 176436 199452
rect 176290 197024 176346 197033
rect 176290 196959 176346 196968
rect 176488 191185 176516 199532
rect 176474 191176 176530 191185
rect 176474 191111 176530 191120
rect 176198 188456 176254 188465
rect 176198 188391 176254 188400
rect 176672 188057 176700 199736
rect 176844 199718 176896 199724
rect 176936 199776 176988 199782
rect 176936 199718 176988 199724
rect 177166 199776 177218 199782
rect 177362 199764 177390 200124
rect 177454 199866 177482 200124
rect 177546 199968 177574 200124
rect 177652 200110 177804 200138
rect 177546 199940 177620 199968
rect 177454 199838 177528 199866
rect 177166 199718 177218 199724
rect 177316 199736 177390 199764
rect 176750 198112 176806 198121
rect 176750 198047 176806 198056
rect 176764 197577 176792 198047
rect 176750 197568 176806 197577
rect 176750 197503 176806 197512
rect 176856 193118 176884 199718
rect 176844 193112 176896 193118
rect 176844 193054 176896 193060
rect 176844 188420 176896 188426
rect 176844 188362 176896 188368
rect 176752 188352 176804 188358
rect 176752 188294 176804 188300
rect 176658 188048 176714 188057
rect 176658 187983 176714 187992
rect 176660 187944 176712 187950
rect 176660 187886 176712 187892
rect 176108 185020 176160 185026
rect 176108 184962 176160 184968
rect 175924 184748 175976 184754
rect 175924 184690 175976 184696
rect 175648 149932 175700 149938
rect 175648 149874 175700 149880
rect 175372 149796 175424 149802
rect 175372 149738 175424 149744
rect 174082 146296 174138 146305
rect 174082 146231 174138 146240
rect 173898 146160 173954 146169
rect 173898 146095 173954 146104
rect 175556 146124 175608 146130
rect 175556 146066 175608 146072
rect 173808 144764 173860 144770
rect 173808 144706 173860 144712
rect 172980 143336 173032 143342
rect 172980 143278 173032 143284
rect 172520 140684 172572 140690
rect 172520 140626 172572 140632
rect 172992 139890 173020 143278
rect 173532 141704 173584 141710
rect 173532 141646 173584 141652
rect 173544 139890 173572 141646
rect 173820 140162 173848 144706
rect 175464 143472 175516 143478
rect 175464 143414 175516 143420
rect 174636 143404 174688 143410
rect 174636 143346 174688 143352
rect 168820 139862 169156 139890
rect 169372 139862 169708 139890
rect 169924 139862 170260 139890
rect 170476 139862 170812 139890
rect 171028 139874 171180 139890
rect 171028 139868 171192 139874
rect 171028 139862 171140 139868
rect 171580 139862 171916 139890
rect 172132 139862 172468 139890
rect 172684 139862 173020 139890
rect 173236 139862 173572 139890
rect 173774 140134 173848 140162
rect 173774 139876 173802 140134
rect 174648 139890 174676 143346
rect 175188 141772 175240 141778
rect 175188 141714 175240 141720
rect 175200 139890 175228 141714
rect 175476 140162 175504 143414
rect 174340 139862 174676 139890
rect 174892 139862 175228 139890
rect 175430 140134 175504 140162
rect 175430 139876 175458 140134
rect 175568 139890 175596 146066
rect 176568 143268 176620 143274
rect 176568 143210 176620 143216
rect 176580 140162 176608 143210
rect 176672 141681 176700 187886
rect 176658 141672 176714 141681
rect 176658 141607 176714 141616
rect 176764 141273 176792 188294
rect 176856 150346 176884 188362
rect 176948 150414 176976 199718
rect 177316 188329 177344 199736
rect 177396 199572 177448 199578
rect 177396 199514 177448 199520
rect 177408 198422 177436 199514
rect 177396 198416 177448 198422
rect 177396 198358 177448 198364
rect 177500 188465 177528 199838
rect 177592 199510 177620 199940
rect 177672 199912 177724 199918
rect 177672 199854 177724 199860
rect 177684 199578 177712 199854
rect 177672 199572 177724 199578
rect 177672 199514 177724 199520
rect 177580 199504 177632 199510
rect 177580 199446 177632 199452
rect 177486 188456 177542 188465
rect 177486 188391 177542 188400
rect 177776 188358 177804 200110
rect 177868 196858 177896 200602
rect 178222 200424 178278 200433
rect 178222 200359 178278 200368
rect 178868 200388 178920 200394
rect 178040 200252 178092 200258
rect 178040 200194 178092 200200
rect 177948 199572 178000 199578
rect 177948 199514 178000 199520
rect 177856 196852 177908 196858
rect 177856 196794 177908 196800
rect 177960 188426 177988 199514
rect 178052 199306 178080 200194
rect 178236 199578 178264 200359
rect 178868 200330 178920 200336
rect 178880 200161 178908 200330
rect 178866 200152 178922 200161
rect 178866 200087 178922 200096
rect 178224 199572 178276 199578
rect 178224 199514 178276 199520
rect 178132 199504 178184 199510
rect 178132 199446 178184 199452
rect 178040 199300 178092 199306
rect 178040 199242 178092 199248
rect 177948 188420 178000 188426
rect 177948 188362 178000 188368
rect 177764 188352 177816 188358
rect 177302 188320 177358 188329
rect 177764 188294 177816 188300
rect 177302 188255 177358 188264
rect 178144 187950 178172 199446
rect 178776 198960 178828 198966
rect 178776 198902 178828 198908
rect 178684 198620 178736 198626
rect 178684 198562 178736 198568
rect 178314 195120 178370 195129
rect 178314 195055 178370 195064
rect 178132 187944 178184 187950
rect 178132 187886 178184 187892
rect 178328 176654 178356 195055
rect 178696 192574 178724 198562
rect 178788 195974 178816 198902
rect 178788 195946 178908 195974
rect 178684 192568 178736 192574
rect 178684 192510 178736 192516
rect 178328 176626 178724 176654
rect 176936 150408 176988 150414
rect 176936 150350 176988 150356
rect 176844 150340 176896 150346
rect 176844 150282 176896 150288
rect 178696 148782 178724 176626
rect 178684 148776 178736 148782
rect 178684 148718 178736 148724
rect 178224 147620 178276 147626
rect 178224 147562 178276 147568
rect 178040 147552 178092 147558
rect 178040 147494 178092 147500
rect 177396 143132 177448 143138
rect 177396 143074 177448 143080
rect 176750 141264 176806 141273
rect 176750 141199 176806 141208
rect 176534 140134 176608 140162
rect 175568 139862 175996 139890
rect 176534 139876 176562 140134
rect 177408 139890 177436 143074
rect 177948 142724 178000 142730
rect 177948 142666 178000 142672
rect 177960 139890 177988 142666
rect 178052 140758 178080 147494
rect 178132 146192 178184 146198
rect 178132 146134 178184 146140
rect 178040 140752 178092 140758
rect 178040 140694 178092 140700
rect 177100 139862 177436 139890
rect 177652 139862 177988 139890
rect 178144 139890 178172 146134
rect 178236 142730 178264 147562
rect 178408 146804 178460 146810
rect 178408 146746 178460 146752
rect 178316 146260 178368 146266
rect 178316 146202 178368 146208
rect 178224 142724 178276 142730
rect 178224 142666 178276 142672
rect 178328 139890 178356 146202
rect 178420 143342 178448 146746
rect 178408 143336 178460 143342
rect 178408 143278 178460 143284
rect 178144 139862 178204 139890
rect 178328 139862 178756 139890
rect 171140 139810 171192 139816
rect 178880 139369 178908 195946
rect 180076 147674 180104 200602
rect 183836 200592 183888 200598
rect 183836 200534 183888 200540
rect 186872 200592 186924 200598
rect 186872 200534 186924 200540
rect 181904 200116 181956 200122
rect 181904 200058 181956 200064
rect 180340 199436 180392 199442
rect 180340 199378 180392 199384
rect 180156 198824 180208 198830
rect 180156 198766 180208 198772
rect 179984 147646 180104 147674
rect 179604 146872 179656 146878
rect 179604 146814 179656 146820
rect 179420 145376 179472 145382
rect 179420 145318 179472 145324
rect 179432 143138 179460 145318
rect 179512 144832 179564 144838
rect 179512 144774 179564 144780
rect 179524 143478 179552 144774
rect 179512 143472 179564 143478
rect 179512 143414 179564 143420
rect 179616 143206 179644 146814
rect 179696 146736 179748 146742
rect 179696 146678 179748 146684
rect 179708 143410 179736 146678
rect 179788 145580 179840 145586
rect 179788 145522 179840 145528
rect 179696 143404 179748 143410
rect 179696 143346 179748 143352
rect 179604 143200 179656 143206
rect 179604 143142 179656 143148
rect 179420 143132 179472 143138
rect 179420 143074 179472 143080
rect 179800 142154 179828 145522
rect 179432 142126 179828 142154
rect 178960 140752 179012 140758
rect 178960 140694 179012 140700
rect 178972 139890 179000 140694
rect 179052 140616 179104 140622
rect 179052 140558 179104 140564
rect 179064 140185 179092 140558
rect 179050 140176 179106 140185
rect 179050 140111 179106 140120
rect 179432 139890 179460 142126
rect 178972 139862 179308 139890
rect 179432 139862 179860 139890
rect 124494 139360 124550 139369
rect 124494 139295 124550 139304
rect 125506 139360 125562 139369
rect 125506 139295 125562 139304
rect 125966 139360 126022 139369
rect 125966 139295 126022 139304
rect 126150 139360 126206 139369
rect 126150 139295 126206 139304
rect 127622 139360 127678 139369
rect 127622 139295 127678 139304
rect 130014 139360 130070 139369
rect 130014 139295 130070 139304
rect 131026 139360 131082 139369
rect 131026 139295 131082 139304
rect 132222 139360 132278 139369
rect 132222 139295 132278 139304
rect 149610 139360 149666 139369
rect 149610 139295 149666 139304
rect 150990 139360 151046 139369
rect 150990 139295 151046 139304
rect 155222 139360 155278 139369
rect 155222 139295 155278 139304
rect 155774 139360 155830 139369
rect 155774 139295 155830 139304
rect 159546 139360 159602 139369
rect 159546 139295 159602 139304
rect 159822 139360 159878 139369
rect 159822 139295 159878 139304
rect 165342 139360 165398 139369
rect 165342 139295 165398 139304
rect 178866 139360 178922 139369
rect 179984 139346 180012 147646
rect 180168 142154 180196 198766
rect 180248 196580 180300 196586
rect 180248 196522 180300 196528
rect 180076 142126 180196 142154
rect 180076 140282 180104 142126
rect 180156 140684 180208 140690
rect 180156 140626 180208 140632
rect 180064 140276 180116 140282
rect 180064 140218 180116 140224
rect 180168 139777 180196 140626
rect 180260 140622 180288 196522
rect 180352 145450 180380 199378
rect 181076 198960 181128 198966
rect 181076 198902 181128 198908
rect 180432 197668 180484 197674
rect 180432 197610 180484 197616
rect 180444 145518 180472 197610
rect 181088 157334 181116 198902
rect 181916 198626 181944 200058
rect 182824 199436 182876 199442
rect 182824 199378 182876 199384
rect 181904 198620 181956 198626
rect 181904 198562 181956 198568
rect 181442 198248 181498 198257
rect 181442 198183 181444 198192
rect 181496 198183 181498 198192
rect 181444 198154 181496 198160
rect 181628 197600 181680 197606
rect 181628 197542 181680 197548
rect 181536 192432 181588 192438
rect 181536 192374 181588 192380
rect 181444 192364 181496 192370
rect 181444 192306 181496 192312
rect 181088 157306 181208 157334
rect 180892 148368 180944 148374
rect 180892 148310 180944 148316
rect 180432 145512 180484 145518
rect 180432 145454 180484 145460
rect 180340 145444 180392 145450
rect 180340 145386 180392 145392
rect 180340 141976 180392 141982
rect 180340 141918 180392 141924
rect 180248 140616 180300 140622
rect 180248 140558 180300 140564
rect 180154 139768 180210 139777
rect 180154 139703 180210 139712
rect 180064 139664 180116 139670
rect 180352 139618 180380 141918
rect 180904 139890 180932 148310
rect 181180 139890 181208 157306
rect 181456 140350 181484 192306
rect 181548 143478 181576 192374
rect 181536 143472 181588 143478
rect 181536 143414 181588 143420
rect 181444 140344 181496 140350
rect 181444 140286 181496 140292
rect 181640 140049 181668 197542
rect 182456 143200 182508 143206
rect 182456 143142 182508 143148
rect 182088 142996 182140 143002
rect 182088 142938 182140 142944
rect 182100 142730 182128 142938
rect 182088 142724 182140 142730
rect 182088 142666 182140 142672
rect 182468 142154 182496 143142
rect 182284 142126 182496 142154
rect 182088 141908 182140 141914
rect 182088 141850 182140 141856
rect 182100 141030 182128 141850
rect 182088 141024 182140 141030
rect 182088 140966 182140 140972
rect 182100 140162 182128 140966
rect 182284 140593 182312 142126
rect 182836 140962 182864 199378
rect 183006 197160 183062 197169
rect 183006 197095 183062 197104
rect 182916 194404 182968 194410
rect 182916 194346 182968 194352
rect 182824 140956 182876 140962
rect 182824 140898 182876 140904
rect 182270 140584 182326 140593
rect 182270 140519 182326 140528
rect 182054 140134 182128 140162
rect 181626 140040 181682 140049
rect 181626 139975 181682 139984
rect 180904 139862 180964 139890
rect 181180 139862 181516 139890
rect 182054 139876 182082 140134
rect 182284 139890 182312 140519
rect 182836 139890 182864 140898
rect 182928 140486 182956 194346
rect 183020 144906 183048 197095
rect 183100 193180 183152 193186
rect 183100 193122 183152 193128
rect 183008 144900 183060 144906
rect 183008 144842 183060 144848
rect 183112 142798 183140 193122
rect 183192 152312 183244 152318
rect 183192 152254 183244 152260
rect 183100 142792 183152 142798
rect 183100 142734 183152 142740
rect 183204 141846 183232 152254
rect 183744 142656 183796 142662
rect 183744 142598 183796 142604
rect 183756 142186 183784 142598
rect 183744 142180 183796 142186
rect 183744 142122 183796 142128
rect 183192 141840 183244 141846
rect 183192 141782 183244 141788
rect 182916 140480 182968 140486
rect 182916 140422 182968 140428
rect 183756 140162 183784 142122
rect 183710 140134 183784 140162
rect 183466 140040 183522 140049
rect 183466 139975 183522 139984
rect 182284 139862 182620 139890
rect 182836 139862 183172 139890
rect 180116 139612 180412 139618
rect 180064 139606 180412 139612
rect 180076 139590 180412 139606
rect 181180 139534 181208 139862
rect 183480 139806 183508 139975
rect 183710 139876 183738 140134
rect 183468 139800 183520 139806
rect 183468 139742 183520 139748
rect 181168 139528 181220 139534
rect 183848 139505 183876 200534
rect 186884 200190 186912 200534
rect 186780 200184 186832 200190
rect 186780 200126 186832 200132
rect 186872 200184 186924 200190
rect 186872 200126 186924 200132
rect 186596 199572 186648 199578
rect 186596 199514 186648 199520
rect 186412 199096 186464 199102
rect 186412 199038 186464 199044
rect 186424 198830 186452 199038
rect 186412 198824 186464 198830
rect 186412 198766 186464 198772
rect 186410 194848 186466 194857
rect 186410 194783 186466 194792
rect 184204 194676 184256 194682
rect 184204 194618 184256 194624
rect 184216 150278 184244 194618
rect 185952 153196 186004 153202
rect 185952 153138 186004 153144
rect 185584 153128 185636 153134
rect 185584 153070 185636 153076
rect 184296 153060 184348 153066
rect 184296 153002 184348 153008
rect 184204 150272 184256 150278
rect 184204 150214 184256 150220
rect 184112 148640 184164 148646
rect 184112 148582 184164 148588
rect 184124 140554 184152 148582
rect 184112 140548 184164 140554
rect 184112 140490 184164 140496
rect 184308 140214 184336 153002
rect 184388 152856 184440 152862
rect 184388 152798 184440 152804
rect 184296 140208 184348 140214
rect 184296 140150 184348 140156
rect 184400 139942 184428 152798
rect 184756 152720 184808 152726
rect 184756 152662 184808 152668
rect 184572 152380 184624 152386
rect 184572 152322 184624 152328
rect 184480 143132 184532 143138
rect 184480 143074 184532 143080
rect 184388 139936 184440 139942
rect 184388 139878 184440 139884
rect 184018 139632 184074 139641
rect 184492 139618 184520 143074
rect 184584 140962 184612 152322
rect 184664 149728 184716 149734
rect 184664 149670 184716 149676
rect 184572 140956 184624 140962
rect 184572 140898 184624 140904
rect 184676 140146 184704 149670
rect 184768 140758 184796 152662
rect 184756 140752 184808 140758
rect 184756 140694 184808 140700
rect 184664 140140 184716 140146
rect 184664 140082 184716 140088
rect 184664 139732 184716 139738
rect 184664 139674 184716 139680
rect 184676 139641 184704 139674
rect 184074 139590 184520 139618
rect 184662 139632 184718 139641
rect 184572 139596 184624 139602
rect 184018 139567 184074 139576
rect 184662 139567 184718 139576
rect 184572 139538 184624 139544
rect 184584 139505 184612 139538
rect 185596 139534 185624 153070
rect 185676 152924 185728 152930
rect 185676 152866 185728 152872
rect 185688 146962 185716 152866
rect 185860 152448 185912 152454
rect 185860 152390 185912 152396
rect 185688 146934 185808 146962
rect 185676 143404 185728 143410
rect 185676 143346 185728 143352
rect 185584 139528 185636 139534
rect 181168 139470 181220 139476
rect 183834 139496 183890 139505
rect 183834 139431 183890 139440
rect 184386 139496 184442 139505
rect 184570 139496 184626 139505
rect 184442 139454 184520 139482
rect 184386 139431 184442 139440
rect 180154 139360 180210 139369
rect 179984 139318 180154 139346
rect 178866 139295 178922 139304
rect 184492 139346 184520 139454
rect 185044 139466 185532 139482
rect 185584 139470 185636 139476
rect 184570 139431 184626 139440
rect 185032 139460 185532 139466
rect 185084 139454 185532 139460
rect 185032 139402 185084 139408
rect 185504 139346 185532 139454
rect 185688 139346 185716 143346
rect 185780 140418 185808 146934
rect 185768 140412 185820 140418
rect 185768 140354 185820 140360
rect 185872 140185 185900 152390
rect 185964 143342 185992 153138
rect 186044 152992 186096 152998
rect 186044 152934 186096 152940
rect 185952 143336 186004 143342
rect 185952 143278 186004 143284
rect 185952 142180 186004 142186
rect 185952 142122 186004 142128
rect 185858 140176 185914 140185
rect 185858 140111 185914 140120
rect 185964 140026 185992 142122
rect 185918 139998 185992 140026
rect 185918 139876 185946 139998
rect 186056 139398 186084 152934
rect 186136 152788 186188 152794
rect 186136 152730 186188 152736
rect 186148 139466 186176 152730
rect 186424 144430 186452 194783
rect 186412 144424 186464 144430
rect 186412 144366 186464 144372
rect 186226 140176 186282 140185
rect 186226 140111 186282 140120
rect 186240 139777 186268 140111
rect 186226 139768 186282 139777
rect 186226 139703 186282 139712
rect 186136 139460 186188 139466
rect 186136 139402 186188 139408
rect 184492 139318 184828 139346
rect 185504 139318 185716 139346
rect 186044 139392 186096 139398
rect 186044 139334 186096 139340
rect 180154 139295 180210 139304
rect 177762 80744 177818 80753
rect 131948 80708 132000 80714
rect 131948 80650 132000 80656
rect 132132 80708 132184 80714
rect 177652 80702 177762 80730
rect 177946 80744 178002 80753
rect 177818 80702 177896 80730
rect 177762 80679 177818 80688
rect 132132 80650 132184 80656
rect 131854 80472 131910 80481
rect 131854 80407 131910 80416
rect 131868 80374 131896 80407
rect 131856 80368 131908 80374
rect 124126 80336 124182 80345
rect 131856 80310 131908 80316
rect 124126 80271 124182 80280
rect 131028 80300 131080 80306
rect 124034 78432 124090 78441
rect 124034 78367 124090 78376
rect 123392 77920 123444 77926
rect 123392 77862 123444 77868
rect 124048 74361 124076 78367
rect 124034 74352 124090 74361
rect 124034 74287 124090 74296
rect 124140 72865 124168 80271
rect 131028 80242 131080 80248
rect 127532 80232 127584 80238
rect 127532 80174 127584 80180
rect 126980 79892 127032 79898
rect 126980 79834 127032 79840
rect 125692 79552 125744 79558
rect 125692 79494 125744 79500
rect 125600 79484 125652 79490
rect 125600 79426 125652 79432
rect 125612 76090 125640 79426
rect 124864 76084 124916 76090
rect 124864 76026 124916 76032
rect 125600 76084 125652 76090
rect 125600 76026 125652 76032
rect 124126 72856 124182 72865
rect 124126 72791 124182 72800
rect 123116 71324 123168 71330
rect 123116 71266 123168 71272
rect 122564 69760 122616 69766
rect 122564 69702 122616 69708
rect 121460 4140 121512 4146
rect 121460 4082 121512 4088
rect 123484 4140 123536 4146
rect 123484 4082 123536 4088
rect 122288 4072 122340 4078
rect 122288 4014 122340 4020
rect 120724 3528 120776 3534
rect 120724 3470 120776 3476
rect 120736 3330 120764 3470
rect 120724 3324 120776 3330
rect 120724 3266 120776 3272
rect 122300 480 122328 4014
rect 123496 480 123524 4082
rect 124876 4078 124904 76026
rect 125704 73234 125732 79494
rect 126992 78266 127020 79834
rect 127440 79552 127492 79558
rect 127440 79494 127492 79500
rect 127452 78742 127480 79494
rect 127544 79490 127572 80174
rect 130842 79520 130898 79529
rect 127532 79484 127584 79490
rect 130842 79455 130898 79464
rect 127532 79426 127584 79432
rect 128360 79416 128412 79422
rect 128360 79358 128412 79364
rect 127440 78736 127492 78742
rect 127440 78678 127492 78684
rect 126980 78260 127032 78266
rect 126980 78202 127032 78208
rect 127164 78192 127216 78198
rect 127164 78134 127216 78140
rect 127176 76702 127204 78134
rect 127164 76696 127216 76702
rect 127164 76638 127216 76644
rect 124956 73228 125008 73234
rect 124956 73170 125008 73176
rect 125692 73228 125744 73234
rect 125692 73170 125744 73176
rect 124968 4146 124996 73170
rect 124956 4140 125008 4146
rect 124956 4082 125008 4088
rect 124864 4072 124916 4078
rect 124864 4014 124916 4020
rect 125876 4072 125928 4078
rect 125876 4014 125928 4020
rect 124680 3868 124732 3874
rect 124680 3810 124732 3816
rect 124692 480 124720 3810
rect 125888 480 125916 4014
rect 128176 3596 128228 3602
rect 128176 3538 128228 3544
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 126992 480 127020 3470
rect 128188 480 128216 3538
rect 128372 490 128400 79358
rect 130384 79348 130436 79354
rect 130384 79290 130436 79296
rect 129832 77988 129884 77994
rect 129832 77930 129884 77936
rect 129740 73772 129792 73778
rect 129740 73714 129792 73720
rect 128452 69624 128504 69630
rect 128452 69566 128504 69572
rect 128464 3534 128492 69566
rect 128452 3528 128504 3534
rect 128452 3470 128504 3476
rect 129752 3210 129780 73714
rect 129844 3618 129872 77930
rect 129924 74724 129976 74730
rect 129924 74666 129976 74672
rect 129936 72350 129964 74666
rect 129924 72344 129976 72350
rect 129924 72286 129976 72292
rect 129936 4078 129964 72286
rect 129924 4072 129976 4078
rect 129924 4014 129976 4020
rect 129844 3590 129964 3618
rect 130396 3602 130424 79290
rect 130660 78056 130712 78062
rect 130660 77998 130712 78004
rect 130672 77858 130700 77998
rect 130660 77852 130712 77858
rect 130660 77794 130712 77800
rect 130752 75676 130804 75682
rect 130752 75618 130804 75624
rect 130764 67634 130792 75618
rect 130856 72468 130884 79455
rect 131040 79422 131068 80242
rect 131960 80102 131988 80650
rect 132144 80481 132172 80650
rect 132224 80640 132276 80646
rect 132224 80582 132276 80588
rect 177868 80594 177896 80702
rect 178406 80744 178462 80753
rect 177946 80679 177948 80688
rect 178000 80679 178002 80688
rect 178040 80708 178092 80714
rect 177948 80650 178000 80656
rect 182546 80744 182602 80753
rect 178406 80679 178462 80688
rect 178592 80708 178644 80714
rect 178040 80650 178092 80656
rect 132130 80472 132186 80481
rect 132236 80442 132264 80582
rect 177868 80566 177988 80594
rect 132130 80407 132186 80416
rect 132224 80436 132276 80442
rect 132224 80378 132276 80384
rect 177764 80232 177816 80238
rect 177764 80174 177816 80180
rect 177856 80232 177908 80238
rect 177856 80174 177908 80180
rect 131948 80096 132000 80102
rect 131948 80038 132000 80044
rect 132052 80022 132388 80050
rect 131762 79928 131818 79937
rect 131762 79863 131818 79872
rect 131028 79416 131080 79422
rect 131028 79358 131080 79364
rect 131026 78704 131082 78713
rect 131026 78639 131082 78648
rect 131040 77654 131068 78639
rect 131304 78532 131356 78538
rect 131304 78474 131356 78480
rect 131028 77648 131080 77654
rect 131028 77590 131080 77596
rect 131040 75682 131068 77590
rect 131118 76664 131174 76673
rect 131118 76599 131174 76608
rect 131028 75676 131080 75682
rect 131028 75618 131080 75624
rect 130856 72440 131068 72468
rect 130764 67606 130976 67634
rect 129936 3398 129964 3590
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 130948 3466 130976 67606
rect 131040 3942 131068 72440
rect 131028 3936 131080 3942
rect 131028 3878 131080 3884
rect 130936 3460 130988 3466
rect 130936 3402 130988 3408
rect 129924 3392 129976 3398
rect 129924 3334 129976 3340
rect 129752 3182 130608 3210
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128372 462 128952 490
rect 130580 480 130608 3182
rect 128924 354 128952 462
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131132 354 131160 76599
rect 131316 64874 131344 78474
rect 131580 77988 131632 77994
rect 131580 77930 131632 77936
rect 131592 76673 131620 77930
rect 131578 76664 131634 76673
rect 131578 76599 131634 76608
rect 131224 64846 131344 64874
rect 131224 3534 131252 64846
rect 131212 3528 131264 3534
rect 131212 3470 131264 3476
rect 131776 3330 131804 79863
rect 132052 78577 132080 80022
rect 132466 79948 132494 80036
rect 132236 79920 132494 79948
rect 132236 79665 132264 79920
rect 132558 79880 132586 80036
rect 132328 79852 132586 79880
rect 132222 79656 132278 79665
rect 132222 79591 132278 79600
rect 132222 79520 132278 79529
rect 132222 79455 132278 79464
rect 132236 78713 132264 79455
rect 132222 78704 132278 78713
rect 132222 78639 132278 78648
rect 132038 78568 132094 78577
rect 132038 78503 132094 78512
rect 132328 78266 132356 79852
rect 132650 79744 132678 80036
rect 132742 79966 132770 80036
rect 132834 79971 132862 80036
rect 132730 79960 132782 79966
rect 132730 79902 132782 79908
rect 132820 79962 132876 79971
rect 132820 79897 132876 79906
rect 132926 79898 132954 80036
rect 132914 79892 132966 79898
rect 132914 79834 132966 79840
rect 133018 79812 133046 80036
rect 133110 79966 133138 80036
rect 133202 79971 133230 80036
rect 133098 79960 133150 79966
rect 133098 79902 133150 79908
rect 133188 79962 133244 79971
rect 133188 79897 133244 79906
rect 133018 79784 133092 79812
rect 133064 79744 133092 79784
rect 133294 79744 133322 80036
rect 133386 79966 133414 80036
rect 133374 79960 133426 79966
rect 133374 79902 133426 79908
rect 133478 79898 133506 80036
rect 133570 79971 133598 80036
rect 133556 79962 133612 79971
rect 133662 79966 133690 80036
rect 133466 79892 133518 79898
rect 133556 79897 133612 79906
rect 133650 79960 133702 79966
rect 133650 79902 133702 79908
rect 133466 79834 133518 79840
rect 133754 79778 133782 80036
rect 133846 79966 133874 80036
rect 133834 79960 133886 79966
rect 133938 79937 133966 80036
rect 134030 79966 134058 80036
rect 134122 79966 134150 80036
rect 134018 79960 134070 79966
rect 133834 79902 133886 79908
rect 133924 79928 133980 79937
rect 134018 79902 134070 79908
rect 134110 79960 134162 79966
rect 134110 79902 134162 79908
rect 133924 79863 133980 79872
rect 134214 79830 134242 80036
rect 134306 79937 134334 80036
rect 134292 79928 134348 79937
rect 134292 79863 134348 79872
rect 133880 79824 133932 79830
rect 132604 79716 132678 79744
rect 132788 79716 133092 79744
rect 133248 79716 133322 79744
rect 133420 79756 133472 79762
rect 132408 79688 132460 79694
rect 132408 79630 132460 79636
rect 132420 79286 132448 79630
rect 132408 79280 132460 79286
rect 132408 79222 132460 79228
rect 132408 78804 132460 78810
rect 132408 78746 132460 78752
rect 132420 78538 132448 78746
rect 132500 78736 132552 78742
rect 132500 78678 132552 78684
rect 132512 78538 132540 78678
rect 132604 78606 132632 79716
rect 132684 79416 132736 79422
rect 132684 79358 132736 79364
rect 132696 78606 132724 79358
rect 132592 78600 132644 78606
rect 132592 78542 132644 78548
rect 132684 78600 132736 78606
rect 132684 78542 132736 78548
rect 132408 78532 132460 78538
rect 132408 78474 132460 78480
rect 132500 78532 132552 78538
rect 132500 78474 132552 78480
rect 132316 78260 132368 78266
rect 132316 78202 132368 78208
rect 131856 76356 131908 76362
rect 131856 76298 131908 76304
rect 131868 4146 131896 76298
rect 132592 75200 132644 75206
rect 132592 75142 132644 75148
rect 132684 75200 132736 75206
rect 132684 75142 132736 75148
rect 132604 74934 132632 75142
rect 132592 74928 132644 74934
rect 132592 74870 132644 74876
rect 132696 60654 132724 75142
rect 132788 63510 132816 79716
rect 133052 79620 133104 79626
rect 133052 79562 133104 79568
rect 132868 79552 132920 79558
rect 132868 79494 132920 79500
rect 132880 77858 132908 79494
rect 132868 77852 132920 77858
rect 132868 77794 132920 77800
rect 132776 63504 132828 63510
rect 132776 63446 132828 63452
rect 132684 60648 132736 60654
rect 132684 60590 132736 60596
rect 132880 40730 132908 77794
rect 132960 77716 133012 77722
rect 132960 77658 133012 77664
rect 132972 73778 133000 77658
rect 132960 73772 133012 73778
rect 132960 73714 133012 73720
rect 133064 53786 133092 79562
rect 133248 73817 133276 79716
rect 133754 79750 133828 79778
rect 133880 79766 133932 79772
rect 133972 79824 134024 79830
rect 133972 79766 134024 79772
rect 134202 79824 134254 79830
rect 134202 79766 134254 79772
rect 133420 79698 133472 79704
rect 133326 79656 133382 79665
rect 133326 79591 133328 79600
rect 133380 79591 133382 79600
rect 133432 79608 133460 79698
rect 133696 79688 133748 79694
rect 133696 79630 133748 79636
rect 133604 79620 133656 79626
rect 133432 79580 133552 79608
rect 133328 79562 133380 79568
rect 133234 73808 133290 73817
rect 133234 73743 133290 73752
rect 133340 71774 133368 79562
rect 133340 71746 133460 71774
rect 133432 64190 133460 71746
rect 133524 70394 133552 79580
rect 133604 79562 133656 79568
rect 133616 79529 133644 79562
rect 133602 79520 133658 79529
rect 133602 79455 133658 79464
rect 133604 78736 133656 78742
rect 133604 78678 133656 78684
rect 133616 72962 133644 78678
rect 133604 72956 133656 72962
rect 133604 72898 133656 72904
rect 133524 70366 133644 70394
rect 133420 64184 133472 64190
rect 133420 64126 133472 64132
rect 133616 56574 133644 70366
rect 133708 69562 133736 79630
rect 133800 75206 133828 79750
rect 133892 78742 133920 79766
rect 133880 78736 133932 78742
rect 133880 78678 133932 78684
rect 133984 78674 134012 79766
rect 134064 79756 134116 79762
rect 134398 79744 134426 80036
rect 134490 79898 134518 80036
rect 134478 79892 134530 79898
rect 134478 79834 134530 79840
rect 134582 79744 134610 80036
rect 134674 79966 134702 80036
rect 134662 79960 134714 79966
rect 134662 79902 134714 79908
rect 134662 79824 134714 79830
rect 134662 79766 134714 79772
rect 134064 79698 134116 79704
rect 134352 79716 134426 79744
rect 134536 79716 134610 79744
rect 133972 78668 134024 78674
rect 133972 78610 134024 78616
rect 133970 78568 134026 78577
rect 133970 78503 134026 78512
rect 133788 75200 133840 75206
rect 133788 75142 133840 75148
rect 133984 70394 134012 78503
rect 134076 77761 134104 79698
rect 134246 79656 134302 79665
rect 134156 79620 134208 79626
rect 134352 79626 134380 79716
rect 134536 79676 134564 79716
rect 134444 79648 134564 79676
rect 134246 79591 134302 79600
rect 134340 79620 134392 79626
rect 134156 79562 134208 79568
rect 134168 77858 134196 79562
rect 134156 77852 134208 77858
rect 134156 77794 134208 77800
rect 134062 77752 134118 77761
rect 134062 77687 134118 77696
rect 134260 76566 134288 79591
rect 134340 79562 134392 79568
rect 134340 79484 134392 79490
rect 134340 79426 134392 79432
rect 134248 76560 134300 76566
rect 134248 76502 134300 76508
rect 134352 75914 134380 79426
rect 134444 78826 134472 79648
rect 134674 79642 134702 79766
rect 134766 79762 134794 80036
rect 134858 79966 134886 80036
rect 134846 79960 134898 79966
rect 134846 79902 134898 79908
rect 134950 79898 134978 80036
rect 134938 79892 134990 79898
rect 134938 79834 134990 79840
rect 134754 79756 134806 79762
rect 135042 79744 135070 80036
rect 135134 79778 135162 80036
rect 135226 79937 135254 80036
rect 135318 79966 135346 80036
rect 135306 79960 135358 79966
rect 135212 79928 135268 79937
rect 135306 79902 135358 79908
rect 135212 79863 135268 79872
rect 135134 79750 135208 79778
rect 134754 79698 134806 79704
rect 134996 79716 135070 79744
rect 134892 79688 134944 79694
rect 134674 79614 134840 79642
rect 134892 79630 134944 79636
rect 134616 79552 134668 79558
rect 134668 79512 134748 79540
rect 134616 79494 134668 79500
rect 134444 78798 134656 78826
rect 134524 78736 134576 78742
rect 134524 78678 134576 78684
rect 134432 77852 134484 77858
rect 134432 77794 134484 77800
rect 134076 75886 134380 75914
rect 134076 74225 134104 75886
rect 134248 75676 134300 75682
rect 134248 75618 134300 75624
rect 134062 74216 134118 74225
rect 134062 74151 134118 74160
rect 134156 71392 134208 71398
rect 134156 71334 134208 71340
rect 133892 70366 134012 70394
rect 133696 69556 133748 69562
rect 133696 69498 133748 69504
rect 133604 56568 133656 56574
rect 133604 56510 133656 56516
rect 133052 53780 133104 53786
rect 133052 53722 133104 53728
rect 132868 40724 132920 40730
rect 132868 40666 132920 40672
rect 133892 39370 133920 70366
rect 133880 39364 133932 39370
rect 133880 39306 133932 39312
rect 134168 7614 134196 71334
rect 134260 51066 134288 75618
rect 134340 74996 134392 75002
rect 134340 74938 134392 74944
rect 134352 66094 134380 74938
rect 134340 66088 134392 66094
rect 134340 66030 134392 66036
rect 134444 60722 134472 77794
rect 134432 60716 134484 60722
rect 134432 60658 134484 60664
rect 134248 51060 134300 51066
rect 134248 51002 134300 51008
rect 134156 7608 134208 7614
rect 134156 7550 134208 7556
rect 131856 4140 131908 4146
rect 131856 4082 131908 4088
rect 134536 4010 134564 78678
rect 134628 71602 134656 78798
rect 134720 75682 134748 79512
rect 134708 75676 134760 75682
rect 134708 75618 134760 75624
rect 134616 71596 134668 71602
rect 134616 71538 134668 71544
rect 134812 71398 134840 79614
rect 134800 71392 134852 71398
rect 134800 71334 134852 71340
rect 134904 70394 134932 79630
rect 134996 77042 135024 79716
rect 135180 79665 135208 79750
rect 135410 79676 135438 80036
rect 135166 79656 135222 79665
rect 135364 79648 135438 79676
rect 135166 79591 135222 79600
rect 135260 79620 135312 79626
rect 135260 79562 135312 79568
rect 135076 79484 135128 79490
rect 135076 79426 135128 79432
rect 134984 77036 135036 77042
rect 134984 76978 135036 76984
rect 135088 75993 135116 79426
rect 135166 77752 135222 77761
rect 135166 77687 135222 77696
rect 135074 75984 135130 75993
rect 135074 75919 135130 75928
rect 135180 75002 135208 77687
rect 135168 74996 135220 75002
rect 135168 74938 135220 74944
rect 135272 72826 135300 79562
rect 135364 77625 135392 79648
rect 135502 79608 135530 80036
rect 135594 79830 135622 80036
rect 135582 79824 135634 79830
rect 135582 79766 135634 79772
rect 135686 79778 135714 80036
rect 135778 79898 135806 80036
rect 135766 79892 135818 79898
rect 135766 79834 135818 79840
rect 135686 79750 135760 79778
rect 135732 79665 135760 79750
rect 135870 79744 135898 80036
rect 135962 79898 135990 80036
rect 136054 79898 136082 80036
rect 135950 79892 136002 79898
rect 135950 79834 136002 79840
rect 136042 79892 136094 79898
rect 136042 79834 136094 79840
rect 135824 79716 135898 79744
rect 136146 79744 136174 80036
rect 136238 79966 136266 80036
rect 136330 79966 136358 80036
rect 136226 79960 136278 79966
rect 136226 79902 136278 79908
rect 136318 79960 136370 79966
rect 136318 79902 136370 79908
rect 136422 79830 136450 80036
rect 136514 79937 136542 80036
rect 136606 79966 136634 80036
rect 136594 79960 136646 79966
rect 136500 79928 136556 79937
rect 136594 79902 136646 79908
rect 136500 79863 136556 79872
rect 136410 79824 136462 79830
rect 136410 79766 136462 79772
rect 136698 79744 136726 80036
rect 136790 79937 136818 80036
rect 136776 79928 136832 79937
rect 136776 79863 136832 79872
rect 136882 79778 136910 80036
rect 136974 79966 137002 80036
rect 137066 79966 137094 80036
rect 137158 79971 137186 80036
rect 136962 79960 137014 79966
rect 136962 79902 137014 79908
rect 137054 79960 137106 79966
rect 137054 79902 137106 79908
rect 137144 79962 137200 79971
rect 137250 79966 137278 80036
rect 137144 79897 137200 79906
rect 137238 79960 137290 79966
rect 137342 79937 137370 80036
rect 137238 79902 137290 79908
rect 137328 79928 137384 79937
rect 137434 79898 137462 80036
rect 137526 79966 137554 80036
rect 137514 79960 137566 79966
rect 137514 79902 137566 79908
rect 137328 79863 137384 79872
rect 137422 79892 137474 79898
rect 136836 79762 136910 79778
rect 136146 79716 136312 79744
rect 135718 79656 135774 79665
rect 135456 79580 135530 79608
rect 135628 79620 135680 79626
rect 135456 77761 135484 79580
rect 135718 79591 135774 79600
rect 135628 79562 135680 79568
rect 135534 79520 135590 79529
rect 135534 79455 135536 79464
rect 135588 79455 135590 79464
rect 135536 79426 135588 79432
rect 135442 77752 135498 77761
rect 135442 77687 135498 77696
rect 135640 77636 135668 79562
rect 135718 79520 135774 79529
rect 135718 79455 135720 79464
rect 135772 79455 135774 79464
rect 135720 79426 135772 79432
rect 135350 77616 135406 77625
rect 135350 77551 135406 77560
rect 135456 77608 135668 77636
rect 135364 77042 135392 77551
rect 135352 77036 135404 77042
rect 135352 76978 135404 76984
rect 135350 76664 135406 76673
rect 135350 76599 135352 76608
rect 135404 76599 135406 76608
rect 135352 76570 135404 76576
rect 135456 75682 135484 77608
rect 135732 77568 135760 79426
rect 135548 77540 135760 77568
rect 135444 75676 135496 75682
rect 135444 75618 135496 75624
rect 135444 74996 135496 75002
rect 135444 74938 135496 74944
rect 135260 72820 135312 72826
rect 135260 72762 135312 72768
rect 135272 72350 135300 72762
rect 135260 72344 135312 72350
rect 135260 72286 135312 72292
rect 134720 70366 134932 70394
rect 134720 69834 134748 70366
rect 134708 69828 134760 69834
rect 134708 69770 134760 69776
rect 135456 69018 135484 74938
rect 135548 72486 135576 77540
rect 135824 77489 135852 79716
rect 135996 79688 136048 79694
rect 135902 79656 135958 79665
rect 135996 79630 136048 79636
rect 135902 79591 135958 79600
rect 135810 77480 135866 77489
rect 135810 77415 135866 77424
rect 135628 77036 135680 77042
rect 135628 76978 135680 76984
rect 135536 72480 135588 72486
rect 135536 72422 135588 72428
rect 135536 72344 135588 72350
rect 135536 72286 135588 72292
rect 135444 69012 135496 69018
rect 135444 68954 135496 68960
rect 135444 67516 135496 67522
rect 135444 67458 135496 67464
rect 135260 61260 135312 61266
rect 135260 61202 135312 61208
rect 134524 4004 134576 4010
rect 134524 3946 134576 3952
rect 135272 3602 135300 61202
rect 135352 37324 135404 37330
rect 135352 37266 135404 37272
rect 135260 3596 135312 3602
rect 135260 3538 135312 3544
rect 134156 3528 134208 3534
rect 135364 3482 135392 37266
rect 135456 35222 135484 67458
rect 135444 35216 135496 35222
rect 135444 35158 135496 35164
rect 135548 31074 135576 72286
rect 135640 37942 135668 76978
rect 135916 75914 135944 79591
rect 136008 78577 136036 79630
rect 136180 79620 136232 79626
rect 136180 79562 136232 79568
rect 136088 79552 136140 79558
rect 136088 79494 136140 79500
rect 135994 78568 136050 78577
rect 135994 78503 136050 78512
rect 135996 77852 136048 77858
rect 135996 77794 136048 77800
rect 135732 75886 135944 75914
rect 135732 61402 135760 75886
rect 135812 75200 135864 75206
rect 135812 75142 135864 75148
rect 135824 67522 135852 75142
rect 135812 67516 135864 67522
rect 135812 67458 135864 67464
rect 136008 62082 136036 77794
rect 136100 77790 136128 79494
rect 136192 78470 136220 79562
rect 136180 78464 136232 78470
rect 136180 78406 136232 78412
rect 136088 77784 136140 77790
rect 136088 77726 136140 77732
rect 136284 75002 136312 79716
rect 136652 79716 136726 79744
rect 136824 79756 136910 79762
rect 136456 79688 136508 79694
rect 136456 79630 136508 79636
rect 136364 79620 136416 79626
rect 136364 79562 136416 79568
rect 136272 74996 136324 75002
rect 136272 74938 136324 74944
rect 136376 73642 136404 79562
rect 136468 77858 136496 79630
rect 136548 79620 136600 79626
rect 136548 79562 136600 79568
rect 136456 77852 136508 77858
rect 136456 77794 136508 77800
rect 136456 75676 136508 75682
rect 136456 75618 136508 75624
rect 136364 73636 136416 73642
rect 136364 73578 136416 73584
rect 136468 70394 136496 75618
rect 136560 75206 136588 79562
rect 136652 75206 136680 79716
rect 136876 79750 136910 79756
rect 137342 79744 137370 79863
rect 137422 79834 137474 79840
rect 136824 79698 136876 79704
rect 137204 79716 137370 79744
rect 137468 79756 137520 79762
rect 136916 79688 136968 79694
rect 136730 79656 136786 79665
rect 137100 79688 137152 79694
rect 136916 79630 136968 79636
rect 137006 79656 137062 79665
rect 136730 79591 136786 79600
rect 136548 75200 136600 75206
rect 136548 75142 136600 75148
rect 136640 75200 136692 75206
rect 136640 75142 136692 75148
rect 136744 71774 136772 79591
rect 136824 77852 136876 77858
rect 136824 77794 136876 77800
rect 136652 71746 136772 71774
rect 136468 70366 136588 70394
rect 136560 70038 136588 70366
rect 136548 70032 136600 70038
rect 136548 69974 136600 69980
rect 135996 62076 136048 62082
rect 135996 62018 136048 62024
rect 135720 61396 135772 61402
rect 135720 61338 135772 61344
rect 136652 44878 136680 71746
rect 136836 55962 136864 77794
rect 136928 76906 136956 79630
rect 137100 79630 137152 79636
rect 137006 79591 137008 79600
rect 137060 79591 137062 79600
rect 137008 79562 137060 79568
rect 137006 79520 137062 79529
rect 137006 79455 137008 79464
rect 137060 79455 137062 79464
rect 137008 79426 137060 79432
rect 136916 76900 136968 76906
rect 136916 76842 136968 76848
rect 136916 71052 136968 71058
rect 136916 70994 136968 71000
rect 136824 55956 136876 55962
rect 136824 55898 136876 55904
rect 136640 44872 136692 44878
rect 136640 44814 136692 44820
rect 135628 37936 135680 37942
rect 135628 37878 135680 37884
rect 135536 31068 135588 31074
rect 135536 31010 135588 31016
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 134156 3470 134208 3476
rect 132960 3392 133012 3398
rect 132960 3334 133012 3340
rect 131764 3324 131816 3330
rect 131764 3266 131816 3272
rect 132972 480 133000 3334
rect 134168 480 134196 3470
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3538
rect 136928 3534 136956 70994
rect 137112 64870 137140 79630
rect 137204 77858 137232 79716
rect 137468 79698 137520 79704
rect 137374 79656 137430 79665
rect 137284 79620 137336 79626
rect 137374 79591 137430 79600
rect 137284 79562 137336 79568
rect 137296 78062 137324 79562
rect 137284 78056 137336 78062
rect 137284 77998 137336 78004
rect 137192 77852 137244 77858
rect 137192 77794 137244 77800
rect 137388 75914 137416 79591
rect 137480 77178 137508 79698
rect 137618 79676 137646 80036
rect 137710 79744 137738 80036
rect 137802 79898 137830 80036
rect 137790 79892 137842 79898
rect 137790 79834 137842 79840
rect 137894 79778 137922 80036
rect 137986 79937 138014 80036
rect 137972 79928 138028 79937
rect 137972 79863 138028 79872
rect 138078 79778 138106 80036
rect 137894 79750 137968 79778
rect 137710 79716 137784 79744
rect 137618 79648 137692 79676
rect 137664 79529 137692 79648
rect 137650 79520 137706 79529
rect 137650 79455 137706 79464
rect 137468 77172 137520 77178
rect 137468 77114 137520 77120
rect 137296 75886 137416 75914
rect 137192 75200 137244 75206
rect 137192 75142 137244 75148
rect 137204 66230 137232 75142
rect 137296 66910 137324 75886
rect 137664 74934 137692 79455
rect 137756 78810 137784 79716
rect 137836 79688 137888 79694
rect 137836 79630 137888 79636
rect 137744 78804 137796 78810
rect 137744 78746 137796 78752
rect 137848 78112 137876 79630
rect 137940 79490 137968 79750
rect 138032 79750 138106 79778
rect 138170 79778 138198 80036
rect 138262 79966 138290 80036
rect 138250 79960 138302 79966
rect 138250 79902 138302 79908
rect 138354 79778 138382 80036
rect 138446 79971 138474 80036
rect 138432 79962 138488 79971
rect 138432 79897 138488 79906
rect 138538 79801 138566 80036
rect 138170 79750 138244 79778
rect 137928 79484 137980 79490
rect 137928 79426 137980 79432
rect 137756 78084 137876 78112
rect 137652 74928 137704 74934
rect 137652 74870 137704 74876
rect 137756 69014 137784 78084
rect 137834 78024 137890 78033
rect 137834 77959 137890 77968
rect 137848 77790 137876 77959
rect 137836 77784 137888 77790
rect 137836 77726 137888 77732
rect 137940 72622 137968 79426
rect 138032 77217 138060 79750
rect 138112 79688 138164 79694
rect 138112 79630 138164 79636
rect 138124 77761 138152 79630
rect 138216 77897 138244 79750
rect 138308 79750 138382 79778
rect 138524 79792 138580 79801
rect 138202 77888 138258 77897
rect 138202 77823 138258 77832
rect 138110 77752 138166 77761
rect 138110 77687 138166 77696
rect 138018 77208 138074 77217
rect 138018 77143 138074 77152
rect 138308 76498 138336 79750
rect 138524 79727 138580 79736
rect 138388 79688 138440 79694
rect 138480 79688 138532 79694
rect 138388 79630 138440 79636
rect 138478 79656 138480 79665
rect 138532 79656 138534 79665
rect 138296 76492 138348 76498
rect 138296 76434 138348 76440
rect 138400 73846 138428 79630
rect 138478 79591 138534 79600
rect 138492 78742 138520 79591
rect 138630 79540 138658 80036
rect 138722 79971 138750 80036
rect 138708 79962 138764 79971
rect 138708 79897 138764 79906
rect 138814 79812 138842 80036
rect 138906 79966 138934 80036
rect 138894 79960 138946 79966
rect 138894 79902 138946 79908
rect 138998 79898 139026 80036
rect 139090 79966 139118 80036
rect 139078 79960 139130 79966
rect 139078 79902 139130 79908
rect 138986 79892 139038 79898
rect 138986 79834 139038 79840
rect 138722 79784 138842 79812
rect 138722 79676 138750 79784
rect 139182 79744 139210 80036
rect 139274 79937 139302 80036
rect 139260 79928 139316 79937
rect 139260 79863 139316 79872
rect 139366 79812 139394 80036
rect 139458 79966 139486 80036
rect 139446 79960 139498 79966
rect 139446 79902 139498 79908
rect 139366 79784 139440 79812
rect 139550 79801 139578 80036
rect 139642 79966 139670 80036
rect 139734 79966 139762 80036
rect 139630 79960 139682 79966
rect 139630 79902 139682 79908
rect 139722 79960 139774 79966
rect 139722 79902 139774 79908
rect 139826 79898 139854 80036
rect 139814 79892 139866 79898
rect 139814 79834 139866 79840
rect 139182 79716 139348 79744
rect 138722 79648 138796 79676
rect 138584 79512 138658 79540
rect 138480 78736 138532 78742
rect 138480 78678 138532 78684
rect 138584 73982 138612 79512
rect 138768 78674 138796 79648
rect 139214 79656 139270 79665
rect 139214 79591 139270 79600
rect 138756 78668 138808 78674
rect 138756 78610 138808 78616
rect 139032 78668 139084 78674
rect 139032 78610 139084 78616
rect 138662 78432 138718 78441
rect 138662 78367 138718 78376
rect 138676 75274 138704 78367
rect 138754 77888 138810 77897
rect 138754 77823 138810 77832
rect 138768 77353 138796 77823
rect 138754 77344 138810 77353
rect 138754 77279 138810 77288
rect 138664 75268 138716 75274
rect 138664 75210 138716 75216
rect 138572 73976 138624 73982
rect 138572 73918 138624 73924
rect 138388 73840 138440 73846
rect 138388 73782 138440 73788
rect 137928 72616 137980 72622
rect 137928 72558 137980 72564
rect 138572 71596 138624 71602
rect 138572 71538 138624 71544
rect 138388 71256 138440 71262
rect 138388 71198 138440 71204
rect 138400 70258 138428 71198
rect 138584 71126 138612 71538
rect 139044 71262 139072 78610
rect 139124 78056 139176 78062
rect 139124 77998 139176 78004
rect 139136 75614 139164 77998
rect 139124 75608 139176 75614
rect 139124 75550 139176 75556
rect 139032 71256 139084 71262
rect 139032 71198 139084 71204
rect 138572 71120 138624 71126
rect 138572 71062 138624 71068
rect 137388 68986 137784 69014
rect 138124 70230 138428 70258
rect 137284 66904 137336 66910
rect 137284 66846 137336 66852
rect 137192 66224 137244 66230
rect 137192 66166 137244 66172
rect 137100 64864 137152 64870
rect 137100 64806 137152 64812
rect 137388 60586 137416 68986
rect 137376 60580 137428 60586
rect 137376 60522 137428 60528
rect 138020 41676 138072 41682
rect 138020 41618 138072 41624
rect 137652 3596 137704 3602
rect 137652 3538 137704 3544
rect 136916 3528 136968 3534
rect 136916 3470 136968 3476
rect 137664 480 137692 3538
rect 138032 3482 138060 41618
rect 138124 3670 138152 70230
rect 138584 64874 138612 71062
rect 138216 64846 138612 64874
rect 138216 8974 138244 64846
rect 139228 62898 139256 79591
rect 139320 71602 139348 79716
rect 139412 78062 139440 79784
rect 139536 79792 139592 79801
rect 139918 79744 139946 80036
rect 140010 79812 140038 80036
rect 140102 79937 140130 80036
rect 140088 79928 140144 79937
rect 140194 79898 140222 80036
rect 140088 79863 140144 79872
rect 140182 79892 140234 79898
rect 140182 79834 140234 79840
rect 140010 79784 140084 79812
rect 139536 79727 139592 79736
rect 139872 79716 139946 79744
rect 139492 79688 139544 79694
rect 139492 79630 139544 79636
rect 139400 78056 139452 78062
rect 139400 77998 139452 78004
rect 139504 77761 139532 79630
rect 139584 79620 139636 79626
rect 139584 79562 139636 79568
rect 139490 77752 139546 77761
rect 139490 77687 139546 77696
rect 139596 77625 139624 79562
rect 139768 79552 139820 79558
rect 139768 79494 139820 79500
rect 139676 78804 139728 78810
rect 139676 78746 139728 78752
rect 139582 77616 139638 77625
rect 139582 77551 139638 77560
rect 139688 75750 139716 78746
rect 139780 78656 139808 79494
rect 139872 78810 139900 79716
rect 140056 79642 140084 79784
rect 140134 79792 140190 79801
rect 140286 79778 140314 80036
rect 140378 79971 140406 80036
rect 140364 79962 140420 79971
rect 140364 79897 140420 79906
rect 140470 79898 140498 80036
rect 140562 79971 140590 80036
rect 140548 79962 140604 79971
rect 140654 79966 140682 80036
rect 140134 79727 140190 79736
rect 140240 79750 140314 79778
rect 140378 79778 140406 79897
rect 140458 79892 140510 79898
rect 140548 79897 140604 79906
rect 140642 79960 140694 79966
rect 140642 79902 140694 79908
rect 140458 79834 140510 79840
rect 140596 79824 140648 79830
rect 140594 79792 140596 79801
rect 140648 79792 140650 79801
rect 140378 79750 140452 79778
rect 139964 79614 140084 79642
rect 139860 78804 139912 78810
rect 139860 78746 139912 78752
rect 139780 78628 139900 78656
rect 139768 78532 139820 78538
rect 139768 78474 139820 78480
rect 139676 75744 139728 75750
rect 139676 75686 139728 75692
rect 139584 73160 139636 73166
rect 139584 73102 139636 73108
rect 139308 71596 139360 71602
rect 139308 71538 139360 71544
rect 139400 64932 139452 64938
rect 139400 64874 139452 64880
rect 139216 62892 139268 62898
rect 139216 62834 139268 62840
rect 138664 55276 138716 55282
rect 138664 55218 138716 55224
rect 138204 8968 138256 8974
rect 138204 8910 138256 8916
rect 138112 3664 138164 3670
rect 138112 3606 138164 3612
rect 138676 3602 138704 55218
rect 139412 6914 139440 64874
rect 139596 10334 139624 73102
rect 139780 54534 139808 78474
rect 139872 66026 139900 78628
rect 139964 66162 139992 79614
rect 140044 79552 140096 79558
rect 140044 79494 140096 79500
rect 140056 79393 140084 79494
rect 140042 79384 140098 79393
rect 140042 79319 140098 79328
rect 140056 73914 140084 79319
rect 140148 78538 140176 79727
rect 140240 79665 140268 79750
rect 140320 79688 140372 79694
rect 140226 79656 140282 79665
rect 140320 79630 140372 79636
rect 140226 79591 140282 79600
rect 140332 79506 140360 79630
rect 140240 79478 140360 79506
rect 140136 78532 140188 78538
rect 140136 78474 140188 78480
rect 140044 73908 140096 73914
rect 140044 73850 140096 73856
rect 140240 70174 140268 79478
rect 140424 79404 140452 79750
rect 140746 79744 140774 80036
rect 140838 79966 140866 80036
rect 140826 79960 140878 79966
rect 140826 79902 140878 79908
rect 140594 79727 140650 79736
rect 140502 79656 140558 79665
rect 140502 79591 140558 79600
rect 140332 79376 140452 79404
rect 140228 70168 140280 70174
rect 140228 70110 140280 70116
rect 139952 66156 140004 66162
rect 139952 66098 140004 66104
rect 139860 66020 139912 66026
rect 139860 65962 139912 65968
rect 139768 54528 139820 54534
rect 139768 54470 139820 54476
rect 139584 10328 139636 10334
rect 139584 10270 139636 10276
rect 139412 6886 139624 6914
rect 138664 3596 138716 3602
rect 138664 3538 138716 3544
rect 138032 3454 138888 3482
rect 138860 480 138888 3454
rect 131734 354 131846 480
rect 131132 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 6886
rect 140332 6186 140360 79376
rect 140516 73166 140544 79591
rect 140608 76362 140636 79727
rect 140700 79716 140774 79744
rect 140930 79744 140958 80036
rect 141022 79966 141050 80036
rect 141010 79960 141062 79966
rect 141010 79902 141062 79908
rect 141114 79778 141142 80036
rect 141206 79966 141234 80036
rect 141194 79960 141246 79966
rect 141194 79902 141246 79908
rect 141298 79898 141326 80036
rect 141286 79892 141338 79898
rect 141286 79834 141338 79840
rect 141068 79762 141142 79778
rect 141056 79756 141142 79762
rect 140930 79716 141004 79744
rect 140596 76356 140648 76362
rect 140596 76298 140648 76304
rect 140700 74322 140728 79716
rect 140780 79620 140832 79626
rect 140780 79562 140832 79568
rect 140792 78577 140820 79562
rect 140870 79384 140926 79393
rect 140870 79319 140926 79328
rect 140778 78568 140834 78577
rect 140778 78503 140834 78512
rect 140688 74316 140740 74322
rect 140688 74258 140740 74264
rect 140504 73160 140556 73166
rect 140504 73102 140556 73108
rect 140780 66292 140832 66298
rect 140780 66234 140832 66240
rect 140320 6180 140372 6186
rect 140320 6122 140372 6128
rect 140792 1306 140820 66234
rect 140884 3874 140912 79319
rect 140976 77625 141004 79716
rect 141108 79750 141142 79756
rect 141056 79698 141108 79704
rect 141148 79688 141200 79694
rect 141390 79676 141418 80036
rect 141482 79898 141510 80036
rect 141574 79966 141602 80036
rect 141562 79960 141614 79966
rect 141562 79902 141614 79908
rect 141666 79898 141694 80036
rect 141470 79892 141522 79898
rect 141470 79834 141522 79840
rect 141654 79892 141706 79898
rect 141654 79834 141706 79840
rect 141758 79801 141786 80036
rect 141850 79966 141878 80036
rect 141838 79960 141890 79966
rect 141838 79902 141890 79908
rect 141942 79812 141970 80036
rect 142034 79937 142062 80036
rect 142020 79928 142076 79937
rect 142020 79863 142076 79872
rect 141744 79792 141800 79801
rect 141896 79784 141970 79812
rect 141800 79736 141832 79744
rect 141744 79727 141832 79736
rect 141758 79716 141832 79727
rect 141390 79648 141464 79676
rect 141148 79630 141200 79636
rect 141056 79620 141108 79626
rect 141056 79562 141108 79568
rect 141068 78198 141096 79562
rect 141160 79422 141188 79630
rect 141240 79552 141292 79558
rect 141240 79494 141292 79500
rect 141332 79552 141384 79558
rect 141332 79494 141384 79500
rect 141148 79416 141200 79422
rect 141148 79358 141200 79364
rect 141056 78192 141108 78198
rect 141056 78134 141108 78140
rect 141054 77752 141110 77761
rect 141054 77687 141110 77696
rect 140962 77616 141018 77625
rect 140962 77551 141018 77560
rect 140964 77512 141016 77518
rect 140964 77454 141016 77460
rect 140976 66978 141004 77454
rect 141068 76770 141096 77687
rect 141056 76764 141108 76770
rect 141056 76706 141108 76712
rect 141160 70394 141188 79358
rect 141252 76945 141280 79494
rect 141344 79393 141372 79494
rect 141330 79384 141386 79393
rect 141330 79319 141386 79328
rect 141344 77518 141372 79319
rect 141332 77512 141384 77518
rect 141332 77454 141384 77460
rect 141238 76936 141294 76945
rect 141436 76888 141464 79648
rect 141516 79484 141568 79490
rect 141516 79426 141568 79432
rect 141238 76871 141294 76880
rect 141344 76860 141464 76888
rect 141344 75138 141372 76860
rect 141424 76764 141476 76770
rect 141424 76706 141476 76712
rect 141332 75132 141384 75138
rect 141332 75074 141384 75080
rect 141068 70366 141188 70394
rect 141068 67046 141096 70366
rect 141056 67040 141108 67046
rect 141056 66982 141108 66988
rect 140964 66972 141016 66978
rect 140964 66914 141016 66920
rect 140872 3868 140924 3874
rect 140872 3810 140924 3816
rect 141436 3602 141464 76706
rect 141528 72418 141556 79426
rect 141608 79416 141660 79422
rect 141606 79384 141608 79393
rect 141660 79384 141662 79393
rect 141606 79319 141662 79328
rect 141700 79008 141752 79014
rect 141700 78950 141752 78956
rect 141712 78810 141740 78950
rect 141700 78804 141752 78810
rect 141700 78746 141752 78752
rect 141700 78192 141752 78198
rect 141700 78134 141752 78140
rect 141712 77722 141740 78134
rect 141700 77716 141752 77722
rect 141700 77658 141752 77664
rect 141608 73976 141660 73982
rect 141608 73918 141660 73924
rect 141516 72412 141568 72418
rect 141516 72354 141568 72360
rect 141516 71596 141568 71602
rect 141516 71538 141568 71544
rect 141424 3596 141476 3602
rect 141424 3538 141476 3544
rect 141528 3398 141556 71538
rect 141620 69630 141648 73918
rect 141804 70394 141832 79716
rect 141896 78470 141924 79784
rect 141976 79688 142028 79694
rect 142126 79676 142154 80036
rect 142218 79830 142246 80036
rect 142206 79824 142258 79830
rect 142206 79766 142258 79772
rect 142310 79744 142338 80036
rect 142402 79966 142430 80036
rect 142390 79960 142442 79966
rect 142390 79902 142442 79908
rect 142494 79898 142522 80036
rect 142482 79892 142534 79898
rect 142482 79834 142534 79840
rect 142586 79744 142614 80036
rect 142678 79971 142706 80036
rect 142664 79962 142720 79971
rect 142664 79897 142720 79906
rect 142770 79830 142798 80036
rect 142758 79824 142810 79830
rect 142862 79801 142890 80036
rect 142954 79898 142982 80036
rect 143046 79971 143074 80036
rect 143032 79962 143088 79971
rect 142942 79892 142994 79898
rect 143032 79897 143088 79906
rect 142942 79834 142994 79840
rect 142758 79766 142810 79772
rect 142848 79792 142904 79801
rect 142310 79716 142384 79744
rect 142126 79648 142200 79676
rect 141976 79630 142028 79636
rect 141884 78464 141936 78470
rect 141884 78406 141936 78412
rect 141988 73982 142016 79630
rect 142068 79552 142120 79558
rect 142068 79494 142120 79500
rect 141976 73976 142028 73982
rect 141976 73918 142028 73924
rect 142080 70990 142108 79494
rect 142172 74730 142200 79648
rect 142356 78606 142384 79716
rect 142540 79716 142614 79744
rect 143138 79778 143166 80036
rect 143230 79898 143258 80036
rect 143218 79892 143270 79898
rect 143218 79834 143270 79840
rect 143138 79750 143212 79778
rect 142848 79727 142904 79736
rect 142540 79608 142568 79716
rect 143184 79665 143212 79750
rect 143322 79744 143350 80036
rect 143414 79966 143442 80036
rect 143402 79960 143454 79966
rect 143402 79902 143454 79908
rect 143506 79898 143534 80036
rect 143598 79966 143626 80036
rect 143586 79960 143638 79966
rect 143586 79902 143638 79908
rect 143690 79898 143718 80036
rect 143782 79937 143810 80036
rect 143768 79928 143824 79937
rect 143494 79892 143546 79898
rect 143494 79834 143546 79840
rect 143678 79892 143730 79898
rect 143768 79863 143824 79872
rect 143678 79834 143730 79840
rect 143630 79792 143686 79801
rect 143540 79756 143592 79762
rect 143322 79716 143396 79744
rect 142710 79656 142766 79665
rect 142448 79580 142568 79608
rect 142620 79620 142672 79626
rect 142344 78600 142396 78606
rect 142344 78542 142396 78548
rect 142448 77994 142476 79580
rect 143170 79656 143226 79665
rect 142710 79591 142766 79600
rect 142804 79620 142856 79626
rect 142620 79562 142672 79568
rect 142528 79484 142580 79490
rect 142528 79426 142580 79432
rect 142436 77988 142488 77994
rect 142436 77930 142488 77936
rect 142436 77852 142488 77858
rect 142436 77794 142488 77800
rect 142160 74724 142212 74730
rect 142160 74666 142212 74672
rect 142448 74050 142476 77794
rect 142436 74044 142488 74050
rect 142436 73986 142488 73992
rect 142252 73092 142304 73098
rect 142252 73034 142304 73040
rect 142264 72690 142292 73034
rect 142252 72684 142304 72690
rect 142252 72626 142304 72632
rect 142068 70984 142120 70990
rect 142068 70926 142120 70932
rect 142066 70408 142122 70417
rect 141804 70366 142016 70394
rect 141608 69624 141660 69630
rect 141608 69566 141660 69572
rect 141988 67114 142016 70366
rect 142066 70343 142122 70352
rect 141976 67108 142028 67114
rect 141976 67050 142028 67056
rect 142080 67017 142108 70343
rect 142160 69692 142212 69698
rect 142160 69634 142212 69640
rect 142066 67008 142122 67017
rect 142066 66943 142122 66952
rect 142172 66298 142200 69634
rect 142160 66292 142212 66298
rect 142160 66234 142212 66240
rect 142264 65006 142292 72626
rect 142344 71460 142396 71466
rect 142344 71402 142396 71408
rect 142356 71194 142384 71402
rect 142344 71188 142396 71194
rect 142344 71130 142396 71136
rect 142252 65000 142304 65006
rect 142252 64942 142304 64948
rect 142356 64874 142384 71130
rect 142448 70922 142476 73986
rect 142540 72554 142568 79426
rect 142632 77926 142660 79562
rect 142620 77920 142672 77926
rect 142620 77862 142672 77868
rect 142724 76888 142752 79591
rect 143368 79608 143396 79716
rect 143874 79778 143902 80036
rect 143966 79830 143994 80036
rect 143630 79727 143686 79736
rect 143736 79750 143902 79778
rect 143954 79824 144006 79830
rect 143954 79766 144006 79772
rect 144058 79778 144086 80036
rect 144150 79898 144178 80036
rect 144138 79892 144190 79898
rect 144138 79834 144190 79840
rect 144242 79778 144270 80036
rect 144058 79750 144132 79778
rect 143540 79698 143592 79704
rect 143170 79591 143226 79600
rect 142804 79562 142856 79568
rect 143276 79580 143396 79608
rect 142632 76860 142752 76888
rect 142528 72548 142580 72554
rect 142528 72490 142580 72496
rect 142436 70916 142488 70922
rect 142436 70858 142488 70864
rect 142436 69896 142488 69902
rect 142436 69838 142488 69844
rect 142264 64846 142384 64874
rect 142264 55282 142292 64846
rect 142252 55276 142304 55282
rect 142252 55218 142304 55224
rect 142448 37330 142476 69838
rect 142540 61266 142568 72490
rect 142632 69970 142660 76860
rect 142710 75984 142766 75993
rect 142710 75919 142766 75928
rect 142620 69964 142672 69970
rect 142620 69906 142672 69912
rect 142528 61260 142580 61266
rect 142528 61202 142580 61208
rect 142632 41682 142660 69906
rect 142724 69902 142752 75919
rect 142816 71058 142844 79562
rect 142896 79552 142948 79558
rect 142896 79494 142948 79500
rect 142908 78198 142936 79494
rect 143172 79484 143224 79490
rect 143172 79426 143224 79432
rect 142896 78192 142948 78198
rect 142896 78134 142948 78140
rect 142988 77920 143040 77926
rect 142988 77862 143040 77868
rect 142894 76664 142950 76673
rect 142894 76599 142950 76608
rect 142908 72758 142936 76599
rect 142896 72752 142948 72758
rect 142896 72694 142948 72700
rect 142908 71602 142936 72694
rect 142896 71596 142948 71602
rect 142896 71538 142948 71544
rect 143000 71482 143028 77862
rect 143184 76770 143212 79426
rect 143172 76764 143224 76770
rect 143172 76706 143224 76712
rect 143170 75984 143226 75993
rect 143170 75919 143226 75928
rect 142908 71454 143028 71482
rect 143184 71466 143212 75919
rect 143172 71460 143224 71466
rect 142804 71052 142856 71058
rect 142804 70994 142856 71000
rect 142804 70916 142856 70922
rect 142804 70858 142856 70864
rect 142712 69896 142764 69902
rect 142712 69838 142764 69844
rect 142620 41676 142672 41682
rect 142620 41618 142672 41624
rect 142436 37324 142488 37330
rect 142436 37266 142488 37272
rect 142816 9654 142844 70858
rect 142804 9648 142856 9654
rect 142804 9590 142856 9596
rect 142908 6914 142936 71454
rect 143172 71402 143224 71408
rect 143276 70394 143304 79580
rect 143448 79484 143500 79490
rect 143448 79426 143500 79432
rect 143460 77858 143488 79426
rect 143552 78713 143580 79698
rect 143538 78704 143594 78713
rect 143538 78639 143594 78648
rect 143448 77852 143500 77858
rect 143448 77794 143500 77800
rect 143448 76764 143500 76770
rect 143448 76706 143500 76712
rect 143460 73098 143488 76706
rect 143540 74520 143592 74526
rect 143540 74462 143592 74468
rect 143552 73846 143580 74462
rect 143540 73840 143592 73846
rect 143540 73782 143592 73788
rect 143448 73092 143500 73098
rect 143448 73034 143500 73040
rect 143000 70366 143304 70394
rect 143000 69698 143028 70366
rect 142988 69692 143040 69698
rect 142988 69634 143040 69640
rect 143644 19990 143672 79727
rect 143736 77790 143764 79750
rect 143816 79688 143868 79694
rect 143814 79656 143816 79665
rect 144000 79688 144052 79694
rect 143868 79656 143870 79665
rect 144000 79630 144052 79636
rect 143814 79591 143870 79600
rect 143724 77784 143776 77790
rect 143724 77726 143776 77732
rect 143724 74520 143776 74526
rect 143724 74462 143776 74468
rect 143736 74186 143764 74462
rect 143724 74180 143776 74186
rect 143724 74122 143776 74128
rect 143736 69698 143764 74122
rect 143724 69692 143776 69698
rect 143724 69634 143776 69640
rect 143828 52902 143856 79591
rect 144012 67590 144040 79630
rect 144104 74526 144132 79750
rect 144196 79750 144270 79778
rect 144092 74520 144144 74526
rect 144092 74462 144144 74468
rect 144196 73846 144224 79750
rect 144334 79676 144362 80036
rect 144426 79801 144454 80036
rect 144518 79937 144546 80036
rect 144504 79928 144560 79937
rect 144610 79898 144638 80036
rect 144702 79937 144730 80036
rect 144794 79966 144822 80036
rect 144886 79966 144914 80036
rect 144782 79960 144834 79966
rect 144688 79928 144744 79937
rect 144504 79863 144560 79872
rect 144598 79892 144650 79898
rect 144782 79902 144834 79908
rect 144874 79960 144926 79966
rect 144874 79902 144926 79908
rect 144688 79863 144744 79872
rect 144598 79834 144650 79840
rect 144412 79792 144468 79801
rect 144702 79778 144730 79863
rect 144828 79824 144880 79830
rect 144702 79750 144776 79778
rect 144828 79766 144880 79772
rect 144412 79727 144468 79736
rect 144288 79648 144362 79676
rect 144644 79688 144696 79694
rect 144288 74458 144316 79648
rect 144644 79630 144696 79636
rect 144368 79552 144420 79558
rect 144368 79494 144420 79500
rect 144552 79552 144604 79558
rect 144552 79494 144604 79500
rect 144380 78742 144408 79494
rect 144460 79348 144512 79354
rect 144460 79290 144512 79296
rect 144368 78736 144420 78742
rect 144368 78678 144420 78684
rect 144368 77784 144420 77790
rect 144368 77726 144420 77732
rect 144276 74452 144328 74458
rect 144276 74394 144328 74400
rect 144184 73840 144236 73846
rect 144184 73782 144236 73788
rect 144000 67584 144052 67590
rect 144000 67526 144052 67532
rect 144012 64874 144040 67526
rect 144012 64846 144224 64874
rect 143816 52896 143868 52902
rect 143816 52838 143868 52844
rect 144196 47598 144224 64846
rect 144288 59362 144316 74394
rect 144380 66230 144408 77726
rect 144368 66224 144420 66230
rect 144368 66166 144420 66172
rect 144276 59356 144328 59362
rect 144276 59298 144328 59304
rect 144184 47592 144236 47598
rect 144184 47534 144236 47540
rect 144472 40050 144500 79290
rect 144564 78577 144592 79494
rect 144550 78568 144606 78577
rect 144550 78503 144606 78512
rect 144656 74497 144684 79630
rect 144642 74488 144698 74497
rect 144642 74423 144698 74432
rect 144748 70394 144776 79750
rect 144840 79393 144868 79766
rect 144978 79744 145006 80036
rect 144932 79716 145006 79744
rect 145070 79744 145098 80036
rect 145162 79937 145190 80036
rect 145148 79928 145204 79937
rect 145148 79863 145204 79872
rect 145254 79744 145282 80036
rect 145346 79801 145374 80036
rect 145070 79716 145144 79744
rect 144826 79384 144882 79393
rect 144826 79319 144882 79328
rect 144932 77654 144960 79716
rect 145012 79484 145064 79490
rect 145012 79426 145064 79432
rect 145024 79150 145052 79426
rect 145012 79144 145064 79150
rect 145012 79086 145064 79092
rect 144920 77648 144972 77654
rect 144920 77590 144972 77596
rect 145024 77500 145052 79086
rect 144932 77472 145052 77500
rect 144932 70394 144960 77472
rect 145116 75834 145144 79716
rect 145208 79716 145282 79744
rect 145332 79792 145388 79801
rect 145332 79727 145388 79736
rect 145438 79744 145466 80036
rect 145530 79898 145558 80036
rect 145518 79892 145570 79898
rect 145518 79834 145570 79840
rect 145622 79778 145650 80036
rect 145714 79966 145742 80036
rect 145806 79966 145834 80036
rect 145702 79960 145754 79966
rect 145702 79902 145754 79908
rect 145794 79960 145846 79966
rect 145794 79902 145846 79908
rect 145898 79812 145926 80036
rect 145990 79966 146018 80036
rect 146082 79966 146110 80036
rect 146174 79971 146202 80036
rect 145978 79960 146030 79966
rect 145978 79902 146030 79908
rect 146070 79960 146122 79966
rect 146070 79902 146122 79908
rect 146160 79962 146216 79971
rect 146266 79966 146294 80036
rect 146160 79897 146216 79906
rect 146254 79960 146306 79966
rect 146254 79902 146306 79908
rect 146358 79898 146386 80036
rect 146346 79892 146398 79898
rect 146346 79834 146398 79840
rect 146024 79824 146076 79830
rect 145898 79784 145972 79812
rect 145576 79762 145650 79778
rect 145564 79756 145650 79762
rect 145438 79716 145512 79744
rect 145208 79642 145236 79716
rect 145378 79656 145434 79665
rect 145208 79614 145328 79642
rect 145196 79552 145248 79558
rect 145196 79494 145248 79500
rect 145024 75806 145144 75834
rect 145024 74526 145052 75806
rect 145012 74520 145064 74526
rect 145012 74462 145064 74468
rect 145024 74254 145052 74462
rect 145012 74248 145064 74254
rect 145012 74190 145064 74196
rect 144748 70366 144868 70394
rect 144932 70366 145144 70394
rect 144460 40044 144512 40050
rect 144460 39986 144512 39992
rect 143632 19984 143684 19990
rect 143632 19926 143684 19932
rect 143540 9648 143592 9654
rect 143540 9590 143592 9596
rect 142448 6886 142936 6914
rect 141516 3392 141568 3398
rect 141516 3334 141568 3340
rect 140792 1278 141280 1306
rect 141252 480 141280 1278
rect 142448 480 142476 6886
rect 143552 480 143580 9590
rect 144840 4826 144868 70366
rect 145116 64874 145144 70366
rect 145024 64846 145144 64874
rect 145024 25566 145052 64846
rect 145208 46238 145236 79494
rect 145300 79393 145328 79614
rect 145378 79591 145434 79600
rect 145286 79384 145342 79393
rect 145286 79319 145342 79328
rect 145300 76906 145328 79319
rect 145288 76900 145340 76906
rect 145288 76842 145340 76848
rect 145392 75546 145420 79591
rect 145484 76514 145512 79716
rect 145616 79750 145650 79756
rect 145564 79698 145616 79704
rect 145656 79688 145708 79694
rect 145708 79648 145788 79676
rect 145656 79630 145708 79636
rect 145656 79552 145708 79558
rect 145656 79494 145708 79500
rect 145668 77353 145696 79494
rect 145654 77344 145710 77353
rect 145654 77279 145710 77288
rect 145484 76486 145604 76514
rect 145472 76356 145524 76362
rect 145472 76298 145524 76304
rect 145484 75886 145512 76298
rect 145472 75880 145524 75886
rect 145472 75822 145524 75828
rect 145380 75540 145432 75546
rect 145380 75482 145432 75488
rect 145392 75274 145420 75482
rect 145380 75268 145432 75274
rect 145380 75210 145432 75216
rect 145380 74520 145432 74526
rect 145380 74462 145432 74468
rect 145392 69018 145420 74462
rect 145484 70394 145512 75822
rect 145576 75342 145604 76486
rect 145564 75336 145616 75342
rect 145564 75278 145616 75284
rect 145576 72298 145604 75278
rect 145668 72486 145696 77279
rect 145760 76809 145788 79648
rect 145746 76800 145802 76809
rect 145746 76735 145802 76744
rect 145944 76362 145972 79784
rect 146024 79766 146076 79772
rect 146116 79824 146168 79830
rect 146116 79766 146168 79772
rect 146206 79792 146262 79801
rect 145932 76356 145984 76362
rect 145932 76298 145984 76304
rect 146036 76265 146064 79766
rect 146128 78130 146156 79766
rect 146206 79727 146262 79736
rect 146300 79756 146352 79762
rect 146220 79257 146248 79727
rect 146300 79698 146352 79704
rect 146206 79248 146262 79257
rect 146206 79183 146262 79192
rect 146116 78124 146168 78130
rect 146116 78066 146168 78072
rect 146128 77518 146156 78066
rect 146116 77512 146168 77518
rect 146116 77454 146168 77460
rect 146220 77364 146248 79183
rect 146312 79082 146340 79698
rect 146450 79642 146478 80036
rect 146542 79898 146570 80036
rect 146634 79903 146662 80036
rect 146726 79966 146754 80036
rect 146714 79960 146766 79966
rect 146530 79892 146582 79898
rect 146530 79834 146582 79840
rect 146620 79894 146676 79903
rect 146714 79902 146766 79908
rect 146620 79829 146676 79838
rect 146668 79756 146720 79762
rect 146668 79698 146720 79704
rect 146404 79614 146478 79642
rect 146576 79620 146628 79626
rect 146300 79076 146352 79082
rect 146300 79018 146352 79024
rect 146312 78946 146340 79018
rect 146300 78940 146352 78946
rect 146300 78882 146352 78888
rect 146404 78690 146432 79614
rect 146576 79562 146628 79568
rect 146128 77336 146248 77364
rect 146312 78662 146432 78690
rect 146022 76256 146078 76265
rect 146022 76191 146078 76200
rect 145748 75268 145800 75274
rect 145748 75210 145800 75216
rect 145656 72480 145708 72486
rect 145656 72422 145708 72428
rect 145576 72270 145696 72298
rect 145484 70366 145604 70394
rect 145380 69012 145432 69018
rect 145380 68954 145432 68960
rect 145196 46232 145248 46238
rect 145196 46174 145248 46180
rect 145104 40044 145156 40050
rect 145104 39986 145156 39992
rect 145012 25560 145064 25566
rect 145012 25502 145064 25508
rect 145116 16574 145144 39986
rect 145576 36582 145604 70366
rect 145668 39370 145696 72270
rect 145760 55894 145788 75210
rect 145748 55888 145800 55894
rect 145748 55830 145800 55836
rect 146128 43654 146156 77336
rect 146312 77246 146340 78662
rect 146390 78568 146446 78577
rect 146390 78503 146446 78512
rect 146300 77240 146352 77246
rect 146300 77182 146352 77188
rect 146208 76900 146260 76906
rect 146208 76842 146260 76848
rect 146116 43648 146168 43654
rect 146116 43590 146168 43596
rect 145656 39364 145708 39370
rect 145656 39306 145708 39312
rect 145564 36576 145616 36582
rect 145564 36518 145616 36524
rect 146220 17270 146248 76842
rect 146312 75750 146340 77182
rect 146300 75744 146352 75750
rect 146300 75686 146352 75692
rect 146404 65550 146432 78503
rect 146588 78266 146616 79562
rect 146680 79150 146708 79698
rect 146818 79642 146846 80036
rect 146910 79937 146938 80036
rect 147002 79966 147030 80036
rect 147094 79966 147122 80036
rect 147186 79966 147214 80036
rect 146990 79960 147042 79966
rect 146896 79928 146952 79937
rect 146990 79902 147042 79908
rect 147082 79960 147134 79966
rect 147082 79902 147134 79908
rect 147174 79960 147226 79966
rect 147174 79902 147226 79908
rect 146896 79863 146952 79872
rect 147278 79778 147306 80036
rect 147370 79971 147398 80036
rect 147356 79962 147412 79971
rect 147462 79966 147490 80036
rect 147554 79966 147582 80036
rect 147356 79897 147412 79906
rect 147450 79960 147502 79966
rect 147450 79902 147502 79908
rect 147542 79960 147594 79966
rect 147646 79937 147674 80036
rect 147542 79902 147594 79908
rect 147632 79928 147688 79937
rect 147632 79863 147688 79872
rect 147232 79762 147306 79778
rect 146944 79756 146996 79762
rect 146944 79698 146996 79704
rect 147220 79756 147306 79762
rect 147272 79750 147306 79756
rect 147402 79792 147458 79801
rect 147738 79778 147766 80036
rect 147830 79898 147858 80036
rect 147922 79966 147950 80036
rect 147910 79960 147962 79966
rect 148014 79937 148042 80036
rect 148106 79966 148134 80036
rect 148094 79960 148146 79966
rect 147910 79902 147962 79908
rect 148000 79928 148056 79937
rect 147818 79892 147870 79898
rect 148094 79902 148146 79908
rect 148198 79903 148226 80036
rect 148000 79863 148056 79872
rect 148184 79894 148240 79903
rect 148290 79898 148318 80036
rect 148382 79898 148410 80036
rect 147818 79834 147870 79840
rect 148184 79829 148240 79838
rect 148278 79892 148330 79898
rect 148278 79834 148330 79840
rect 148370 79892 148422 79898
rect 148370 79834 148422 79840
rect 147738 79762 147812 79778
rect 147402 79727 147458 79736
rect 147496 79756 147548 79762
rect 147220 79698 147272 79704
rect 146818 79614 146892 79642
rect 146760 79484 146812 79490
rect 146760 79426 146812 79432
rect 146772 79393 146800 79426
rect 146758 79384 146814 79393
rect 146758 79319 146814 79328
rect 146668 79144 146720 79150
rect 146668 79086 146720 79092
rect 146576 78260 146628 78266
rect 146576 78202 146628 78208
rect 146772 75682 146800 79319
rect 146864 76673 146892 79614
rect 146850 76664 146906 76673
rect 146850 76599 146906 76608
rect 146760 75676 146812 75682
rect 146760 75618 146812 75624
rect 146668 73160 146720 73166
rect 146956 73154 146984 79698
rect 147036 79688 147088 79694
rect 147036 79630 147088 79636
rect 147128 79688 147180 79694
rect 147128 79630 147180 79636
rect 147048 79082 147076 79630
rect 147140 79286 147168 79630
rect 147220 79620 147272 79626
rect 147220 79562 147272 79568
rect 147128 79280 147180 79286
rect 147232 79257 147260 79562
rect 147416 79558 147444 79727
rect 147738 79756 147824 79762
rect 147738 79750 147772 79756
rect 147496 79698 147548 79704
rect 147772 79698 147824 79704
rect 148232 79756 148284 79762
rect 148232 79698 148284 79704
rect 147404 79552 147456 79558
rect 147404 79494 147456 79500
rect 147404 79416 147456 79422
rect 147508 79393 147536 79698
rect 147864 79688 147916 79694
rect 147862 79656 147864 79665
rect 147916 79656 147918 79665
rect 147772 79620 147824 79626
rect 148138 79656 148194 79665
rect 147862 79591 147918 79600
rect 147956 79620 148008 79626
rect 147772 79562 147824 79568
rect 147588 79552 147640 79558
rect 147588 79494 147640 79500
rect 147404 79358 147456 79364
rect 147494 79384 147550 79393
rect 147416 79257 147444 79358
rect 147494 79319 147550 79328
rect 147128 79222 147180 79228
rect 147218 79248 147274 79257
rect 147036 79076 147088 79082
rect 147036 79018 147088 79024
rect 147036 78940 147088 78946
rect 147036 78882 147088 78888
rect 146720 73126 146984 73154
rect 146668 73102 146720 73108
rect 146680 72418 146708 73102
rect 146668 72412 146720 72418
rect 146668 72354 146720 72360
rect 146758 71768 146814 71777
rect 146758 71703 146814 71712
rect 146772 70394 146800 71703
rect 146772 70366 146984 70394
rect 146392 65544 146444 65550
rect 146392 65486 146444 65492
rect 146208 17264 146260 17270
rect 146208 17206 146260 17212
rect 145116 16546 145512 16574
rect 144828 4820 144880 4826
rect 144828 4762 144880 4768
rect 144736 3936 144788 3942
rect 144736 3878 144788 3884
rect 144748 480 144776 3878
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146956 3806 146984 70366
rect 147048 69902 147076 78882
rect 147140 76566 147168 79222
rect 147218 79183 147274 79192
rect 147402 79248 147458 79257
rect 147402 79183 147458 79192
rect 147220 79076 147272 79082
rect 147220 79018 147272 79024
rect 147128 76560 147180 76566
rect 147128 76502 147180 76508
rect 147232 75070 147260 79018
rect 147310 78704 147366 78713
rect 147310 78639 147366 78648
rect 147220 75064 147272 75070
rect 147220 75006 147272 75012
rect 147036 69896 147088 69902
rect 147036 69838 147088 69844
rect 147232 69698 147260 75006
rect 147036 69692 147088 69698
rect 147036 69634 147088 69640
rect 147220 69692 147272 69698
rect 147220 69634 147272 69640
rect 146944 3800 146996 3806
rect 146944 3742 146996 3748
rect 147048 3330 147076 69634
rect 147128 69012 147180 69018
rect 147128 68954 147180 68960
rect 147140 3738 147168 68954
rect 147220 66224 147272 66230
rect 147220 66166 147272 66172
rect 147128 3732 147180 3738
rect 147128 3674 147180 3680
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 147036 3324 147088 3330
rect 147036 3266 147088 3272
rect 147140 480 147168 3538
rect 147232 3058 147260 66166
rect 147324 60042 147352 78639
rect 147404 72412 147456 72418
rect 147404 72354 147456 72360
rect 147416 64190 147444 72354
rect 147404 64184 147456 64190
rect 147404 64126 147456 64132
rect 147312 60036 147364 60042
rect 147312 59978 147364 59984
rect 147508 36922 147536 79319
rect 147496 36916 147548 36922
rect 147496 36858 147548 36864
rect 147600 32706 147628 79494
rect 147680 79212 147732 79218
rect 147680 79154 147732 79160
rect 147692 53174 147720 79154
rect 147784 78810 147812 79562
rect 147772 78804 147824 78810
rect 147772 78746 147824 78752
rect 147784 57254 147812 78746
rect 147876 75614 147904 79591
rect 148138 79591 148194 79600
rect 147956 79562 148008 79568
rect 147968 79286 147996 79562
rect 148046 79384 148102 79393
rect 148046 79319 148102 79328
rect 147956 79280 148008 79286
rect 147956 79222 148008 79228
rect 147864 75608 147916 75614
rect 147864 75550 147916 75556
rect 148060 74118 148088 79319
rect 148152 75478 148180 79591
rect 148244 79218 148272 79698
rect 148324 79688 148376 79694
rect 148474 79676 148502 80036
rect 148324 79630 148376 79636
rect 148428 79648 148502 79676
rect 148232 79212 148284 79218
rect 148232 79154 148284 79160
rect 148336 78334 148364 79630
rect 148324 78328 148376 78334
rect 148324 78270 148376 78276
rect 148336 77654 148364 78270
rect 148324 77648 148376 77654
rect 148324 77590 148376 77596
rect 148324 77512 148376 77518
rect 148324 77454 148376 77460
rect 148140 75472 148192 75478
rect 148140 75414 148192 75420
rect 148048 74112 148100 74118
rect 148048 74054 148100 74060
rect 148060 72146 148088 74054
rect 148048 72140 148100 72146
rect 148048 72082 148100 72088
rect 148152 71774 148180 75414
rect 147876 71746 148180 71774
rect 147876 69834 147904 71746
rect 147864 69828 147916 69834
rect 147864 69770 147916 69776
rect 147772 57248 147824 57254
rect 147772 57190 147824 57196
rect 147680 53168 147732 53174
rect 147680 53110 147732 53116
rect 147588 32700 147640 32706
rect 147588 32642 147640 32648
rect 148336 3534 148364 77454
rect 148428 77042 148456 79648
rect 148566 79608 148594 80036
rect 148658 79937 148686 80036
rect 148644 79928 148700 79937
rect 148644 79863 148700 79872
rect 148750 79778 148778 80036
rect 148842 79966 148870 80036
rect 148934 79966 148962 80036
rect 148830 79960 148882 79966
rect 148830 79902 148882 79908
rect 148922 79960 148974 79966
rect 148922 79902 148974 79908
rect 148876 79824 148928 79830
rect 148874 79792 148876 79801
rect 149026 79812 149054 80036
rect 149118 79966 149146 80036
rect 149210 79966 149238 80036
rect 149106 79960 149158 79966
rect 149106 79902 149158 79908
rect 149198 79960 149250 79966
rect 149198 79902 149250 79908
rect 149152 79824 149204 79830
rect 148928 79792 148930 79801
rect 148750 79750 148824 79778
rect 148692 79688 148744 79694
rect 148692 79630 148744 79636
rect 148520 79580 148594 79608
rect 148520 78033 148548 79580
rect 148600 79484 148652 79490
rect 148600 79426 148652 79432
rect 148506 78024 148562 78033
rect 148506 77959 148562 77968
rect 148612 77897 148640 79426
rect 148704 79393 148732 79630
rect 148690 79384 148746 79393
rect 148690 79319 148746 79328
rect 148690 79248 148746 79257
rect 148690 79183 148746 79192
rect 148704 79014 148732 79183
rect 148692 79008 148744 79014
rect 148692 78950 148744 78956
rect 148796 78674 148824 79750
rect 149026 79784 149100 79812
rect 148874 79727 148930 79736
rect 149072 79694 149100 79784
rect 149152 79766 149204 79772
rect 149060 79688 149112 79694
rect 149060 79630 149112 79636
rect 148966 79248 149022 79257
rect 148966 79183 149022 79192
rect 148796 78646 148916 78674
rect 148598 77888 148654 77897
rect 148598 77823 148654 77832
rect 148508 77648 148560 77654
rect 148508 77590 148560 77596
rect 148416 77036 148468 77042
rect 148416 76978 148468 76984
rect 148428 65686 148456 76978
rect 148520 70394 148548 77590
rect 148612 71774 148640 77823
rect 148888 76974 148916 78646
rect 148876 76968 148928 76974
rect 148876 76910 148928 76916
rect 148784 72140 148836 72146
rect 148784 72082 148836 72088
rect 148612 71746 148732 71774
rect 148520 70366 148640 70394
rect 148416 65680 148468 65686
rect 148416 65622 148468 65628
rect 148416 59356 148468 59362
rect 148416 59298 148468 59304
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148428 3058 148456 59298
rect 148508 52896 148560 52902
rect 148508 52838 148560 52844
rect 148520 3942 148548 52838
rect 148612 36854 148640 70366
rect 148704 44946 148732 71746
rect 148796 49162 148824 72082
rect 148888 71126 148916 76910
rect 148876 71120 148928 71126
rect 148876 71062 148928 71068
rect 148980 58818 149008 79183
rect 149060 78940 149112 78946
rect 149060 78882 149112 78888
rect 148968 58812 149020 58818
rect 148968 58754 149020 58760
rect 148784 49156 148836 49162
rect 148784 49098 148836 49104
rect 148692 44940 148744 44946
rect 148692 44882 148744 44888
rect 148600 36848 148652 36854
rect 148600 36790 148652 36796
rect 149072 18902 149100 78882
rect 149164 78402 149192 79766
rect 149302 79744 149330 80036
rect 149394 79971 149422 80036
rect 149380 79962 149436 79971
rect 149380 79897 149436 79906
rect 149486 79898 149514 80036
rect 149474 79892 149526 79898
rect 149474 79834 149526 79840
rect 149426 79792 149482 79801
rect 149302 79716 149376 79744
rect 149578 79778 149606 80036
rect 149670 79966 149698 80036
rect 149762 79966 149790 80036
rect 149854 79966 149882 80036
rect 149658 79960 149710 79966
rect 149658 79902 149710 79908
rect 149750 79960 149802 79966
rect 149750 79902 149802 79908
rect 149842 79960 149894 79966
rect 149842 79902 149894 79908
rect 149704 79824 149756 79830
rect 149578 79750 149652 79778
rect 149704 79766 149756 79772
rect 149946 79778 149974 80036
rect 150038 79971 150066 80036
rect 150024 79962 150080 79971
rect 150024 79897 150080 79906
rect 150130 79898 150158 80036
rect 150222 79937 150250 80036
rect 150208 79928 150264 79937
rect 150118 79892 150170 79898
rect 150208 79863 150264 79872
rect 150118 79834 150170 79840
rect 150314 79778 150342 80036
rect 150406 79971 150434 80036
rect 150392 79962 150448 79971
rect 150392 79897 150448 79906
rect 150498 79778 150526 80036
rect 150590 79937 150618 80036
rect 150682 79966 150710 80036
rect 150670 79960 150722 79966
rect 150576 79928 150632 79937
rect 150670 79902 150722 79908
rect 150576 79863 150632 79872
rect 150622 79792 150678 79801
rect 149426 79727 149482 79736
rect 149244 79620 149296 79626
rect 149244 79562 149296 79568
rect 149256 78878 149284 79562
rect 149244 78872 149296 78878
rect 149244 78814 149296 78820
rect 149152 78396 149204 78402
rect 149152 78338 149204 78344
rect 149164 76770 149192 78338
rect 149152 76764 149204 76770
rect 149152 76706 149204 76712
rect 149256 47734 149284 78814
rect 149348 76265 149376 79716
rect 149440 79676 149468 79727
rect 149440 79648 149560 79676
rect 149426 79248 149482 79257
rect 149426 79183 149482 79192
rect 149334 76256 149390 76265
rect 149334 76191 149390 76200
rect 149440 71774 149468 79183
rect 149532 78169 149560 79648
rect 149518 78160 149574 78169
rect 149518 78095 149574 78104
rect 149532 76634 149560 78095
rect 149520 76628 149572 76634
rect 149520 76570 149572 76576
rect 149624 76401 149652 79750
rect 149610 76392 149666 76401
rect 149610 76327 149666 76336
rect 149716 76276 149744 79766
rect 149796 79756 149848 79762
rect 149946 79750 150020 79778
rect 150314 79762 150388 79778
rect 150314 79756 150400 79762
rect 150314 79750 150348 79756
rect 149796 79698 149848 79704
rect 149808 79665 149836 79698
rect 149888 79688 149940 79694
rect 149794 79656 149850 79665
rect 149888 79630 149940 79636
rect 149794 79591 149850 79600
rect 149796 76764 149848 76770
rect 149796 76706 149848 76712
rect 149624 76248 149744 76276
rect 149624 75478 149652 76248
rect 149612 75472 149664 75478
rect 149612 75414 149664 75420
rect 149440 71746 149744 71774
rect 149244 47728 149296 47734
rect 149244 47670 149296 47676
rect 149244 47592 149296 47598
rect 149244 47534 149296 47540
rect 149060 18896 149112 18902
rect 149060 18838 149112 18844
rect 149256 16574 149284 47534
rect 149256 16546 149560 16574
rect 148508 3936 148560 3942
rect 148508 3878 148560 3884
rect 147220 3052 147272 3058
rect 147220 2994 147272 3000
rect 148324 3052 148376 3058
rect 148324 2994 148376 3000
rect 148416 3052 148468 3058
rect 148416 2994 148468 3000
rect 148336 480 148364 2994
rect 149532 480 149560 16546
rect 149716 3874 149744 71746
rect 149808 51882 149836 76706
rect 149900 75410 149928 79630
rect 149992 78946 150020 79750
rect 150498 79750 150572 79778
rect 150348 79698 150400 79704
rect 150440 79688 150492 79694
rect 150070 79656 150126 79665
rect 150440 79630 150492 79636
rect 150070 79591 150126 79600
rect 149980 78940 150032 78946
rect 149980 78882 150032 78888
rect 149980 76628 150032 76634
rect 149980 76570 150032 76576
rect 149888 75404 149940 75410
rect 149888 75346 149940 75352
rect 149900 64326 149928 75346
rect 149888 64320 149940 64326
rect 149888 64262 149940 64268
rect 149796 51876 149848 51882
rect 149796 51818 149848 51824
rect 149992 49094 150020 76570
rect 150084 70394 150112 79591
rect 150164 79552 150216 79558
rect 150452 79529 150480 79630
rect 150164 79494 150216 79500
rect 150254 79520 150310 79529
rect 150176 75546 150204 79494
rect 150254 79455 150310 79464
rect 150438 79520 150494 79529
rect 150438 79455 150494 79464
rect 150164 75540 150216 75546
rect 150164 75482 150216 75488
rect 150268 74322 150296 79455
rect 150346 79248 150402 79257
rect 150346 79183 150402 79192
rect 150256 74316 150308 74322
rect 150256 74258 150308 74264
rect 150084 70366 150204 70394
rect 150176 64874 150204 70366
rect 150084 64846 150204 64874
rect 149980 49088 150032 49094
rect 149980 49030 150032 49036
rect 150084 23050 150112 64846
rect 150072 23044 150124 23050
rect 150072 22986 150124 22992
rect 150360 9246 150388 79183
rect 150544 78441 150572 79750
rect 150622 79727 150678 79736
rect 150774 79744 150802 80036
rect 150866 79971 150894 80036
rect 150852 79962 150908 79971
rect 150852 79897 150908 79906
rect 150958 79898 150986 80036
rect 150946 79892 150998 79898
rect 150946 79834 150998 79840
rect 150898 79792 150954 79801
rect 150636 79506 150664 79727
rect 150774 79716 150848 79744
rect 151050 79778 151078 80036
rect 151142 79937 151170 80036
rect 151234 79966 151262 80036
rect 151326 79971 151354 80036
rect 151222 79960 151274 79966
rect 151128 79928 151184 79937
rect 151222 79902 151274 79908
rect 151312 79962 151368 79971
rect 151418 79966 151446 80036
rect 151312 79897 151368 79906
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151128 79863 151184 79872
rect 151176 79824 151228 79830
rect 151050 79750 151124 79778
rect 151176 79766 151228 79772
rect 151266 79792 151322 79801
rect 150898 79727 150954 79736
rect 150636 79478 150756 79506
rect 150624 78736 150676 78742
rect 150624 78678 150676 78684
rect 150530 78432 150586 78441
rect 150530 78367 150586 78376
rect 150544 77353 150572 78367
rect 150530 77344 150586 77353
rect 150530 77279 150586 77288
rect 150636 67046 150664 78678
rect 150728 70394 150756 79478
rect 150820 71534 150848 79716
rect 150912 74254 150940 79727
rect 150992 79620 151044 79626
rect 150992 79562 151044 79568
rect 151004 79150 151032 79562
rect 151096 79393 151124 79750
rect 151082 79384 151138 79393
rect 151082 79319 151138 79328
rect 150992 79144 151044 79150
rect 150992 79086 151044 79092
rect 150990 77344 151046 77353
rect 150990 77279 151046 77288
rect 151004 76786 151032 77279
rect 151096 76906 151124 79319
rect 151188 78742 151216 79766
rect 151510 79744 151538 80036
rect 151266 79727 151322 79736
rect 151176 78736 151228 78742
rect 151176 78678 151228 78684
rect 151280 78674 151308 79727
rect 151464 79716 151538 79744
rect 151360 79688 151412 79694
rect 151360 79630 151412 79636
rect 151372 79529 151400 79630
rect 151358 79520 151414 79529
rect 151358 79455 151414 79464
rect 151268 78668 151320 78674
rect 151268 78610 151320 78616
rect 151084 76900 151136 76906
rect 151084 76842 151136 76848
rect 151004 76758 151216 76786
rect 150900 74248 150952 74254
rect 150900 74190 150952 74196
rect 150808 71528 150860 71534
rect 150808 71470 150860 71476
rect 150820 70922 150848 71470
rect 150808 70916 150860 70922
rect 150808 70858 150860 70864
rect 150728 70378 151124 70394
rect 150728 70372 151136 70378
rect 150728 70366 151084 70372
rect 151084 70314 151136 70320
rect 150624 67040 150676 67046
rect 150624 66982 150676 66988
rect 151096 10538 151124 70314
rect 151188 43586 151216 76758
rect 151268 70916 151320 70922
rect 151268 70858 151320 70864
rect 151280 57390 151308 70858
rect 151372 70394 151400 79455
rect 151464 78577 151492 79716
rect 151602 79676 151630 80036
rect 151694 79801 151722 80036
rect 151786 79937 151814 80036
rect 151772 79928 151828 79937
rect 151878 79898 151906 80036
rect 151772 79863 151828 79872
rect 151866 79892 151918 79898
rect 151866 79834 151918 79840
rect 151680 79792 151736 79801
rect 151970 79744 151998 80036
rect 152062 79966 152090 80036
rect 152050 79960 152102 79966
rect 152050 79902 152102 79908
rect 152154 79812 152182 80036
rect 152246 79830 152274 80036
rect 151680 79727 151736 79736
rect 151556 79648 151630 79676
rect 151924 79716 151998 79744
rect 152108 79784 152182 79812
rect 152234 79824 152286 79830
rect 152232 79792 152234 79801
rect 152286 79792 152288 79801
rect 151726 79656 151782 79665
rect 151450 78568 151506 78577
rect 151450 78503 151506 78512
rect 151556 77314 151584 79648
rect 151726 79591 151782 79600
rect 151820 79620 151872 79626
rect 151636 78668 151688 78674
rect 151636 78610 151688 78616
rect 151544 77308 151596 77314
rect 151544 77250 151596 77256
rect 151452 77240 151504 77246
rect 151452 77182 151504 77188
rect 151464 76838 151492 77182
rect 151452 76832 151504 76838
rect 151452 76774 151504 76780
rect 151372 70366 151492 70394
rect 151268 57384 151320 57390
rect 151268 57326 151320 57332
rect 151176 43580 151228 43586
rect 151176 43522 151228 43528
rect 151464 12034 151492 70366
rect 151648 17542 151676 78610
rect 151740 74186 151768 79591
rect 151820 79562 151872 79568
rect 151728 74180 151780 74186
rect 151728 74122 151780 74128
rect 151832 71738 151860 79562
rect 151924 79218 151952 79716
rect 151912 79212 151964 79218
rect 151912 79154 151964 79160
rect 151910 79112 151966 79121
rect 151910 79047 151966 79056
rect 151820 71732 151872 71738
rect 151820 71674 151872 71680
rect 151832 71466 151860 71674
rect 151820 71460 151872 71466
rect 151820 71402 151872 71408
rect 151924 47666 151952 79047
rect 152004 78668 152056 78674
rect 152004 78610 152056 78616
rect 151912 47660 151964 47666
rect 151912 47602 151964 47608
rect 152016 35426 152044 78610
rect 152108 74390 152136 79784
rect 152232 79727 152288 79736
rect 152338 79744 152366 80036
rect 152430 79966 152458 80036
rect 152418 79960 152470 79966
rect 152418 79902 152470 79908
rect 152522 79812 152550 80036
rect 152614 79971 152642 80036
rect 152600 79962 152656 79971
rect 152600 79897 152656 79906
rect 152706 79898 152734 80036
rect 152798 79903 152826 80036
rect 152890 79966 152918 80036
rect 152982 79966 153010 80036
rect 152878 79960 152930 79966
rect 152694 79892 152746 79898
rect 152694 79834 152746 79840
rect 152784 79894 152840 79903
rect 152878 79902 152930 79908
rect 152970 79960 153022 79966
rect 152970 79902 153022 79908
rect 152784 79829 152840 79838
rect 152970 79824 153022 79830
rect 152476 79784 152550 79812
rect 152890 79784 152970 79812
rect 152338 79716 152412 79744
rect 152188 79688 152240 79694
rect 152188 79630 152240 79636
rect 152096 74384 152148 74390
rect 152096 74326 152148 74332
rect 152108 72146 152136 74326
rect 152200 73982 152228 79630
rect 152280 79212 152332 79218
rect 152280 79154 152332 79160
rect 152188 73976 152240 73982
rect 152188 73918 152240 73924
rect 152188 73840 152240 73846
rect 152188 73782 152240 73788
rect 152096 72140 152148 72146
rect 152096 72082 152148 72088
rect 152004 35420 152056 35426
rect 152004 35362 152056 35368
rect 151636 17536 151688 17542
rect 151636 17478 151688 17484
rect 152200 16574 152228 73782
rect 152292 70242 152320 79154
rect 152384 75993 152412 79716
rect 152476 79665 152504 79784
rect 152890 79778 152918 79784
rect 152844 79750 152918 79778
rect 152970 79766 153022 79772
rect 153074 79778 153102 80036
rect 153166 79898 153194 80036
rect 153154 79892 153206 79898
rect 153154 79834 153206 79840
rect 153074 79750 153148 79778
rect 152648 79688 152700 79694
rect 152462 79656 152518 79665
rect 152648 79630 152700 79636
rect 152462 79591 152518 79600
rect 152556 79620 152608 79626
rect 152370 75984 152426 75993
rect 152370 75919 152426 75928
rect 152476 70394 152504 79591
rect 152556 79562 152608 79568
rect 152568 71330 152596 79562
rect 152660 79354 152688 79630
rect 152648 79348 152700 79354
rect 152648 79290 152700 79296
rect 152660 76770 152688 79290
rect 152648 76764 152700 76770
rect 152648 76706 152700 76712
rect 152844 74633 152872 79750
rect 153016 79688 153068 79694
rect 152922 79656 152978 79665
rect 153016 79630 153068 79636
rect 152922 79591 152978 79600
rect 152830 74624 152886 74633
rect 152830 74559 152886 74568
rect 152936 73846 152964 79591
rect 153028 79121 153056 79630
rect 153120 79529 153148 79750
rect 153258 79744 153286 80036
rect 153212 79716 153286 79744
rect 153350 79744 153378 80036
rect 153442 79966 153470 80036
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 153534 79744 153562 80036
rect 153626 79937 153654 80036
rect 153612 79928 153668 79937
rect 153718 79898 153746 80036
rect 153612 79863 153668 79872
rect 153706 79892 153758 79898
rect 153706 79834 153758 79840
rect 153810 79744 153838 80036
rect 153902 79830 153930 80036
rect 153890 79824 153942 79830
rect 153890 79766 153942 79772
rect 153350 79716 153424 79744
rect 153534 79716 153608 79744
rect 153106 79520 153162 79529
rect 153106 79455 153162 79464
rect 153014 79112 153070 79121
rect 153014 79047 153070 79056
rect 153120 78674 153148 79455
rect 153108 78668 153160 78674
rect 153108 78610 153160 78616
rect 153212 76702 153240 79716
rect 153292 79620 153344 79626
rect 153292 79562 153344 79568
rect 153304 76809 153332 79562
rect 153290 76800 153346 76809
rect 153290 76735 153346 76744
rect 153200 76696 153252 76702
rect 153200 76638 153252 76644
rect 153396 74497 153424 79716
rect 153476 79552 153528 79558
rect 153474 79520 153476 79529
rect 153528 79520 153530 79529
rect 153474 79455 153530 79464
rect 153488 77790 153516 79455
rect 153476 77784 153528 77790
rect 153476 77726 153528 77732
rect 153476 76696 153528 76702
rect 153476 76638 153528 76644
rect 153382 74488 153438 74497
rect 153382 74423 153438 74432
rect 152924 73840 152976 73846
rect 152924 73782 152976 73788
rect 153488 73137 153516 76638
rect 153474 73128 153530 73137
rect 153474 73063 153530 73072
rect 153292 72616 153344 72622
rect 153292 72558 153344 72564
rect 152832 72140 152884 72146
rect 152832 72082 152884 72088
rect 152740 71460 152792 71466
rect 152740 71402 152792 71408
rect 152556 71324 152608 71330
rect 152556 71266 152608 71272
rect 152384 70366 152504 70394
rect 152568 70394 152596 71266
rect 152568 70366 152688 70394
rect 152280 70236 152332 70242
rect 152280 70178 152332 70184
rect 152200 16546 152320 16574
rect 151452 12028 151504 12034
rect 151452 11970 151504 11976
rect 151084 10532 151136 10538
rect 151084 10474 151136 10480
rect 150348 9240 150400 9246
rect 150348 9182 150400 9188
rect 151820 3936 151872 3942
rect 151820 3878 151872 3884
rect 149704 3868 149756 3874
rect 149704 3810 149756 3816
rect 150624 3324 150676 3330
rect 150624 3266 150676 3272
rect 150636 480 150664 3266
rect 151832 480 151860 3878
rect 152292 3482 152320 16546
rect 152384 5098 152412 70366
rect 152556 70236 152608 70242
rect 152556 70178 152608 70184
rect 152462 63064 152518 63073
rect 152462 62999 152518 63008
rect 152372 5092 152424 5098
rect 152372 5034 152424 5040
rect 152476 3602 152504 62999
rect 152568 16114 152596 70178
rect 152660 28558 152688 70366
rect 152752 39642 152780 71402
rect 152844 54670 152872 72082
rect 153304 69766 153332 72558
rect 153580 71398 153608 79716
rect 153672 79716 153838 79744
rect 153994 79744 154022 80036
rect 154086 79812 154114 80036
rect 154178 79966 154206 80036
rect 154270 79966 154298 80036
rect 154362 79966 154390 80036
rect 154454 79966 154482 80036
rect 154166 79960 154218 79966
rect 154166 79902 154218 79908
rect 154258 79960 154310 79966
rect 154258 79902 154310 79908
rect 154350 79960 154402 79966
rect 154350 79902 154402 79908
rect 154442 79960 154494 79966
rect 154442 79902 154494 79908
rect 154212 79824 154264 79830
rect 154086 79784 154160 79812
rect 153994 79716 154068 79744
rect 153672 72622 153700 79716
rect 153842 79656 153898 79665
rect 153752 79620 153804 79626
rect 153842 79591 153898 79600
rect 153936 79620 153988 79626
rect 153752 79562 153804 79568
rect 153764 73030 153792 79562
rect 153856 74474 153884 79591
rect 153936 79562 153988 79568
rect 153948 79529 153976 79562
rect 153934 79520 153990 79529
rect 153934 79455 153990 79464
rect 153948 78674 153976 79455
rect 153936 78668 153988 78674
rect 153936 78610 153988 78616
rect 154040 76673 154068 79716
rect 154026 76664 154082 76673
rect 154026 76599 154082 76608
rect 153856 74446 154068 74474
rect 153752 73024 153804 73030
rect 153752 72966 153804 72972
rect 153660 72616 153712 72622
rect 153660 72558 153712 72564
rect 153568 71392 153620 71398
rect 153568 71334 153620 71340
rect 153580 71194 153608 71334
rect 153568 71188 153620 71194
rect 153568 71130 153620 71136
rect 153568 71052 153620 71058
rect 153568 70994 153620 71000
rect 153580 70009 153608 70994
rect 153566 70000 153622 70009
rect 153566 69935 153622 69944
rect 153292 69760 153344 69766
rect 153292 69702 153344 69708
rect 153764 65618 153792 72966
rect 154040 72894 154068 74446
rect 154028 72888 154080 72894
rect 154028 72830 154080 72836
rect 153936 71188 153988 71194
rect 153936 71130 153988 71136
rect 153844 69760 153896 69766
rect 153844 69702 153896 69708
rect 153752 65612 153804 65618
rect 153752 65554 153804 65560
rect 152832 54664 152884 54670
rect 152832 54606 152884 54612
rect 152740 39636 152792 39642
rect 152740 39578 152792 39584
rect 152648 28552 152700 28558
rect 152648 28494 152700 28500
rect 152556 16108 152608 16114
rect 152556 16050 152608 16056
rect 153856 6390 153884 69702
rect 153948 14754 153976 71130
rect 154040 24410 154068 72830
rect 154132 71058 154160 79784
rect 154396 79824 154448 79830
rect 154212 79766 154264 79772
rect 154302 79792 154358 79801
rect 154224 78713 154252 79766
rect 154396 79766 154448 79772
rect 154302 79727 154358 79736
rect 154316 79694 154344 79727
rect 154304 79688 154356 79694
rect 154304 79630 154356 79636
rect 154210 78704 154266 78713
rect 154210 78639 154266 78648
rect 154316 78588 154344 79630
rect 154224 78560 154344 78588
rect 154224 74118 154252 78560
rect 154302 78160 154358 78169
rect 154302 78095 154358 78104
rect 154212 74112 154264 74118
rect 154212 74054 154264 74060
rect 154210 73128 154266 73137
rect 154210 73063 154266 73072
rect 154120 71052 154172 71058
rect 154120 70994 154172 71000
rect 154118 70000 154174 70009
rect 154118 69935 154174 69944
rect 154132 32638 154160 69935
rect 154224 38214 154252 73063
rect 154316 44878 154344 78095
rect 154408 77897 154436 79766
rect 154546 79744 154574 80036
rect 154638 79898 154666 80036
rect 154730 79971 154758 80036
rect 154716 79962 154772 79971
rect 154822 79966 154850 80036
rect 154626 79892 154678 79898
rect 154716 79897 154772 79906
rect 154810 79960 154862 79966
rect 154810 79902 154862 79908
rect 154626 79834 154678 79840
rect 154914 79835 154942 80036
rect 155006 79966 155034 80036
rect 155098 79971 155126 80036
rect 154994 79960 155046 79966
rect 154994 79902 155046 79908
rect 155084 79962 155140 79971
rect 155190 79966 155218 80036
rect 155084 79897 155140 79906
rect 155178 79960 155230 79966
rect 155178 79902 155230 79908
rect 154900 79826 154956 79835
rect 155282 79801 155310 80036
rect 155374 79898 155402 80036
rect 155362 79892 155414 79898
rect 155362 79834 155414 79840
rect 155466 79830 155494 80036
rect 155454 79824 155506 79830
rect 154500 79716 154574 79744
rect 154764 79756 154816 79762
rect 154900 79761 154956 79770
rect 155130 79792 155186 79801
rect 154500 79665 154528 79716
rect 155130 79727 155186 79736
rect 155268 79792 155324 79801
rect 155558 79812 155586 80036
rect 155650 79937 155678 80036
rect 155636 79928 155692 79937
rect 155636 79863 155692 79872
rect 155558 79784 155632 79812
rect 155454 79766 155506 79772
rect 155268 79727 155324 79736
rect 154764 79698 154816 79704
rect 154672 79688 154724 79694
rect 154486 79656 154542 79665
rect 154672 79630 154724 79636
rect 154486 79591 154542 79600
rect 154578 79520 154634 79529
rect 154578 79455 154634 79464
rect 154488 78668 154540 78674
rect 154488 78610 154540 78616
rect 154394 77888 154450 77897
rect 154394 77823 154450 77832
rect 154396 77784 154448 77790
rect 154396 77726 154448 77732
rect 154304 44872 154356 44878
rect 154304 44814 154356 44820
rect 154408 41002 154436 77726
rect 154396 40996 154448 41002
rect 154396 40938 154448 40944
rect 154212 38208 154264 38214
rect 154212 38150 154264 38156
rect 154120 32632 154172 32638
rect 154120 32574 154172 32580
rect 154028 24404 154080 24410
rect 154028 24346 154080 24352
rect 154500 20262 154528 78610
rect 154592 71670 154620 79455
rect 154580 71664 154632 71670
rect 154580 71606 154632 71612
rect 154684 70310 154712 79630
rect 154776 79257 154804 79698
rect 155144 79676 155172 79727
rect 155500 79688 155552 79694
rect 154854 79656 154910 79665
rect 155144 79648 155264 79676
rect 154854 79591 154910 79600
rect 154948 79620 155000 79626
rect 154762 79248 154818 79257
rect 154762 79183 154818 79192
rect 154868 72962 154896 79591
rect 154948 79562 155000 79568
rect 154856 72956 154908 72962
rect 154856 72898 154908 72904
rect 154672 70304 154724 70310
rect 154672 70246 154724 70252
rect 154960 70106 154988 79562
rect 155132 79552 155184 79558
rect 155132 79494 155184 79500
rect 154948 70100 155000 70106
rect 154948 70042 155000 70048
rect 155144 67590 155172 79494
rect 155236 76702 155264 79648
rect 155604 79665 155632 79784
rect 155742 79744 155770 80036
rect 155834 79937 155862 80036
rect 155820 79928 155876 79937
rect 155926 79898 155954 80036
rect 155820 79863 155876 79872
rect 155914 79892 155966 79898
rect 155914 79834 155966 79840
rect 155696 79716 155770 79744
rect 156018 79744 156046 80036
rect 156110 79971 156138 80036
rect 156096 79962 156152 79971
rect 156096 79897 156152 79906
rect 156202 79898 156230 80036
rect 156294 79966 156322 80036
rect 156386 79966 156414 80036
rect 156478 79971 156506 80036
rect 156282 79960 156334 79966
rect 156282 79902 156334 79908
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156464 79962 156520 79971
rect 156570 79966 156598 80036
rect 156190 79892 156242 79898
rect 156464 79897 156520 79906
rect 156558 79960 156610 79966
rect 156558 79902 156610 79908
rect 156190 79834 156242 79840
rect 156662 79778 156690 80036
rect 156754 79966 156782 80036
rect 156742 79960 156794 79966
rect 156742 79902 156794 79908
rect 156846 79898 156874 80036
rect 156938 79966 156966 80036
rect 156926 79960 156978 79966
rect 156926 79902 156978 79908
rect 156834 79892 156886 79898
rect 156834 79834 156886 79840
rect 157030 79801 157058 80036
rect 156432 79750 156690 79778
rect 157016 79792 157072 79801
rect 156788 79756 156840 79762
rect 156018 79716 156092 79744
rect 155500 79630 155552 79636
rect 155590 79656 155646 79665
rect 155512 77042 155540 79630
rect 155590 79591 155646 79600
rect 155590 79384 155646 79393
rect 155590 79319 155646 79328
rect 155500 77036 155552 77042
rect 155500 76978 155552 76984
rect 155224 76696 155276 76702
rect 155224 76638 155276 76644
rect 155224 71664 155276 71670
rect 155224 71606 155276 71612
rect 155132 67584 155184 67590
rect 155132 67526 155184 67532
rect 154488 20256 154540 20262
rect 154488 20198 154540 20204
rect 155236 20126 155264 71606
rect 155408 70304 155460 70310
rect 155408 70246 155460 70252
rect 155316 70100 155368 70106
rect 155316 70042 155368 70048
rect 155328 42294 155356 70042
rect 155420 46374 155448 70246
rect 155604 50386 155632 79319
rect 155696 74225 155724 79716
rect 155866 79656 155922 79665
rect 155866 79591 155922 79600
rect 155774 79248 155830 79257
rect 155774 79183 155830 79192
rect 155682 74216 155738 74225
rect 155682 74151 155738 74160
rect 155592 50380 155644 50386
rect 155592 50322 155644 50328
rect 155408 46368 155460 46374
rect 155408 46310 155460 46316
rect 155316 42288 155368 42294
rect 155316 42230 155368 42236
rect 155696 34066 155724 74151
rect 155684 34060 155736 34066
rect 155684 34002 155736 34008
rect 155788 20194 155816 79183
rect 155776 20188 155828 20194
rect 155776 20130 155828 20136
rect 155224 20120 155276 20126
rect 155224 20062 155276 20068
rect 154580 19984 154632 19990
rect 154580 19926 154632 19932
rect 154592 16574 154620 19926
rect 155880 18834 155908 79591
rect 155960 76968 156012 76974
rect 155960 76910 156012 76916
rect 155868 18828 155920 18834
rect 155868 18770 155920 18776
rect 154592 16546 155448 16574
rect 153936 14748 153988 14754
rect 153936 14690 153988 14696
rect 153844 6384 153896 6390
rect 153844 6326 153896 6332
rect 152464 3596 152516 3602
rect 152464 3538 152516 3544
rect 152292 3454 153056 3482
rect 153028 480 153056 3454
rect 154212 3052 154264 3058
rect 154212 2994 154264 3000
rect 154224 480 154252 2994
rect 155420 480 155448 16546
rect 155972 14686 156000 76910
rect 156064 75342 156092 79716
rect 156144 79552 156196 79558
rect 156144 79494 156196 79500
rect 156156 78985 156184 79494
rect 156236 79484 156288 79490
rect 156236 79426 156288 79432
rect 156142 78976 156198 78985
rect 156142 78911 156198 78920
rect 156248 78674 156276 79426
rect 156432 79121 156460 79750
rect 157016 79727 157072 79736
rect 157122 79744 157150 80036
rect 157214 79937 157242 80036
rect 157306 79966 157334 80036
rect 157294 79960 157346 79966
rect 157200 79928 157256 79937
rect 157294 79902 157346 79908
rect 157200 79863 157256 79872
rect 157122 79716 157196 79744
rect 156788 79698 156840 79704
rect 156604 79688 156656 79694
rect 156602 79656 156604 79665
rect 156656 79656 156658 79665
rect 156602 79591 156658 79600
rect 156696 79620 156748 79626
rect 156696 79562 156748 79568
rect 156510 79520 156566 79529
rect 156510 79455 156566 79464
rect 156418 79112 156474 79121
rect 156418 79047 156474 79056
rect 156248 78646 156460 78674
rect 156432 75818 156460 78646
rect 156420 75812 156472 75818
rect 156420 75754 156472 75760
rect 156052 75336 156104 75342
rect 156052 75278 156104 75284
rect 156524 73030 156552 79455
rect 156512 73024 156564 73030
rect 156512 72966 156564 72972
rect 156328 72480 156380 72486
rect 156328 72422 156380 72428
rect 156340 64874 156368 72422
rect 156708 71774 156736 79562
rect 156800 75857 156828 79698
rect 156880 79688 156932 79694
rect 156880 79630 156932 79636
rect 156892 78849 156920 79630
rect 157064 79484 157116 79490
rect 157064 79426 157116 79432
rect 156972 79348 157024 79354
rect 156972 79290 157024 79296
rect 156984 79257 157012 79290
rect 156970 79248 157026 79257
rect 156970 79183 157026 79192
rect 156970 79112 157026 79121
rect 156970 79047 157026 79056
rect 156878 78840 156934 78849
rect 156878 78775 156934 78784
rect 156892 76974 156920 78775
rect 156880 76968 156932 76974
rect 156880 76910 156932 76916
rect 156786 75848 156842 75857
rect 156786 75783 156842 75792
rect 156880 75812 156932 75818
rect 156880 75754 156932 75760
rect 156892 75585 156920 75754
rect 156878 75576 156934 75585
rect 156878 75511 156934 75520
rect 156788 75336 156840 75342
rect 156788 75278 156840 75284
rect 156800 74089 156828 75278
rect 156786 74080 156842 74089
rect 156786 74015 156842 74024
rect 156616 71746 156736 71774
rect 156616 70145 156644 71746
rect 156602 70136 156658 70145
rect 156602 70071 156658 70080
rect 156616 67634 156644 70071
rect 156616 67606 156736 67634
rect 156340 64846 156644 64874
rect 156616 16574 156644 64846
rect 156708 25838 156736 67606
rect 156800 36786 156828 74015
rect 156892 64874 156920 75511
rect 156984 72758 157012 79047
rect 157076 73098 157104 79426
rect 157168 75041 157196 79716
rect 157398 79642 157426 80036
rect 157490 79966 157518 80036
rect 157582 79966 157610 80036
rect 157674 79966 157702 80036
rect 157766 79966 157794 80036
rect 157478 79960 157530 79966
rect 157478 79902 157530 79908
rect 157570 79960 157622 79966
rect 157570 79902 157622 79908
rect 157662 79960 157714 79966
rect 157662 79902 157714 79908
rect 157754 79960 157806 79966
rect 157858 79937 157886 80036
rect 157754 79902 157806 79908
rect 157844 79928 157900 79937
rect 157844 79863 157900 79872
rect 157950 79830 157978 80036
rect 158042 79898 158070 80036
rect 158030 79892 158082 79898
rect 158030 79834 158082 79840
rect 157938 79824 157990 79830
rect 157938 79766 157990 79772
rect 158134 79744 158162 80036
rect 158226 79966 158254 80036
rect 158214 79960 158266 79966
rect 158214 79902 158266 79908
rect 158318 79801 158346 80036
rect 158410 79898 158438 80036
rect 158502 79966 158530 80036
rect 158490 79960 158542 79966
rect 158594 79937 158622 80036
rect 158490 79902 158542 79908
rect 158580 79928 158636 79937
rect 158398 79892 158450 79898
rect 158580 79863 158636 79872
rect 158398 79834 158450 79840
rect 158088 79716 158162 79744
rect 158304 79792 158360 79801
rect 158686 79778 158714 80036
rect 158778 79966 158806 80036
rect 158870 79966 158898 80036
rect 158766 79960 158818 79966
rect 158766 79902 158818 79908
rect 158858 79960 158910 79966
rect 158858 79902 158910 79908
rect 158812 79824 158864 79830
rect 158686 79750 158760 79778
rect 158812 79766 158864 79772
rect 158962 79778 158990 80036
rect 159054 79966 159082 80036
rect 159042 79960 159094 79966
rect 159042 79902 159094 79908
rect 159146 79898 159174 80036
rect 159134 79892 159186 79898
rect 159134 79834 159186 79840
rect 158304 79727 158360 79736
rect 157524 79688 157576 79694
rect 157248 79620 157300 79626
rect 157248 79562 157300 79568
rect 157352 79614 157426 79642
rect 157522 79656 157524 79665
rect 157576 79656 157578 79665
rect 157154 75032 157210 75041
rect 157154 74967 157210 74976
rect 157064 73092 157116 73098
rect 157064 73034 157116 73040
rect 156972 72752 157024 72758
rect 156972 72694 157024 72700
rect 156892 64846 157012 64874
rect 156984 42226 157012 64846
rect 156972 42220 157024 42226
rect 156972 42162 157024 42168
rect 156788 36780 156840 36786
rect 156788 36722 156840 36728
rect 157168 31346 157196 74967
rect 157156 31340 157208 31346
rect 157156 31282 157208 31288
rect 156696 25832 156748 25838
rect 156696 25774 156748 25780
rect 156616 16546 156736 16574
rect 155960 14680 156012 14686
rect 155960 14622 156012 14628
rect 156708 3806 156736 16546
rect 157260 7818 157288 79562
rect 157352 73914 157380 79614
rect 157522 79591 157578 79600
rect 157524 79552 157576 79558
rect 157430 79520 157486 79529
rect 157892 79552 157944 79558
rect 157524 79494 157576 79500
rect 157614 79520 157670 79529
rect 157430 79455 157486 79464
rect 157340 73908 157392 73914
rect 157340 73850 157392 73856
rect 157444 72690 157472 79455
rect 157536 75138 157564 79494
rect 157892 79494 157944 79500
rect 157982 79520 158038 79529
rect 157614 79455 157670 79464
rect 157800 79484 157852 79490
rect 157628 77722 157656 79455
rect 157800 79426 157852 79432
rect 157708 79348 157760 79354
rect 157708 79290 157760 79296
rect 157720 78849 157748 79290
rect 157706 78840 157762 78849
rect 157706 78775 157762 78784
rect 157616 77716 157668 77722
rect 157616 77658 157668 77664
rect 157524 75132 157576 75138
rect 157524 75074 157576 75080
rect 157536 74050 157564 75074
rect 157524 74044 157576 74050
rect 157524 73986 157576 73992
rect 157432 72684 157484 72690
rect 157432 72626 157484 72632
rect 157720 72622 157748 78775
rect 157708 72616 157760 72622
rect 157708 72558 157760 72564
rect 157812 72554 157840 79426
rect 157904 79121 157932 79494
rect 158088 79506 158116 79716
rect 158260 79688 158312 79694
rect 158166 79656 158222 79665
rect 158260 79630 158312 79636
rect 158352 79688 158404 79694
rect 158536 79688 158588 79694
rect 158352 79630 158404 79636
rect 158442 79656 158498 79665
rect 158166 79591 158222 79600
rect 158038 79478 158116 79506
rect 158180 79490 158208 79591
rect 158168 79484 158220 79490
rect 157982 79455 158038 79464
rect 158168 79426 158220 79432
rect 157984 79416 158036 79422
rect 157984 79358 158036 79364
rect 158076 79416 158128 79422
rect 158076 79358 158128 79364
rect 158166 79384 158222 79393
rect 157890 79112 157946 79121
rect 157890 79047 157946 79056
rect 157800 72548 157852 72554
rect 157800 72490 157852 72496
rect 157904 70394 157932 79047
rect 157996 72865 158024 79358
rect 158088 78985 158116 79358
rect 158166 79319 158222 79328
rect 158074 78976 158130 78985
rect 158074 78911 158130 78920
rect 158074 74352 158130 74361
rect 158074 74287 158130 74296
rect 157982 72856 158038 72865
rect 157982 72791 158038 72800
rect 157352 70366 157932 70394
rect 157352 24342 157380 70366
rect 157340 24336 157392 24342
rect 157340 24278 157392 24284
rect 157338 21312 157394 21321
rect 157338 21247 157394 21256
rect 157352 16574 157380 21247
rect 157352 16546 157840 16574
rect 157248 7812 157300 7818
rect 157248 7754 157300 7760
rect 156604 3800 156656 3806
rect 156604 3742 156656 3748
rect 156696 3800 156748 3806
rect 156696 3742 156748 3748
rect 156616 480 156644 3742
rect 157812 480 157840 16546
rect 157996 13258 158024 72791
rect 158088 54602 158116 74287
rect 158076 54596 158128 54602
rect 158076 54538 158128 54544
rect 158180 21622 158208 79319
rect 158272 74236 158300 79630
rect 158364 74361 158392 79630
rect 158628 79688 158680 79694
rect 158536 79630 158588 79636
rect 158626 79656 158628 79665
rect 158680 79656 158682 79665
rect 158442 79591 158444 79600
rect 158496 79591 158498 79600
rect 158444 79562 158496 79568
rect 158444 79348 158496 79354
rect 158444 79290 158496 79296
rect 158456 79082 158484 79290
rect 158444 79076 158496 79082
rect 158444 79018 158496 79024
rect 158548 78577 158576 79630
rect 158626 79591 158682 79600
rect 158732 79529 158760 79750
rect 158718 79520 158774 79529
rect 158718 79455 158774 79464
rect 158534 78568 158590 78577
rect 158534 78503 158590 78512
rect 158534 78160 158590 78169
rect 158534 78095 158590 78104
rect 158350 74352 158406 74361
rect 158350 74287 158406 74296
rect 158272 74208 158484 74236
rect 158260 74044 158312 74050
rect 158260 73986 158312 73992
rect 158272 40934 158300 73986
rect 158350 73944 158406 73953
rect 158350 73879 158352 73888
rect 158404 73879 158406 73888
rect 158352 73850 158404 73856
rect 158260 40928 158312 40934
rect 158260 40870 158312 40876
rect 158364 35358 158392 73850
rect 158456 72457 158484 74208
rect 158442 72448 158498 72457
rect 158442 72383 158498 72392
rect 158352 35352 158404 35358
rect 158352 35294 158404 35300
rect 158456 29850 158484 72383
rect 158444 29844 158496 29850
rect 158444 29786 158496 29792
rect 158548 21690 158576 78095
rect 158824 74934 158852 79766
rect 158962 79750 159036 79778
rect 158904 79688 158956 79694
rect 158904 79630 158956 79636
rect 158916 78985 158944 79630
rect 158902 78976 158958 78985
rect 158902 78911 158958 78920
rect 158812 74928 158864 74934
rect 158812 74870 158864 74876
rect 158916 74746 158944 78911
rect 159008 78656 159036 79750
rect 159088 79756 159140 79762
rect 159238 79744 159266 80036
rect 159088 79698 159140 79704
rect 159192 79716 159266 79744
rect 159100 79082 159128 79698
rect 159088 79076 159140 79082
rect 159088 79018 159140 79024
rect 159008 78628 159128 78656
rect 158824 74718 158944 74746
rect 158536 21684 158588 21690
rect 158536 21626 158588 21632
rect 158168 21616 158220 21622
rect 158168 21558 158220 21564
rect 158824 21554 158852 74718
rect 158904 74656 158956 74662
rect 158904 74598 158956 74604
rect 158916 56506 158944 74598
rect 158996 73296 159048 73302
rect 158996 73238 159048 73244
rect 159008 57866 159036 73238
rect 159100 63510 159128 78628
rect 159192 73302 159220 79716
rect 159330 79676 159358 80036
rect 159422 79801 159450 80036
rect 159514 79830 159542 80036
rect 159606 79966 159634 80036
rect 159698 79966 159726 80036
rect 159594 79960 159646 79966
rect 159594 79902 159646 79908
rect 159686 79960 159738 79966
rect 159790 79937 159818 80036
rect 159686 79902 159738 79908
rect 159776 79928 159832 79937
rect 159776 79863 159832 79872
rect 159502 79824 159554 79830
rect 159408 79792 159464 79801
rect 159502 79766 159554 79772
rect 159882 79744 159910 80036
rect 159974 79801 160002 80036
rect 160066 79966 160094 80036
rect 160054 79960 160106 79966
rect 160054 79902 160106 79908
rect 160158 79898 160186 80036
rect 160250 79966 160278 80036
rect 160238 79960 160290 79966
rect 160238 79902 160290 79908
rect 160342 79898 160370 80036
rect 160434 79966 160462 80036
rect 160422 79960 160474 79966
rect 160526 79937 160554 80036
rect 160618 79966 160646 80036
rect 160606 79960 160658 79966
rect 160422 79902 160474 79908
rect 160512 79928 160568 79937
rect 160146 79892 160198 79898
rect 160146 79834 160198 79840
rect 160330 79892 160382 79898
rect 160606 79902 160658 79908
rect 160512 79863 160568 79872
rect 160330 79834 160382 79840
rect 159408 79727 159464 79736
rect 159284 79648 159358 79676
rect 159180 73296 159232 73302
rect 159180 73238 159232 73244
rect 159284 67634 159312 79648
rect 159422 79608 159450 79727
rect 159836 79716 159910 79744
rect 159960 79792 160016 79801
rect 159960 79727 160016 79736
rect 160190 79792 160246 79801
rect 160466 79792 160522 79801
rect 160190 79727 160246 79736
rect 160284 79756 160336 79762
rect 159640 79688 159692 79694
rect 159836 79642 159864 79716
rect 159640 79630 159692 79636
rect 159376 79580 159450 79608
rect 159548 79620 159600 79626
rect 159376 74050 159404 79580
rect 159548 79562 159600 79568
rect 159560 79370 159588 79562
rect 159468 79342 159588 79370
rect 159468 74662 159496 79342
rect 159548 79280 159600 79286
rect 159548 79222 159600 79228
rect 159560 79150 159588 79222
rect 159548 79144 159600 79150
rect 159548 79086 159600 79092
rect 159652 78878 159680 79630
rect 159744 79614 159864 79642
rect 160008 79688 160060 79694
rect 160008 79630 160060 79636
rect 159640 78872 159692 78878
rect 159640 78814 159692 78820
rect 159548 78464 159600 78470
rect 159546 78432 159548 78441
rect 159600 78432 159602 78441
rect 159546 78367 159602 78376
rect 159456 74656 159508 74662
rect 159456 74598 159508 74604
rect 159364 74044 159416 74050
rect 159364 73986 159416 73992
rect 159192 67606 159312 67634
rect 159192 66230 159220 67606
rect 159180 66224 159232 66230
rect 159180 66166 159232 66172
rect 159088 63504 159140 63510
rect 159088 63446 159140 63452
rect 158996 57860 159048 57866
rect 158996 57802 159048 57808
rect 158904 56500 158956 56506
rect 158904 56442 158956 56448
rect 158812 21548 158864 21554
rect 158812 21490 158864 21496
rect 157984 13252 158036 13258
rect 157984 13194 158036 13200
rect 159652 10470 159680 78814
rect 159744 77110 159772 79614
rect 159824 79552 159876 79558
rect 159822 79520 159824 79529
rect 159876 79520 159878 79529
rect 159878 79478 159956 79506
rect 159822 79455 159878 79464
rect 159824 79076 159876 79082
rect 159824 79018 159876 79024
rect 159732 77104 159784 77110
rect 159732 77046 159784 77052
rect 159836 75070 159864 79018
rect 159824 75064 159876 75070
rect 159824 75006 159876 75012
rect 159824 74928 159876 74934
rect 159824 74870 159876 74876
rect 159836 73001 159864 74870
rect 159822 72992 159878 73001
rect 159822 72927 159878 72936
rect 159836 28490 159864 72927
rect 159928 31278 159956 79478
rect 160020 75993 160048 79630
rect 160100 79620 160152 79626
rect 160100 79562 160152 79568
rect 160006 75984 160062 75993
rect 160006 75919 160062 75928
rect 160008 75064 160060 75070
rect 160008 75006 160060 75012
rect 160020 72350 160048 75006
rect 160112 72894 160140 79562
rect 160100 72888 160152 72894
rect 160100 72830 160152 72836
rect 160008 72344 160060 72350
rect 160008 72286 160060 72292
rect 159916 31272 159968 31278
rect 159916 31214 159968 31220
rect 159824 28484 159876 28490
rect 159824 28426 159876 28432
rect 160020 11966 160048 72286
rect 160204 69766 160232 79727
rect 160466 79727 160522 79736
rect 160710 79744 160738 80036
rect 160802 79971 160830 80036
rect 160788 79962 160844 79971
rect 160894 79966 160922 80036
rect 160986 79966 161014 80036
rect 160788 79897 160844 79906
rect 160882 79960 160934 79966
rect 160882 79902 160934 79908
rect 160974 79960 161026 79966
rect 160974 79902 161026 79908
rect 161078 79801 161106 80036
rect 161170 79966 161198 80036
rect 161262 79971 161290 80036
rect 161158 79960 161210 79966
rect 161158 79902 161210 79908
rect 161248 79962 161304 79971
rect 161248 79897 161304 79906
rect 161354 79898 161382 80036
rect 161342 79892 161394 79898
rect 161342 79834 161394 79840
rect 161204 79824 161256 79830
rect 161064 79792 161120 79801
rect 160284 79698 160336 79704
rect 160192 69760 160244 69766
rect 160192 69702 160244 69708
rect 160296 67634 160324 79698
rect 160376 79620 160428 79626
rect 160376 79562 160428 79568
rect 160388 75721 160416 79562
rect 160480 78305 160508 79727
rect 160710 79716 160968 79744
rect 161446 79801 161474 80036
rect 161204 79766 161256 79772
rect 161432 79792 161488 79801
rect 161064 79727 161120 79736
rect 160560 79688 160612 79694
rect 160560 79630 160612 79636
rect 160650 79656 160706 79665
rect 160466 78296 160522 78305
rect 160466 78231 160522 78240
rect 160374 75712 160430 75721
rect 160374 75647 160430 75656
rect 160480 75342 160508 78231
rect 160468 75336 160520 75342
rect 160468 75278 160520 75284
rect 160572 74390 160600 79630
rect 160650 79591 160706 79600
rect 160744 79620 160796 79626
rect 160664 77382 160692 79591
rect 160744 79562 160796 79568
rect 160756 79529 160784 79562
rect 160836 79552 160888 79558
rect 160742 79520 160798 79529
rect 160836 79494 160888 79500
rect 160742 79455 160798 79464
rect 160652 77376 160704 77382
rect 160652 77318 160704 77324
rect 160560 74384 160612 74390
rect 160560 74326 160612 74332
rect 160756 73930 160784 79455
rect 160848 75993 160876 79494
rect 160834 75984 160890 75993
rect 160834 75919 160890 75928
rect 160204 67606 160324 67634
rect 160664 73902 160784 73930
rect 160204 64870 160232 67606
rect 160192 64864 160244 64870
rect 160192 64806 160244 64812
rect 160664 39574 160692 73902
rect 160744 72888 160796 72894
rect 160744 72830 160796 72836
rect 160756 67634 160784 72830
rect 160940 71774 160968 79716
rect 161020 79688 161072 79694
rect 161020 79630 161072 79636
rect 161032 74526 161060 79630
rect 161110 79520 161166 79529
rect 161110 79455 161166 79464
rect 161020 74520 161072 74526
rect 161020 74462 161072 74468
rect 160940 71746 161060 71774
rect 161032 71398 161060 71746
rect 161020 71392 161072 71398
rect 161020 71334 161072 71340
rect 160756 67606 160968 67634
rect 160652 39568 160704 39574
rect 160652 39510 160704 39516
rect 160940 32570 160968 67606
rect 160928 32564 160980 32570
rect 160928 32506 160980 32512
rect 160098 30968 160154 30977
rect 160098 30903 160154 30912
rect 160008 11960 160060 11966
rect 160008 11902 160060 11908
rect 159640 10464 159692 10470
rect 159640 10406 159692 10412
rect 158904 4820 158956 4826
rect 158904 4762 158956 4768
rect 158916 480 158944 4762
rect 160112 480 160140 30903
rect 161032 15978 161060 71334
rect 161124 22982 161152 79455
rect 161216 78577 161244 79766
rect 161296 79756 161348 79762
rect 161538 79778 161566 80036
rect 161630 79937 161658 80036
rect 161722 79966 161750 80036
rect 161710 79960 161762 79966
rect 161616 79928 161672 79937
rect 161710 79902 161762 79908
rect 161616 79863 161672 79872
rect 161664 79824 161716 79830
rect 161538 79750 161612 79778
rect 161664 79766 161716 79772
rect 161814 79778 161842 80036
rect 161906 79898 161934 80036
rect 161998 79966 162026 80036
rect 162090 79966 162118 80036
rect 161986 79960 162038 79966
rect 161986 79902 162038 79908
rect 162078 79960 162130 79966
rect 162078 79902 162130 79908
rect 161894 79892 161946 79898
rect 161894 79834 161946 79840
rect 162182 79812 162210 80036
rect 162274 79966 162302 80036
rect 162262 79960 162314 79966
rect 162262 79902 162314 79908
rect 161984 79792 162040 79801
rect 161432 79727 161488 79736
rect 161296 79698 161348 79704
rect 161202 78568 161258 78577
rect 161202 78503 161258 78512
rect 161202 78296 161258 78305
rect 161308 78282 161336 79698
rect 161386 79656 161442 79665
rect 161386 79591 161442 79600
rect 161258 78254 161336 78282
rect 161202 78231 161258 78240
rect 161112 22976 161164 22982
rect 161112 22918 161164 22924
rect 161216 20058 161244 78231
rect 161296 74384 161348 74390
rect 161296 74326 161348 74332
rect 161204 20052 161256 20058
rect 161204 19994 161256 20000
rect 161308 16046 161336 74326
rect 161400 71330 161428 79591
rect 161584 77246 161612 79750
rect 161572 77240 161624 77246
rect 161572 77182 161624 77188
rect 161676 75818 161704 79766
rect 161814 79750 161888 79778
rect 161754 79656 161810 79665
rect 161754 79591 161810 79600
rect 161768 79014 161796 79591
rect 161756 79008 161808 79014
rect 161756 78950 161808 78956
rect 161664 75812 161716 75818
rect 161664 75754 161716 75760
rect 161480 74520 161532 74526
rect 161480 74462 161532 74468
rect 161388 71324 161440 71330
rect 161388 71266 161440 71272
rect 161296 16040 161348 16046
rect 161296 15982 161348 15988
rect 161020 15972 161072 15978
rect 161020 15914 161072 15920
rect 161400 9178 161428 71266
rect 161492 68950 161520 74462
rect 161860 72010 161888 79750
rect 162136 79784 162210 79812
rect 162136 79778 162164 79784
rect 162040 79750 162164 79778
rect 161984 79727 162040 79736
rect 161940 79688 161992 79694
rect 162366 79676 162394 80036
rect 162458 79778 162486 80036
rect 162550 79898 162578 80036
rect 162538 79892 162590 79898
rect 162538 79834 162590 79840
rect 162642 79778 162670 80036
rect 162734 79971 162762 80036
rect 162720 79962 162776 79971
rect 162720 79897 162776 79906
rect 162826 79898 162854 80036
rect 162814 79892 162866 79898
rect 162814 79834 162866 79840
rect 162918 79778 162946 80036
rect 163010 79898 163038 80036
rect 163102 79937 163130 80036
rect 163088 79928 163144 79937
rect 162998 79892 163050 79898
rect 163194 79898 163222 80036
rect 163286 79966 163314 80036
rect 163274 79960 163326 79966
rect 163274 79902 163326 79908
rect 163378 79898 163406 80036
rect 163470 79966 163498 80036
rect 163458 79960 163510 79966
rect 163562 79937 163590 80036
rect 163458 79902 163510 79908
rect 163548 79928 163604 79937
rect 163088 79863 163144 79872
rect 163182 79892 163234 79898
rect 162998 79834 163050 79840
rect 163182 79834 163234 79840
rect 163366 79892 163418 79898
rect 163548 79863 163604 79872
rect 163366 79834 163418 79840
rect 163318 79792 163374 79801
rect 162458 79750 162532 79778
rect 162642 79750 162716 79778
rect 162918 79750 163084 79778
rect 161940 79630 161992 79636
rect 162214 79656 162270 79665
rect 161952 78470 161980 79630
rect 162032 79620 162084 79626
rect 162214 79591 162270 79600
rect 162320 79648 162394 79676
rect 162504 79665 162532 79750
rect 162584 79688 162636 79694
rect 162490 79656 162546 79665
rect 162032 79562 162084 79568
rect 162044 78742 162072 79562
rect 162124 79552 162176 79558
rect 162124 79494 162176 79500
rect 162032 78736 162084 78742
rect 162032 78678 162084 78684
rect 161940 78464 161992 78470
rect 161940 78406 161992 78412
rect 162136 77042 162164 79494
rect 162228 79150 162256 79591
rect 162216 79144 162268 79150
rect 162216 79086 162268 79092
rect 162320 78928 162348 79648
rect 162584 79630 162636 79636
rect 162490 79591 162546 79600
rect 162492 79552 162544 79558
rect 162398 79520 162454 79529
rect 162492 79494 162544 79500
rect 162398 79455 162454 79464
rect 162412 79422 162440 79455
rect 162400 79416 162452 79422
rect 162400 79358 162452 79364
rect 162228 78900 162348 78928
rect 162124 77036 162176 77042
rect 162124 76978 162176 76984
rect 162032 75336 162084 75342
rect 162032 75278 162084 75284
rect 161848 72004 161900 72010
rect 161848 71946 161900 71952
rect 161480 68944 161532 68950
rect 161480 68886 161532 68892
rect 162044 43518 162072 75278
rect 162122 73128 162178 73137
rect 162122 73063 162178 73072
rect 162136 72457 162164 73063
rect 162122 72448 162178 72457
rect 162228 72418 162256 78900
rect 162400 78464 162452 78470
rect 162400 78406 162452 78412
rect 162412 75426 162440 78406
rect 162504 77081 162532 79494
rect 162596 79393 162624 79630
rect 162582 79384 162638 79393
rect 162582 79319 162638 79328
rect 162584 79144 162636 79150
rect 162584 79086 162636 79092
rect 162490 77072 162546 77081
rect 162490 77007 162546 77016
rect 162490 76936 162546 76945
rect 162490 76871 162546 76880
rect 162320 75398 162440 75426
rect 162122 72383 162178 72392
rect 162216 72412 162268 72418
rect 162216 72354 162268 72360
rect 162124 55888 162176 55894
rect 162124 55830 162176 55836
rect 162032 43512 162084 43518
rect 162032 43454 162084 43460
rect 161388 9172 161440 9178
rect 161388 9114 161440 9120
rect 161294 8936 161350 8945
rect 161294 8871 161350 8880
rect 161308 480 161336 8871
rect 162136 3398 162164 55830
rect 162228 33930 162256 72354
rect 162216 33924 162268 33930
rect 162216 33866 162268 33872
rect 162320 29782 162348 75398
rect 162400 72004 162452 72010
rect 162400 71946 162452 71952
rect 162412 71262 162440 71946
rect 162400 71256 162452 71262
rect 162400 71198 162452 71204
rect 162308 29776 162360 29782
rect 162308 29718 162360 29724
rect 162412 7750 162440 71198
rect 162504 11898 162532 76871
rect 162492 11892 162544 11898
rect 162492 11834 162544 11840
rect 162596 9110 162624 79086
rect 162688 76945 162716 79750
rect 162860 79688 162912 79694
rect 162860 79630 162912 79636
rect 162768 79416 162820 79422
rect 162768 79358 162820 79364
rect 162780 77466 162808 79358
rect 162872 77625 162900 79630
rect 162952 79484 163004 79490
rect 162952 79426 163004 79432
rect 162964 78130 162992 79426
rect 162952 78124 163004 78130
rect 162952 78066 163004 78072
rect 162964 77761 162992 78066
rect 162950 77752 163006 77761
rect 162950 77687 163006 77696
rect 162858 77616 162914 77625
rect 162858 77551 162914 77560
rect 162952 77512 163004 77518
rect 162780 77438 162900 77466
rect 162952 77454 163004 77460
rect 162768 77036 162820 77042
rect 162768 76978 162820 76984
rect 162674 76936 162730 76945
rect 162674 76871 162730 76880
rect 162780 76276 162808 76978
rect 162688 76248 162808 76276
rect 162584 9104 162636 9110
rect 162584 9046 162636 9052
rect 162400 7744 162452 7750
rect 162400 7686 162452 7692
rect 162688 5030 162716 76248
rect 162768 75812 162820 75818
rect 162768 75754 162820 75760
rect 162676 5024 162728 5030
rect 162676 4966 162728 4972
rect 162780 3738 162808 75754
rect 162872 60722 162900 77438
rect 162964 62082 162992 77454
rect 163056 77178 163084 79750
rect 163562 79778 163590 79863
rect 163654 79830 163682 80036
rect 163746 79898 163774 80036
rect 163838 79966 163866 80036
rect 163826 79960 163878 79966
rect 163826 79902 163878 79908
rect 163734 79892 163786 79898
rect 163734 79834 163786 79840
rect 163318 79727 163374 79736
rect 163424 79750 163590 79778
rect 163642 79824 163694 79830
rect 163930 79801 163958 80036
rect 163642 79766 163694 79772
rect 163916 79792 163972 79801
rect 163780 79756 163832 79762
rect 163136 79688 163188 79694
rect 163188 79648 163268 79676
rect 163136 79630 163188 79636
rect 163136 79552 163188 79558
rect 163136 79494 163188 79500
rect 163148 78985 163176 79494
rect 163134 78976 163190 78985
rect 163134 78911 163190 78920
rect 163136 78668 163188 78674
rect 163136 78610 163188 78616
rect 163044 77172 163096 77178
rect 163044 77114 163096 77120
rect 163148 67634 163176 78610
rect 163240 77314 163268 79648
rect 163332 77518 163360 79727
rect 163424 77994 163452 79750
rect 163916 79727 163972 79736
rect 163780 79698 163832 79704
rect 163596 79620 163648 79626
rect 163596 79562 163648 79568
rect 163502 79520 163558 79529
rect 163502 79455 163504 79464
rect 163556 79455 163558 79464
rect 163504 79426 163556 79432
rect 163412 77988 163464 77994
rect 163412 77930 163464 77936
rect 163320 77512 163372 77518
rect 163320 77454 163372 77460
rect 163320 77376 163372 77382
rect 163320 77318 163372 77324
rect 163228 77308 163280 77314
rect 163228 77250 163280 77256
rect 163056 67606 163176 67634
rect 163332 67634 163360 77318
rect 163608 73681 163636 79562
rect 163688 79552 163740 79558
rect 163688 79494 163740 79500
rect 163594 73672 163650 73681
rect 163594 73607 163650 73616
rect 163700 71466 163728 79494
rect 163792 78674 163820 79698
rect 164022 79676 164050 80036
rect 164114 79898 164142 80036
rect 164206 79937 164234 80036
rect 164192 79928 164248 79937
rect 164102 79892 164154 79898
rect 164192 79863 164248 79872
rect 164102 79834 164154 79840
rect 164148 79756 164200 79762
rect 164148 79698 164200 79704
rect 163976 79648 164050 79676
rect 163780 78668 163832 78674
rect 163780 78610 163832 78616
rect 163778 78568 163834 78577
rect 163778 78503 163834 78512
rect 163688 71460 163740 71466
rect 163688 71402 163740 71408
rect 163792 67634 163820 78503
rect 163976 71806 164004 79648
rect 164056 79552 164108 79558
rect 164054 79520 164056 79529
rect 164108 79520 164110 79529
rect 164054 79455 164110 79464
rect 164160 77296 164188 79698
rect 164298 79676 164326 80036
rect 164390 79830 164418 80036
rect 164482 79898 164510 80036
rect 164470 79892 164522 79898
rect 164470 79834 164522 79840
rect 164378 79824 164430 79830
rect 164574 79778 164602 80036
rect 164666 79830 164694 80036
rect 164378 79766 164430 79772
rect 164528 79750 164602 79778
rect 164654 79824 164706 79830
rect 164758 79801 164786 80036
rect 164654 79766 164706 79772
rect 164744 79792 164800 79801
rect 164252 79648 164326 79676
rect 164424 79688 164476 79694
rect 164252 78946 164280 79648
rect 164424 79630 164476 79636
rect 164240 78940 164292 78946
rect 164240 78882 164292 78888
rect 164332 78668 164384 78674
rect 164332 78610 164384 78616
rect 164160 77268 164280 77296
rect 164146 77208 164202 77217
rect 164146 77143 164202 77152
rect 163964 71800 164016 71806
rect 164016 71748 164096 71774
rect 163964 71746 164096 71748
rect 163964 71742 164016 71746
rect 163964 71460 164016 71466
rect 163964 71402 164016 71408
rect 163332 67606 163452 67634
rect 163792 67606 163912 67634
rect 163056 67522 163084 67606
rect 163044 67516 163096 67522
rect 163044 67458 163096 67464
rect 162952 62076 163004 62082
rect 162952 62018 163004 62024
rect 162860 60716 162912 60722
rect 162860 60658 162912 60664
rect 163424 33998 163452 67606
rect 163412 33992 163464 33998
rect 163412 33934 163464 33940
rect 163884 28422 163912 67606
rect 163872 28416 163924 28422
rect 163872 28358 163924 28364
rect 163976 14618 164004 71402
rect 163964 14612 164016 14618
rect 163964 14554 164016 14560
rect 164068 13190 164096 71746
rect 164160 14550 164188 77143
rect 164252 72214 164280 77268
rect 164240 72208 164292 72214
rect 164240 72150 164292 72156
rect 164240 72072 164292 72078
rect 164240 72014 164292 72020
rect 164252 31210 164280 72014
rect 164344 71738 164372 78610
rect 164332 71732 164384 71738
rect 164332 71674 164384 71680
rect 164436 70394 164464 79630
rect 164528 78674 164556 79750
rect 164744 79727 164800 79736
rect 164608 79688 164660 79694
rect 164850 79676 164878 80036
rect 164942 79937 164970 80036
rect 165034 79966 165062 80036
rect 165126 79966 165154 80036
rect 165022 79960 165074 79966
rect 164928 79928 164984 79937
rect 165022 79902 165074 79908
rect 165114 79960 165166 79966
rect 165114 79902 165166 79908
rect 164928 79863 164984 79872
rect 164942 79812 164970 79863
rect 165218 79830 165246 80036
rect 165310 79898 165338 80036
rect 165298 79892 165350 79898
rect 165298 79834 165350 79840
rect 165206 79824 165258 79830
rect 164942 79784 165016 79812
rect 164988 79744 165016 79784
rect 165402 79778 165430 80036
rect 165494 79937 165522 80036
rect 165480 79928 165536 79937
rect 165480 79863 165536 79872
rect 165586 79778 165614 80036
rect 165206 79766 165258 79772
rect 165356 79750 165430 79778
rect 165540 79750 165614 79778
rect 164988 79716 165108 79744
rect 164608 79630 164660 79636
rect 164712 79648 164878 79676
rect 164620 79393 164648 79630
rect 164606 79384 164662 79393
rect 164606 79319 164662 79328
rect 164516 78668 164568 78674
rect 164516 78610 164568 78616
rect 164620 77790 164648 79319
rect 164608 77784 164660 77790
rect 164608 77726 164660 77732
rect 164608 77648 164660 77654
rect 164608 77590 164660 77596
rect 164620 72078 164648 77590
rect 164712 73166 164740 79648
rect 164792 79552 164844 79558
rect 164792 79494 164844 79500
rect 164804 78169 164832 79494
rect 164976 79348 165028 79354
rect 164976 79290 165028 79296
rect 164884 79144 164936 79150
rect 164884 79086 164936 79092
rect 164790 78160 164846 78169
rect 164790 78095 164846 78104
rect 164792 78056 164844 78062
rect 164792 77998 164844 78004
rect 164804 75070 164832 77998
rect 164896 77654 164924 79086
rect 164988 79082 165016 79290
rect 164976 79076 165028 79082
rect 164976 79018 165028 79024
rect 164974 78432 165030 78441
rect 164974 78367 165030 78376
rect 164884 77648 164936 77654
rect 164884 77590 164936 77596
rect 164792 75064 164844 75070
rect 164792 75006 164844 75012
rect 164700 73160 164752 73166
rect 164700 73102 164752 73108
rect 164608 72072 164660 72078
rect 164608 72014 164660 72020
rect 164344 70366 164464 70394
rect 164344 69018 164372 70366
rect 164332 69012 164384 69018
rect 164332 68954 164384 68960
rect 164804 64874 164832 75006
rect 164804 64846 164924 64874
rect 164896 43450 164924 64846
rect 164884 43444 164936 43450
rect 164884 43386 164936 43392
rect 164988 38146 165016 78367
rect 165080 46306 165108 79716
rect 165160 79688 165212 79694
rect 165160 79630 165212 79636
rect 165172 79257 165200 79630
rect 165252 79620 165304 79626
rect 165252 79562 165304 79568
rect 165158 79248 165214 79257
rect 165158 79183 165214 79192
rect 165172 77654 165200 79183
rect 165264 78849 165292 79562
rect 165250 78840 165306 78849
rect 165250 78775 165306 78784
rect 165356 78520 165384 79750
rect 165436 79552 165488 79558
rect 165436 79494 165488 79500
rect 165264 78492 165384 78520
rect 165264 78033 165292 78492
rect 165342 78432 165398 78441
rect 165342 78367 165398 78376
rect 165250 78024 165306 78033
rect 165250 77959 165306 77968
rect 165160 77648 165212 77654
rect 165160 77590 165212 77596
rect 165252 73160 165304 73166
rect 165252 73102 165304 73108
rect 165160 71596 165212 71602
rect 165160 71538 165212 71544
rect 165068 46300 165120 46306
rect 165068 46242 165120 46248
rect 164976 38140 165028 38146
rect 164976 38082 165028 38088
rect 164240 31204 164292 31210
rect 164240 31146 164292 31152
rect 165172 27130 165200 71538
rect 165160 27124 165212 27130
rect 165160 27066 165212 27072
rect 165264 22914 165292 73102
rect 165252 22908 165304 22914
rect 165252 22850 165304 22856
rect 165356 17474 165384 78367
rect 165448 73681 165476 79494
rect 165540 78062 165568 79750
rect 165678 79676 165706 80036
rect 165770 79830 165798 80036
rect 165862 79937 165890 80036
rect 165954 79966 165982 80036
rect 165942 79960 165994 79966
rect 165848 79928 165904 79937
rect 165942 79902 165994 79908
rect 166046 79898 166074 80036
rect 166138 79966 166166 80036
rect 166126 79960 166178 79966
rect 166126 79902 166178 79908
rect 165848 79863 165904 79872
rect 166034 79892 166086 79898
rect 166034 79834 166086 79840
rect 165758 79824 165810 79830
rect 165758 79766 165810 79772
rect 165896 79824 165948 79830
rect 165896 79766 165948 79772
rect 166078 79792 166134 79801
rect 165678 79648 165752 79676
rect 165620 79552 165672 79558
rect 165620 79494 165672 79500
rect 165632 79150 165660 79494
rect 165620 79144 165672 79150
rect 165620 79086 165672 79092
rect 165620 78940 165672 78946
rect 165620 78882 165672 78888
rect 165528 78056 165580 78062
rect 165528 77998 165580 78004
rect 165434 73672 165490 73681
rect 165434 73607 165490 73616
rect 165528 72208 165580 72214
rect 165528 72150 165580 72156
rect 165436 71732 165488 71738
rect 165436 71674 165488 71680
rect 165448 71194 165476 71674
rect 165436 71188 165488 71194
rect 165436 71130 165488 71136
rect 165344 17468 165396 17474
rect 165344 17410 165396 17416
rect 164148 14544 164200 14550
rect 164148 14486 164200 14492
rect 164056 13184 164108 13190
rect 164056 13126 164108 13132
rect 165448 6254 165476 71130
rect 165540 6322 165568 72150
rect 165632 71602 165660 78882
rect 165724 75410 165752 79648
rect 165804 79620 165856 79626
rect 165804 79562 165856 79568
rect 165816 77858 165844 79562
rect 165804 77852 165856 77858
rect 165804 77794 165856 77800
rect 165712 75404 165764 75410
rect 165712 75346 165764 75352
rect 165908 74526 165936 79766
rect 166230 79744 166258 80036
rect 166322 79801 166350 80036
rect 166414 79966 166442 80036
rect 166506 79966 166534 80036
rect 166402 79960 166454 79966
rect 166402 79902 166454 79908
rect 166494 79960 166546 79966
rect 166598 79937 166626 80036
rect 166494 79902 166546 79908
rect 166584 79928 166640 79937
rect 166584 79863 166640 79872
rect 166078 79727 166134 79736
rect 166092 79676 166120 79727
rect 166000 79648 166120 79676
rect 166184 79716 166258 79744
rect 166308 79792 166364 79801
rect 166308 79727 166364 79736
rect 166000 79234 166028 79648
rect 166000 79206 166120 79234
rect 165988 75404 166040 75410
rect 165988 75346 166040 75352
rect 165896 74520 165948 74526
rect 165896 74462 165948 74468
rect 166000 71738 166028 75346
rect 166092 75342 166120 79206
rect 166080 75336 166132 75342
rect 166080 75278 166132 75284
rect 165988 71732 166040 71738
rect 165988 71674 166040 71680
rect 165620 71596 165672 71602
rect 165620 71538 165672 71544
rect 166184 70394 166212 79716
rect 166448 79688 166500 79694
rect 166598 79676 166626 79863
rect 166690 79778 166718 80036
rect 166782 79966 166810 80036
rect 166770 79960 166822 79966
rect 166770 79902 166822 79908
rect 166874 79898 166902 80036
rect 166966 79971 166994 80036
rect 166952 79962 167008 79971
rect 166862 79892 166914 79898
rect 166952 79897 167008 79906
rect 166862 79834 166914 79840
rect 166690 79750 166948 79778
rect 166598 79648 166672 79676
rect 166448 79630 166500 79636
rect 166356 79620 166408 79626
rect 166356 79562 166408 79568
rect 166264 77308 166316 77314
rect 166264 77250 166316 77256
rect 165908 70366 166212 70394
rect 165908 70174 165936 70366
rect 165896 70168 165948 70174
rect 165896 70110 165948 70116
rect 166276 60654 166304 77250
rect 166368 71874 166396 79562
rect 166460 78033 166488 79630
rect 166540 79484 166592 79490
rect 166540 79426 166592 79432
rect 166552 79257 166580 79426
rect 166538 79248 166594 79257
rect 166538 79183 166594 79192
rect 166446 78024 166502 78033
rect 166446 77959 166502 77968
rect 166552 72298 166580 79183
rect 166644 78928 166672 79648
rect 166816 79620 166868 79626
rect 166816 79562 166868 79568
rect 166644 78900 166764 78928
rect 166630 78840 166686 78849
rect 166630 78775 166686 78784
rect 166644 77926 166672 78775
rect 166632 77920 166684 77926
rect 166632 77862 166684 77868
rect 166736 77772 166764 78900
rect 166460 72270 166580 72298
rect 166644 77744 166764 77772
rect 166356 71868 166408 71874
rect 166356 71810 166408 71816
rect 166356 71732 166408 71738
rect 166356 71674 166408 71680
rect 166368 70922 166396 71674
rect 166356 70916 166408 70922
rect 166356 70858 166408 70864
rect 166264 60648 166316 60654
rect 166264 60590 166316 60596
rect 166368 40866 166396 70858
rect 166356 40860 166408 40866
rect 166356 40802 166408 40808
rect 166460 32502 166488 72270
rect 166540 70304 166592 70310
rect 166540 70246 166592 70252
rect 166552 69630 166580 70246
rect 166540 69624 166592 69630
rect 166540 69566 166592 69572
rect 166448 32496 166500 32502
rect 166448 32438 166500 32444
rect 166552 17406 166580 69566
rect 166644 21418 166672 77744
rect 166828 75936 166856 79562
rect 166920 75993 166948 79750
rect 167058 79744 167086 80036
rect 167150 79898 167178 80036
rect 167242 79966 167270 80036
rect 167230 79960 167282 79966
rect 167230 79902 167282 79908
rect 167138 79892 167190 79898
rect 167138 79834 167190 79840
rect 167334 79812 167362 80036
rect 167426 79898 167454 80036
rect 167518 79966 167546 80036
rect 167506 79960 167558 79966
rect 167506 79902 167558 79908
rect 167414 79892 167466 79898
rect 167414 79834 167466 79840
rect 167012 79716 167086 79744
rect 167288 79784 167362 79812
rect 166736 75908 166856 75936
rect 166906 75984 166962 75993
rect 166906 75919 166962 75928
rect 166736 70310 166764 75908
rect 167012 75274 167040 79716
rect 167092 79620 167144 79626
rect 167092 79562 167144 79568
rect 167000 75268 167052 75274
rect 167000 75210 167052 75216
rect 166816 74520 166868 74526
rect 166816 74462 166868 74468
rect 166724 70304 166776 70310
rect 166724 70246 166776 70252
rect 166724 70168 166776 70174
rect 166724 70110 166776 70116
rect 166632 21412 166684 21418
rect 166632 21354 166684 21360
rect 166540 17400 166592 17406
rect 166540 17342 166592 17348
rect 165620 17264 165672 17270
rect 165620 17206 165672 17212
rect 165632 16574 165660 17206
rect 165632 16546 166120 16574
rect 165528 6316 165580 6322
rect 165528 6258 165580 6264
rect 165436 6248 165488 6254
rect 165436 6190 165488 6196
rect 162768 3732 162820 3738
rect 162768 3674 162820 3680
rect 163688 3664 163740 3670
rect 163688 3606 163740 3612
rect 162492 3460 162544 3466
rect 162492 3402 162544 3408
rect 162124 3392 162176 3398
rect 162124 3334 162176 3340
rect 162504 480 162532 3402
rect 163700 480 163728 3606
rect 164884 3392 164936 3398
rect 164884 3334 164936 3340
rect 164896 480 164924 3334
rect 166092 480 166120 16546
rect 166736 11830 166764 70110
rect 166828 15910 166856 74462
rect 166908 71868 166960 71874
rect 166908 71810 166960 71816
rect 166920 70106 166948 71810
rect 166908 70100 166960 70106
rect 166908 70042 166960 70048
rect 166816 15904 166868 15910
rect 166816 15846 166868 15852
rect 166724 11824 166776 11830
rect 166724 11766 166776 11772
rect 166920 10402 166948 70042
rect 167104 59362 167132 79562
rect 167184 79552 167236 79558
rect 167184 79494 167236 79500
rect 167196 79393 167224 79494
rect 167182 79384 167238 79393
rect 167182 79319 167238 79328
rect 167196 78470 167224 79319
rect 167184 78464 167236 78470
rect 167184 78406 167236 78412
rect 167182 76528 167238 76537
rect 167182 76463 167238 76472
rect 167196 62014 167224 76463
rect 167288 75721 167316 79784
rect 167610 79778 167638 80036
rect 167702 79937 167730 80036
rect 167688 79928 167744 79937
rect 167794 79898 167822 80036
rect 167886 79966 167914 80036
rect 167978 79966 168006 80036
rect 167874 79960 167926 79966
rect 167874 79902 167926 79908
rect 167966 79960 168018 79966
rect 167966 79902 168018 79908
rect 167688 79863 167744 79872
rect 167782 79892 167834 79898
rect 167782 79834 167834 79840
rect 167460 79756 167512 79762
rect 167460 79698 167512 79704
rect 167564 79750 167638 79778
rect 167920 79824 167972 79830
rect 167920 79766 167972 79772
rect 167828 79756 167880 79762
rect 167472 79393 167500 79698
rect 167458 79384 167514 79393
rect 167458 79319 167514 79328
rect 167460 79008 167512 79014
rect 167460 78950 167512 78956
rect 167274 75712 167330 75721
rect 167274 75647 167330 75656
rect 167472 72486 167500 78950
rect 167564 75886 167592 79750
rect 167828 79698 167880 79704
rect 167644 79688 167696 79694
rect 167644 79630 167696 79636
rect 167734 79656 167790 79665
rect 167552 75880 167604 75886
rect 167552 75822 167604 75828
rect 167564 75410 167592 75822
rect 167552 75404 167604 75410
rect 167552 75346 167604 75352
rect 167460 72480 167512 72486
rect 167460 72422 167512 72428
rect 167656 67634 167684 79630
rect 167734 79591 167790 79600
rect 167748 68338 167776 79591
rect 167840 76129 167868 79698
rect 167826 76120 167882 76129
rect 167826 76055 167882 76064
rect 167932 75954 167960 79766
rect 168070 79744 168098 80036
rect 168162 79971 168190 80036
rect 168148 79962 168204 79971
rect 168148 79897 168204 79906
rect 168254 79778 168282 80036
rect 168024 79716 168098 79744
rect 168208 79750 168282 79778
rect 168346 79778 168374 80036
rect 168438 79937 168466 80036
rect 168530 79966 168558 80036
rect 168518 79960 168570 79966
rect 168424 79928 168480 79937
rect 168518 79902 168570 79908
rect 168424 79863 168480 79872
rect 168470 79792 168526 79801
rect 168346 79750 168420 79778
rect 167920 75948 167972 75954
rect 167920 75890 167972 75896
rect 168024 75857 168052 79716
rect 168208 79665 168236 79750
rect 168288 79688 168340 79694
rect 168194 79656 168250 79665
rect 168116 79614 168194 79642
rect 168010 75848 168066 75857
rect 168010 75783 168066 75792
rect 168116 75698 168144 79614
rect 168288 79630 168340 79636
rect 168194 79591 168250 79600
rect 168194 79384 168250 79393
rect 168194 79319 168250 79328
rect 167932 75670 168144 75698
rect 167736 68332 167788 68338
rect 167736 68274 167788 68280
rect 167656 67606 167868 67634
rect 167184 62008 167236 62014
rect 167184 61950 167236 61956
rect 167092 59356 167144 59362
rect 167092 59298 167144 59304
rect 167840 56574 167868 67606
rect 167828 56568 167880 56574
rect 167828 56510 167880 56516
rect 167000 43648 167052 43654
rect 167000 43590 167052 43596
rect 167012 16574 167040 43590
rect 167932 33862 167960 75670
rect 168012 75404 168064 75410
rect 168012 75346 168064 75352
rect 167920 33856 167972 33862
rect 167920 33798 167972 33804
rect 168024 29714 168052 75346
rect 168104 75268 168156 75274
rect 168104 75210 168156 75216
rect 168116 70378 168144 75210
rect 168104 70372 168156 70378
rect 168104 70314 168156 70320
rect 168012 29708 168064 29714
rect 168012 29650 168064 29656
rect 168116 17338 168144 70314
rect 168208 24274 168236 79319
rect 168300 79257 168328 79630
rect 168286 79248 168342 79257
rect 168286 79183 168342 79192
rect 168392 75993 168420 79750
rect 168622 79744 168650 80036
rect 168714 79971 168742 80036
rect 168700 79962 168756 79971
rect 168806 79966 168834 80036
rect 168700 79897 168756 79906
rect 168794 79960 168846 79966
rect 168794 79902 168846 79908
rect 168898 79812 168926 80036
rect 168470 79727 168526 79736
rect 168484 76634 168512 79727
rect 168576 79716 168650 79744
rect 168852 79784 168926 79812
rect 168472 76628 168524 76634
rect 168472 76570 168524 76576
rect 168378 75984 168434 75993
rect 168288 75948 168340 75954
rect 168378 75919 168434 75928
rect 168288 75890 168340 75896
rect 168300 70242 168328 75890
rect 168576 75562 168604 79716
rect 168748 79484 168800 79490
rect 168748 79426 168800 79432
rect 168484 75534 168604 75562
rect 168288 70236 168340 70242
rect 168288 70178 168340 70184
rect 168196 24268 168248 24274
rect 168196 24210 168248 24216
rect 168104 17332 168156 17338
rect 168104 17274 168156 17280
rect 167012 16546 167224 16574
rect 166908 10396 166960 10402
rect 166908 10338 166960 10344
rect 167196 480 167224 16546
rect 168300 9042 168328 70178
rect 168484 60734 168512 75534
rect 168656 75200 168708 75206
rect 168656 75142 168708 75148
rect 168564 74656 168616 74662
rect 168564 74598 168616 74604
rect 168392 60706 168512 60734
rect 168392 52426 168420 60706
rect 168576 57934 168604 74598
rect 168668 64802 168696 75142
rect 168760 74458 168788 79426
rect 168748 74452 168800 74458
rect 168748 74394 168800 74400
rect 168852 67634 168880 79784
rect 168990 79744 169018 80036
rect 169082 79966 169110 80036
rect 169070 79960 169122 79966
rect 169070 79902 169122 79908
rect 169174 79744 169202 80036
rect 168944 79716 169018 79744
rect 169128 79716 169202 79744
rect 168944 75954 168972 79716
rect 169022 79656 169078 79665
rect 169022 79591 169024 79600
rect 169076 79591 169078 79600
rect 169024 79562 169076 79568
rect 169036 78334 169064 79562
rect 169024 78328 169076 78334
rect 169024 78270 169076 78276
rect 168932 75948 168984 75954
rect 168932 75890 168984 75896
rect 169128 75206 169156 79716
rect 169266 79676 169294 80036
rect 169358 79966 169386 80036
rect 169346 79960 169398 79966
rect 169450 79937 169478 80036
rect 169542 79966 169570 80036
rect 169530 79960 169582 79966
rect 169346 79902 169398 79908
rect 169436 79928 169492 79937
rect 169530 79902 169582 79908
rect 169634 79898 169662 80036
rect 169726 79966 169754 80036
rect 169818 79971 169846 80036
rect 169714 79960 169766 79966
rect 169714 79902 169766 79908
rect 169804 79962 169860 79971
rect 169436 79863 169492 79872
rect 169622 79892 169674 79898
rect 169804 79897 169860 79906
rect 169910 79898 169938 80036
rect 169622 79834 169674 79840
rect 169898 79892 169950 79898
rect 169898 79834 169950 79840
rect 169574 79792 169630 79801
rect 169574 79727 169630 79736
rect 169220 79648 169294 79676
rect 169392 79688 169444 79694
rect 169390 79656 169392 79665
rect 169484 79688 169536 79694
rect 169444 79656 169446 79665
rect 169116 75200 169168 75206
rect 169116 75142 169168 75148
rect 169220 74662 169248 79648
rect 169484 79630 169536 79636
rect 169390 79591 169446 79600
rect 169392 79552 169444 79558
rect 169392 79494 169444 79500
rect 169404 79393 169432 79494
rect 169390 79384 169446 79393
rect 169390 79319 169446 79328
rect 169300 76628 169352 76634
rect 169300 76570 169352 76576
rect 169208 74656 169260 74662
rect 169208 74598 169260 74604
rect 168852 67606 169064 67634
rect 168656 64796 168708 64802
rect 168656 64738 168708 64744
rect 168564 57928 168616 57934
rect 168564 57870 168616 57876
rect 169036 55214 169064 67606
rect 169312 60734 169340 76570
rect 169404 73710 169432 79319
rect 169392 73704 169444 73710
rect 169392 73646 169444 73652
rect 169496 71398 169524 79630
rect 169588 79626 169616 79727
rect 169666 79656 169722 79665
rect 169576 79620 169628 79626
rect 170002 79642 170030 80036
rect 170094 79971 170122 80036
rect 170080 79962 170136 79971
rect 170080 79897 170136 79906
rect 170186 79898 170214 80036
rect 170278 79966 170306 80036
rect 170370 79966 170398 80036
rect 170266 79960 170318 79966
rect 170266 79902 170318 79908
rect 170358 79960 170410 79966
rect 170462 79937 170490 80036
rect 170358 79902 170410 79908
rect 170448 79928 170504 79937
rect 170174 79892 170226 79898
rect 170448 79863 170504 79872
rect 170174 79834 170226 79840
rect 170404 79824 170456 79830
rect 170126 79792 170182 79801
rect 170404 79766 170456 79772
rect 170126 79727 170128 79736
rect 170180 79727 170182 79736
rect 170128 79698 170180 79704
rect 170416 79665 170444 79766
rect 170554 79676 170582 80036
rect 170646 79830 170674 80036
rect 170738 79966 170766 80036
rect 170830 79966 170858 80036
rect 170922 79966 170950 80036
rect 170726 79960 170778 79966
rect 170726 79902 170778 79908
rect 170818 79960 170870 79966
rect 170818 79902 170870 79908
rect 170910 79960 170962 79966
rect 170910 79902 170962 79908
rect 170634 79824 170686 79830
rect 171014 79801 171042 80036
rect 171106 79830 171134 80036
rect 171094 79824 171146 79830
rect 170634 79766 170686 79772
rect 171000 79792 171056 79801
rect 171094 79766 171146 79772
rect 171198 79778 171226 80036
rect 171290 79898 171318 80036
rect 171382 79937 171410 80036
rect 171368 79928 171424 79937
rect 171278 79892 171330 79898
rect 171368 79863 171424 79872
rect 171278 79834 171330 79840
rect 171474 79778 171502 80036
rect 171566 79937 171594 80036
rect 171552 79928 171608 79937
rect 171658 79898 171686 80036
rect 171552 79863 171608 79872
rect 171646 79892 171698 79898
rect 171198 79750 171272 79778
rect 171000 79727 171056 79736
rect 170402 79656 170458 79665
rect 169666 79591 169722 79600
rect 169852 79620 169904 79626
rect 169576 79562 169628 79568
rect 169588 78062 169616 79562
rect 169576 78056 169628 78062
rect 169576 77998 169628 78004
rect 169576 75948 169628 75954
rect 169576 75890 169628 75896
rect 169484 71392 169536 71398
rect 169484 71334 169536 71340
rect 169220 60706 169340 60734
rect 169024 55208 169076 55214
rect 169024 55150 169076 55156
rect 168380 52420 168432 52426
rect 168380 52362 168432 52368
rect 169220 46238 169248 60706
rect 168380 46232 168432 46238
rect 168380 46174 168432 46180
rect 169208 46232 169260 46238
rect 169208 46174 169260 46180
rect 168288 9036 168340 9042
rect 168288 8978 168340 8984
rect 168392 3670 168420 46174
rect 169496 39506 169524 71334
rect 169588 70310 169616 75890
rect 169576 70304 169628 70310
rect 169576 70246 169628 70252
rect 169484 39500 169536 39506
rect 169484 39442 169536 39448
rect 168472 39364 168524 39370
rect 168472 39306 168524 39312
rect 168380 3664 168432 3670
rect 168380 3606 168432 3612
rect 168484 3482 168512 39306
rect 169588 28354 169616 70246
rect 169680 31142 169708 79591
rect 170002 79614 170260 79642
rect 169852 79562 169904 79568
rect 169760 79484 169812 79490
rect 169760 79426 169812 79432
rect 169772 79121 169800 79426
rect 169758 79112 169814 79121
rect 169758 79047 169814 79056
rect 169668 31136 169720 31142
rect 169668 31078 169720 31084
rect 169576 28348 169628 28354
rect 169576 28290 169628 28296
rect 169772 7682 169800 79047
rect 169864 76537 169892 79562
rect 170128 79552 170180 79558
rect 170128 79494 170180 79500
rect 169942 79248 169998 79257
rect 169942 79183 169998 79192
rect 169850 76528 169906 76537
rect 169850 76463 169906 76472
rect 169852 75948 169904 75954
rect 169852 75890 169904 75896
rect 169864 35290 169892 75890
rect 169956 58682 169984 79183
rect 170140 76158 170168 79494
rect 170232 78538 170260 79614
rect 170554 79648 170720 79676
rect 170402 79591 170458 79600
rect 170312 79280 170364 79286
rect 170312 79222 170364 79228
rect 170220 78532 170272 78538
rect 170220 78474 170272 78480
rect 170324 77518 170352 79222
rect 170312 77512 170364 77518
rect 170312 77454 170364 77460
rect 170128 76152 170180 76158
rect 170128 76094 170180 76100
rect 170416 60734 170444 79591
rect 170496 79552 170548 79558
rect 170496 79494 170548 79500
rect 170588 79552 170640 79558
rect 170588 79494 170640 79500
rect 170508 78985 170536 79494
rect 170600 79393 170628 79494
rect 170586 79384 170642 79393
rect 170586 79319 170642 79328
rect 170494 78976 170550 78985
rect 170494 78911 170550 78920
rect 170048 60706 170444 60734
rect 169944 58676 169996 58682
rect 169944 58618 169996 58624
rect 170048 38078 170076 60706
rect 170036 38072 170088 38078
rect 170036 38014 170088 38020
rect 170404 36576 170456 36582
rect 170404 36518 170456 36524
rect 169852 35284 169904 35290
rect 169852 35226 169904 35232
rect 169760 7676 169812 7682
rect 169760 7618 169812 7624
rect 169576 3664 169628 3670
rect 169576 3606 169628 3612
rect 168392 3454 168512 3482
rect 168392 480 168420 3454
rect 169588 480 169616 3606
rect 170416 3330 170444 36518
rect 170508 33794 170536 78911
rect 170600 75954 170628 79319
rect 170692 78418 170720 79648
rect 171140 79620 171192 79626
rect 171140 79562 171192 79568
rect 170956 79552 171008 79558
rect 170956 79494 171008 79500
rect 170968 79257 170996 79494
rect 171048 79484 171100 79490
rect 171048 79426 171100 79432
rect 170954 79248 171010 79257
rect 170772 79212 170824 79218
rect 170954 79183 171010 79192
rect 170772 79154 170824 79160
rect 170784 78606 170812 79154
rect 170772 78600 170824 78606
rect 170772 78542 170824 78548
rect 170692 78390 170904 78418
rect 170876 76498 170904 78390
rect 170864 76492 170916 76498
rect 170864 76434 170916 76440
rect 170680 76424 170732 76430
rect 170680 76366 170732 76372
rect 170692 76158 170720 76366
rect 170772 76356 170824 76362
rect 170772 76298 170824 76304
rect 170680 76152 170732 76158
rect 170784 76129 170812 76298
rect 170680 76094 170732 76100
rect 170770 76120 170826 76129
rect 170588 75948 170640 75954
rect 170588 75890 170640 75896
rect 170692 49026 170720 76094
rect 170770 76055 170826 76064
rect 170680 49020 170732 49026
rect 170680 48962 170732 48968
rect 170784 39438 170812 76055
rect 170772 39432 170824 39438
rect 170772 39374 170824 39380
rect 170876 36718 170904 76434
rect 170864 36712 170916 36718
rect 170864 36654 170916 36660
rect 170496 33788 170548 33794
rect 170496 33730 170548 33736
rect 170968 17270 170996 79183
rect 170956 17264 171008 17270
rect 170956 17206 171008 17212
rect 171060 4894 171088 79426
rect 171152 71233 171180 79562
rect 171244 78946 171272 79750
rect 171428 79750 171502 79778
rect 171566 79778 171594 79863
rect 171646 79834 171698 79840
rect 171566 79750 171640 79778
rect 171322 79656 171378 79665
rect 171322 79591 171378 79600
rect 171232 78940 171284 78946
rect 171232 78882 171284 78888
rect 171244 76090 171272 78882
rect 171336 78849 171364 79591
rect 171428 79286 171456 79750
rect 171508 79688 171560 79694
rect 171508 79630 171560 79636
rect 171416 79280 171468 79286
rect 171416 79222 171468 79228
rect 171322 78840 171378 78849
rect 171322 78775 171378 78784
rect 171324 77308 171376 77314
rect 171324 77250 171376 77256
rect 171232 76084 171284 76090
rect 171232 76026 171284 76032
rect 171230 75984 171286 75993
rect 171230 75919 171286 75928
rect 171138 71224 171194 71233
rect 171138 71159 171194 71168
rect 171244 28286 171272 75919
rect 171336 29646 171364 77250
rect 171428 36650 171456 79222
rect 171520 78713 171548 79630
rect 171612 79218 171640 79750
rect 171750 79744 171778 80036
rect 171842 79966 171870 80036
rect 171830 79960 171882 79966
rect 171830 79902 171882 79908
rect 171704 79716 171778 79744
rect 171600 79212 171652 79218
rect 171600 79154 171652 79160
rect 171704 79121 171732 79716
rect 171934 79676 171962 80036
rect 172026 79801 172054 80036
rect 172012 79792 172068 79801
rect 172118 79778 172146 80036
rect 172210 79966 172238 80036
rect 172198 79960 172250 79966
rect 172198 79902 172250 79908
rect 172302 79898 172330 80036
rect 172394 79937 172422 80036
rect 172486 79966 172514 80036
rect 172474 79960 172526 79966
rect 172380 79928 172436 79937
rect 172290 79892 172342 79898
rect 172474 79902 172526 79908
rect 172380 79863 172436 79872
rect 172290 79834 172342 79840
rect 172428 79824 172480 79830
rect 172118 79750 172284 79778
rect 172428 79766 172480 79772
rect 172012 79727 172068 79736
rect 172060 79688 172112 79694
rect 171782 79656 171838 79665
rect 171934 79648 172008 79676
rect 171782 79591 171784 79600
rect 171836 79591 171838 79600
rect 171784 79562 171836 79568
rect 171796 79422 171824 79562
rect 171876 79552 171928 79558
rect 171876 79494 171928 79500
rect 171784 79416 171836 79422
rect 171784 79358 171836 79364
rect 171888 79286 171916 79494
rect 171876 79280 171928 79286
rect 171980 79257 172008 79648
rect 172060 79630 172112 79636
rect 171876 79222 171928 79228
rect 171966 79248 172022 79257
rect 171966 79183 172022 79192
rect 171690 79112 171746 79121
rect 171690 79047 171746 79056
rect 171506 78704 171562 78713
rect 171506 78639 171562 78648
rect 171520 75410 171548 78639
rect 171704 77314 171732 79047
rect 171968 78804 172020 78810
rect 171968 78746 172020 78752
rect 171980 78713 172008 78746
rect 171966 78704 172022 78713
rect 171966 78639 172022 78648
rect 171876 78192 171928 78198
rect 171876 78134 171928 78140
rect 171692 77308 171744 77314
rect 171692 77250 171744 77256
rect 171784 76696 171836 76702
rect 171784 76638 171836 76644
rect 171600 76084 171652 76090
rect 171600 76026 171652 76032
rect 171508 75404 171560 75410
rect 171508 75346 171560 75352
rect 171612 60734 171640 76026
rect 171796 76022 171824 76638
rect 171784 76016 171836 76022
rect 171784 75958 171836 75964
rect 171520 60706 171640 60734
rect 171520 42158 171548 60706
rect 171508 42152 171560 42158
rect 171508 42094 171560 42100
rect 171416 36644 171468 36650
rect 171416 36586 171468 36592
rect 171324 29640 171376 29646
rect 171324 29582 171376 29588
rect 171232 28280 171284 28286
rect 171232 28222 171284 28228
rect 171888 26994 171916 78134
rect 172072 75993 172100 79630
rect 172256 79393 172284 79750
rect 172336 79688 172388 79694
rect 172336 79630 172388 79636
rect 172242 79384 172298 79393
rect 172152 79348 172204 79354
rect 172242 79319 172298 79328
rect 172152 79290 172204 79296
rect 172058 75984 172114 75993
rect 172058 75919 172114 75928
rect 171968 75336 172020 75342
rect 171968 75278 172020 75284
rect 171980 70038 172008 75278
rect 172164 70281 172192 79290
rect 172348 79218 172376 79630
rect 172244 79212 172296 79218
rect 172244 79154 172296 79160
rect 172336 79212 172388 79218
rect 172336 79154 172388 79160
rect 172150 70272 172206 70281
rect 172150 70207 172206 70216
rect 171968 70032 172020 70038
rect 171968 69974 172020 69980
rect 171876 26988 171928 26994
rect 171876 26930 171928 26936
rect 171784 25560 171836 25566
rect 171784 25502 171836 25508
rect 171048 4888 171100 4894
rect 171048 4830 171100 4836
rect 170772 3800 170824 3806
rect 170772 3742 170824 3748
rect 170404 3324 170456 3330
rect 170404 3266 170456 3272
rect 170784 480 170812 3742
rect 171796 3534 171824 25502
rect 172256 14482 172284 79154
rect 172348 78198 172376 79154
rect 172336 78192 172388 78198
rect 172336 78134 172388 78140
rect 172334 78024 172390 78033
rect 172334 77959 172390 77968
rect 172244 14476 172296 14482
rect 172244 14418 172296 14424
rect 172348 13122 172376 77959
rect 172440 74361 172468 79766
rect 172578 79744 172606 80036
rect 172670 79830 172698 80036
rect 172762 79971 172790 80036
rect 172748 79962 172804 79971
rect 172748 79897 172804 79906
rect 172854 79898 172882 80036
rect 172946 79898 172974 80036
rect 173038 79966 173066 80036
rect 173026 79960 173078 79966
rect 173026 79902 173078 79908
rect 173130 79898 173158 80036
rect 173222 79898 173250 80036
rect 172842 79892 172894 79898
rect 172842 79834 172894 79840
rect 172934 79892 172986 79898
rect 172934 79834 172986 79840
rect 173118 79892 173170 79898
rect 173118 79834 173170 79840
rect 173210 79892 173262 79898
rect 173210 79834 173262 79840
rect 172658 79824 172710 79830
rect 173314 79778 173342 80036
rect 173406 79830 173434 80036
rect 172658 79766 172710 79772
rect 173176 79762 173342 79778
rect 173394 79824 173446 79830
rect 173498 79801 173526 80036
rect 173590 79966 173618 80036
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173682 79898 173710 80036
rect 173774 79971 173802 80036
rect 173760 79962 173816 79971
rect 173670 79892 173722 79898
rect 173760 79897 173816 79906
rect 173670 79834 173722 79840
rect 173394 79766 173446 79772
rect 173484 79792 173540 79801
rect 172532 79716 172606 79744
rect 172980 79756 173032 79762
rect 172532 79014 172560 79716
rect 172980 79698 173032 79704
rect 173072 79756 173124 79762
rect 173072 79698 173124 79704
rect 173164 79756 173342 79762
rect 173216 79750 173342 79756
rect 173484 79727 173540 79736
rect 173716 79756 173768 79762
rect 173164 79698 173216 79704
rect 172704 79688 172756 79694
rect 172610 79656 172666 79665
rect 172704 79630 172756 79636
rect 172888 79688 172940 79694
rect 172888 79630 172940 79636
rect 172610 79591 172666 79600
rect 172520 79008 172572 79014
rect 172520 78950 172572 78956
rect 172520 77308 172572 77314
rect 172520 77250 172572 77256
rect 172426 74352 172482 74361
rect 172426 74287 172482 74296
rect 172428 73908 172480 73914
rect 172428 73850 172480 73856
rect 172440 73817 172468 73850
rect 172426 73808 172482 73817
rect 172426 73743 172482 73752
rect 172336 13116 172388 13122
rect 172336 13058 172388 13064
rect 172440 3806 172468 73743
rect 172532 24206 172560 77250
rect 172624 32434 172652 79591
rect 172716 75857 172744 79630
rect 172796 79484 172848 79490
rect 172796 79426 172848 79432
rect 172808 76090 172836 79426
rect 172796 76084 172848 76090
rect 172796 76026 172848 76032
rect 172702 75848 172758 75857
rect 172702 75783 172758 75792
rect 172900 75274 172928 79630
rect 172992 79393 173020 79698
rect 172978 79384 173034 79393
rect 172978 79319 173034 79328
rect 172888 75268 172940 75274
rect 172888 75210 172940 75216
rect 172992 75206 173020 79319
rect 172980 75200 173032 75206
rect 173084 75177 173112 79698
rect 173164 79620 173216 79626
rect 173164 79562 173216 79568
rect 173256 79620 173308 79626
rect 173256 79562 173308 79568
rect 173348 79620 173400 79626
rect 173498 79608 173526 79727
rect 173716 79698 173768 79704
rect 173498 79580 173572 79608
rect 173348 79562 173400 79568
rect 173176 79286 173204 79562
rect 173268 79393 173296 79562
rect 173254 79384 173310 79393
rect 173254 79319 173310 79328
rect 173164 79280 173216 79286
rect 173164 79222 173216 79228
rect 173268 78402 173296 79319
rect 173360 78742 173388 79562
rect 173440 79484 173492 79490
rect 173440 79426 173492 79432
rect 173348 78736 173400 78742
rect 173348 78678 173400 78684
rect 173256 78396 173308 78402
rect 173256 78338 173308 78344
rect 173360 77314 173388 78678
rect 173348 77308 173400 77314
rect 173348 77250 173400 77256
rect 173452 76786 173480 79426
rect 173176 76758 173480 76786
rect 172980 75142 173032 75148
rect 173070 75168 173126 75177
rect 173070 75103 173126 75112
rect 173176 66162 173204 76758
rect 173346 76664 173402 76673
rect 173346 76599 173402 76608
rect 173360 67634 173388 76599
rect 173360 67606 173480 67634
rect 173164 66156 173216 66162
rect 173164 66098 173216 66104
rect 173452 40798 173480 67606
rect 173440 40792 173492 40798
rect 173440 40734 173492 40740
rect 173544 38010 173572 79580
rect 173624 79076 173676 79082
rect 173624 79018 173676 79024
rect 173636 77450 173664 79018
rect 173624 77444 173676 77450
rect 173624 77386 173676 77392
rect 173728 75449 173756 79698
rect 173866 79642 173894 80036
rect 173958 79830 173986 80036
rect 174050 79966 174078 80036
rect 174038 79960 174090 79966
rect 174038 79902 174090 79908
rect 174142 79903 174170 80036
rect 174128 79894 174184 79903
rect 173946 79824 173998 79830
rect 174128 79829 174184 79838
rect 173946 79766 173998 79772
rect 174234 79744 174262 80036
rect 174326 79966 174354 80036
rect 174418 79966 174446 80036
rect 174510 79971 174538 80036
rect 174314 79960 174366 79966
rect 174314 79902 174366 79908
rect 174406 79960 174458 79966
rect 174406 79902 174458 79908
rect 174496 79962 174552 79971
rect 174496 79897 174552 79906
rect 174602 79898 174630 80036
rect 174694 79971 174722 80036
rect 174680 79962 174736 79971
rect 174786 79966 174814 80036
rect 174590 79892 174642 79898
rect 174680 79897 174736 79906
rect 174774 79960 174826 79966
rect 174878 79937 174906 80036
rect 174774 79902 174826 79908
rect 174864 79928 174920 79937
rect 174864 79863 174920 79872
rect 174590 79834 174642 79840
rect 174728 79824 174780 79830
rect 174878 79812 174906 79863
rect 174728 79766 174780 79772
rect 174832 79784 174906 79812
rect 174360 79756 174412 79762
rect 174234 79716 174308 79744
rect 173992 79688 174044 79694
rect 173866 79614 173940 79642
rect 173992 79630 174044 79636
rect 174082 79656 174138 79665
rect 173912 79393 173940 79614
rect 173898 79384 173954 79393
rect 173898 79319 173954 79328
rect 173808 78396 173860 78402
rect 173808 78338 173860 78344
rect 173900 78396 173952 78402
rect 173900 78338 173952 78344
rect 173714 75440 173770 75449
rect 173714 75375 173770 75384
rect 173716 75268 173768 75274
rect 173716 75210 173768 75216
rect 173728 75002 173756 75210
rect 173716 74996 173768 75002
rect 173716 74938 173768 74944
rect 173532 38004 173584 38010
rect 173532 37946 173584 37952
rect 172612 32428 172664 32434
rect 172612 32370 172664 32376
rect 173728 25702 173756 74938
rect 173716 25696 173768 25702
rect 173716 25638 173768 25644
rect 172520 24200 172572 24206
rect 172520 24142 172572 24148
rect 173820 6186 173848 78338
rect 173912 47598 173940 78338
rect 174004 75313 174032 79630
rect 174082 79591 174084 79600
rect 174136 79591 174138 79600
rect 174084 79562 174136 79568
rect 174176 79416 174228 79422
rect 174176 79358 174228 79364
rect 174084 79008 174136 79014
rect 174084 78950 174136 78956
rect 174096 76673 174124 78950
rect 174082 76664 174138 76673
rect 174082 76599 174138 76608
rect 174188 75410 174216 79358
rect 174280 79082 174308 79716
rect 174360 79698 174412 79704
rect 174452 79756 174504 79762
rect 174452 79698 174504 79704
rect 174544 79756 174596 79762
rect 174544 79698 174596 79704
rect 174372 79665 174400 79698
rect 174358 79656 174414 79665
rect 174358 79591 174414 79600
rect 174372 79422 174400 79591
rect 174360 79416 174412 79422
rect 174360 79358 174412 79364
rect 174268 79076 174320 79082
rect 174268 79018 174320 79024
rect 174176 75404 174228 75410
rect 174176 75346 174228 75352
rect 173990 75304 174046 75313
rect 173990 75239 174046 75248
rect 174280 67634 174308 79018
rect 174358 78704 174414 78713
rect 174358 78639 174414 78648
rect 174372 75274 174400 78639
rect 174360 75268 174412 75274
rect 174360 75210 174412 75216
rect 174464 68785 174492 79698
rect 174556 79393 174584 79698
rect 174542 79384 174598 79393
rect 174542 79319 174598 79328
rect 174556 78402 174584 79319
rect 174740 79014 174768 79766
rect 174832 79694 174860 79784
rect 174970 79744 174998 80036
rect 175062 79966 175090 80036
rect 175050 79960 175102 79966
rect 175154 79937 175182 80036
rect 175246 79966 175274 80036
rect 175234 79960 175286 79966
rect 175050 79902 175102 79908
rect 175140 79928 175196 79937
rect 175234 79902 175286 79908
rect 175140 79863 175196 79872
rect 174924 79716 174998 79744
rect 175094 79792 175150 79801
rect 175094 79727 175150 79736
rect 174820 79688 174872 79694
rect 174924 79665 174952 79716
rect 174820 79630 174872 79636
rect 174910 79656 174966 79665
rect 174910 79591 174966 79600
rect 175004 79620 175056 79626
rect 175004 79562 175056 79568
rect 174820 79552 174872 79558
rect 174872 79512 174952 79540
rect 174820 79494 174872 79500
rect 174820 79416 174872 79422
rect 174820 79358 174872 79364
rect 174728 79008 174780 79014
rect 174728 78950 174780 78956
rect 174544 78396 174596 78402
rect 174544 78338 174596 78344
rect 174728 78396 174780 78402
rect 174728 78338 174780 78344
rect 174740 76566 174768 78338
rect 174544 76560 174596 76566
rect 174544 76502 174596 76508
rect 174728 76560 174780 76566
rect 174728 76502 174780 76508
rect 174450 68776 174506 68785
rect 174450 68711 174506 68720
rect 174280 67606 174400 67634
rect 174372 60734 174400 67606
rect 174004 60706 174400 60734
rect 173900 47592 173952 47598
rect 173900 47534 173952 47540
rect 174004 22846 174032 60706
rect 173992 22840 174044 22846
rect 173992 22782 174044 22788
rect 174556 11762 174584 76502
rect 174726 75304 174782 75313
rect 174726 75239 174782 75248
rect 174740 39370 174768 75239
rect 174832 42090 174860 79358
rect 174924 72282 174952 79512
rect 174912 72276 174964 72282
rect 174912 72218 174964 72224
rect 174820 42084 174872 42090
rect 174820 42026 174872 42032
rect 174728 39364 174780 39370
rect 174728 39306 174780 39312
rect 174924 26926 174952 72218
rect 174912 26920 174964 26926
rect 174912 26862 174964 26868
rect 175016 25634 175044 79562
rect 175108 79354 175136 79727
rect 175338 79676 175366 80036
rect 175430 79966 175458 80036
rect 175522 79966 175550 80036
rect 175418 79960 175470 79966
rect 175418 79902 175470 79908
rect 175510 79960 175562 79966
rect 175510 79902 175562 79908
rect 175464 79756 175516 79762
rect 175614 79744 175642 80036
rect 175706 79898 175734 80036
rect 175798 79966 175826 80036
rect 175786 79960 175838 79966
rect 175786 79902 175838 79908
rect 175694 79892 175746 79898
rect 175694 79834 175746 79840
rect 175464 79698 175516 79704
rect 175568 79716 175642 79744
rect 175740 79756 175792 79762
rect 175338 79648 175412 79676
rect 175188 79620 175240 79626
rect 175188 79562 175240 79568
rect 175096 79348 175148 79354
rect 175096 79290 175148 79296
rect 175200 79257 175228 79562
rect 175280 79552 175332 79558
rect 175280 79494 175332 79500
rect 175292 79422 175320 79494
rect 175280 79416 175332 79422
rect 175280 79358 175332 79364
rect 175186 79248 175242 79257
rect 175186 79183 175242 79192
rect 175096 79008 175148 79014
rect 175096 78950 175148 78956
rect 175108 74361 175136 78950
rect 175200 77081 175228 79183
rect 175292 78402 175320 79358
rect 175384 79014 175412 79648
rect 175372 79008 175424 79014
rect 175372 78950 175424 78956
rect 175280 78396 175332 78402
rect 175280 78338 175332 78344
rect 175280 78192 175332 78198
rect 175280 78134 175332 78140
rect 175186 77072 175242 77081
rect 175186 77007 175242 77016
rect 175186 76800 175242 76809
rect 175186 76735 175242 76744
rect 175094 74352 175150 74361
rect 175094 74287 175150 74296
rect 175004 25628 175056 25634
rect 175004 25570 175056 25576
rect 174544 11756 174596 11762
rect 174544 11698 174596 11704
rect 175108 7614 175136 74287
rect 175096 7608 175148 7614
rect 175096 7550 175148 7556
rect 173808 6180 173860 6186
rect 173808 6122 173860 6128
rect 175200 4826 175228 76735
rect 175292 10334 175320 78134
rect 175384 37942 175412 78950
rect 175476 75177 175504 79698
rect 175568 75721 175596 79716
rect 175890 79744 175918 80036
rect 175982 79971 176010 80036
rect 175968 79962 176024 79971
rect 176074 79966 176102 80036
rect 175968 79897 176024 79906
rect 176062 79960 176114 79966
rect 176166 79937 176194 80036
rect 176062 79902 176114 79908
rect 176152 79928 176208 79937
rect 176258 79898 176286 80036
rect 176152 79863 176208 79872
rect 176246 79892 176298 79898
rect 176246 79834 176298 79840
rect 176016 79824 176068 79830
rect 175740 79698 175792 79704
rect 175844 79716 175918 79744
rect 176014 79792 176016 79801
rect 176350 79801 176378 80036
rect 176068 79792 176070 79801
rect 176014 79727 176070 79736
rect 176198 79792 176254 79801
rect 176198 79727 176254 79736
rect 176336 79792 176392 79801
rect 176336 79727 176392 79736
rect 176442 79744 176470 80036
rect 176534 79898 176562 80036
rect 176522 79892 176574 79898
rect 176522 79834 176574 79840
rect 176626 79830 176654 80036
rect 176614 79824 176666 79830
rect 176614 79766 176666 79772
rect 176718 79744 176746 80036
rect 176810 79898 176838 80036
rect 176902 79898 176930 80036
rect 176798 79892 176850 79898
rect 176798 79834 176850 79840
rect 176890 79892 176942 79898
rect 176890 79834 176942 79840
rect 176994 79778 177022 80036
rect 177086 79898 177114 80036
rect 177074 79892 177126 79898
rect 177074 79834 177126 79840
rect 176856 79750 177022 79778
rect 175648 79620 175700 79626
rect 175648 79562 175700 79568
rect 175660 79393 175688 79562
rect 175646 79384 175702 79393
rect 175646 79319 175702 79328
rect 175660 78402 175688 79319
rect 175648 78396 175700 78402
rect 175648 78338 175700 78344
rect 175554 75712 175610 75721
rect 175554 75647 175610 75656
rect 175462 75168 175518 75177
rect 175462 75103 175518 75112
rect 175752 71774 175780 79698
rect 175844 77625 175872 79716
rect 176016 79688 176068 79694
rect 176016 79630 176068 79636
rect 176106 79656 176162 79665
rect 175924 79552 175976 79558
rect 175924 79494 175976 79500
rect 175936 79393 175964 79494
rect 175922 79384 175978 79393
rect 175922 79319 175978 79328
rect 175830 77616 175886 77625
rect 175830 77551 175886 77560
rect 175830 77344 175886 77353
rect 175830 77279 175886 77288
rect 175660 71746 175780 71774
rect 175660 67454 175688 71746
rect 175844 69970 175872 77279
rect 175832 69964 175884 69970
rect 175832 69906 175884 69912
rect 175648 67448 175700 67454
rect 175648 67390 175700 67396
rect 175372 37936 175424 37942
rect 175372 37878 175424 37884
rect 175936 18698 175964 79319
rect 176028 77586 176056 79630
rect 176106 79591 176162 79600
rect 176120 79490 176148 79591
rect 176108 79484 176160 79490
rect 176108 79426 176160 79432
rect 176212 78849 176240 79727
rect 176442 79716 176516 79744
rect 176718 79716 176792 79744
rect 176382 79656 176438 79665
rect 176382 79591 176384 79600
rect 176436 79591 176438 79600
rect 176384 79562 176436 79568
rect 176292 79484 176344 79490
rect 176292 79426 176344 79432
rect 176198 78840 176254 78849
rect 176198 78775 176254 78784
rect 176108 78396 176160 78402
rect 176108 78338 176160 78344
rect 176016 77580 176068 77586
rect 176016 77522 176068 77528
rect 176120 53106 176148 78338
rect 176212 78198 176240 78775
rect 176304 78606 176332 79426
rect 176292 78600 176344 78606
rect 176292 78542 176344 78548
rect 176396 78418 176424 79562
rect 176304 78390 176424 78418
rect 176200 78192 176252 78198
rect 176200 78134 176252 78140
rect 176198 77616 176254 77625
rect 176198 77551 176254 77560
rect 176212 73778 176240 77551
rect 176200 73772 176252 73778
rect 176200 73714 176252 73720
rect 176108 53100 176160 53106
rect 176108 53042 176160 53048
rect 176212 36582 176240 73714
rect 176200 36576 176252 36582
rect 176200 36518 176252 36524
rect 176304 24138 176332 78390
rect 176384 77580 176436 77586
rect 176384 77522 176436 77528
rect 176292 24132 176344 24138
rect 176292 24074 176344 24080
rect 176396 18766 176424 77522
rect 176488 77081 176516 79716
rect 176658 79656 176714 79665
rect 176568 79620 176620 79626
rect 176658 79591 176714 79600
rect 176568 79562 176620 79568
rect 176580 77217 176608 79562
rect 176566 77208 176622 77217
rect 176566 77143 176622 77152
rect 176474 77072 176530 77081
rect 176474 77007 176530 77016
rect 176566 75712 176622 75721
rect 176566 75647 176622 75656
rect 176384 18760 176436 18766
rect 176384 18702 176436 18708
rect 175924 18692 175976 18698
rect 175924 18634 175976 18640
rect 175922 18592 175978 18601
rect 175922 18527 175978 18536
rect 175280 10328 175332 10334
rect 175280 10270 175332 10276
rect 175188 4820 175240 4826
rect 175188 4762 175240 4768
rect 172428 3800 172480 3806
rect 172428 3742 172480 3748
rect 175464 3596 175516 3602
rect 175464 3538 175516 3544
rect 171784 3528 171836 3534
rect 171784 3470 171836 3476
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 171966 3360 172022 3369
rect 171966 3295 172022 3304
rect 171980 480 172008 3295
rect 173176 480 173204 3470
rect 174268 3324 174320 3330
rect 174268 3266 174320 3272
rect 174280 480 174308 3266
rect 175476 480 175504 3538
rect 175936 3058 175964 18527
rect 176580 8974 176608 75647
rect 176672 51746 176700 79591
rect 176764 79257 176792 79716
rect 176750 79248 176806 79257
rect 176750 79183 176806 79192
rect 176752 78668 176804 78674
rect 176752 78610 176804 78616
rect 176764 68814 176792 78610
rect 176856 77897 176884 79750
rect 177178 79744 177206 80036
rect 177270 79812 177298 80036
rect 177362 79937 177390 80036
rect 177348 79928 177404 79937
rect 177348 79863 177404 79872
rect 177454 79880 177482 80036
rect 177546 79948 177574 80036
rect 177672 79960 177724 79966
rect 177546 79937 177620 79948
rect 177546 79928 177634 79937
rect 177546 79920 177578 79928
rect 177454 79852 177528 79880
rect 177672 79902 177724 79908
rect 177578 79863 177634 79872
rect 177270 79784 177436 79812
rect 177500 79801 177528 79852
rect 177178 79716 177252 79744
rect 176936 79688 176988 79694
rect 176936 79630 176988 79636
rect 177028 79688 177080 79694
rect 177028 79630 177080 79636
rect 176842 77888 176898 77897
rect 176842 77823 176898 77832
rect 176844 77580 176896 77586
rect 176844 77522 176896 77528
rect 176856 77081 176884 77522
rect 176842 77072 176898 77081
rect 176842 77007 176898 77016
rect 176856 74934 176884 77007
rect 176844 74928 176896 74934
rect 176844 74870 176896 74876
rect 176752 68808 176804 68814
rect 176752 68750 176804 68756
rect 176948 56438 176976 79630
rect 177040 78169 177068 79630
rect 177120 79620 177172 79626
rect 177120 79562 177172 79568
rect 177026 78160 177082 78169
rect 177026 78095 177082 78104
rect 177040 76226 177068 78095
rect 177132 77586 177160 79562
rect 177224 78674 177252 79716
rect 177302 79248 177358 79257
rect 177302 79183 177358 79192
rect 177212 78668 177264 78674
rect 177212 78610 177264 78616
rect 177120 77580 177172 77586
rect 177120 77522 177172 77528
rect 177028 76220 177080 76226
rect 177028 76162 177080 76168
rect 177212 76084 177264 76090
rect 177212 76026 177264 76032
rect 177224 71505 177252 76026
rect 177210 71496 177266 71505
rect 177210 71431 177266 71440
rect 176936 56432 176988 56438
rect 176936 56374 176988 56380
rect 176660 51740 176712 51746
rect 176660 51682 176712 51688
rect 177316 40730 177344 79183
rect 177408 77625 177436 79784
rect 177486 79792 177542 79801
rect 177486 79727 177542 79736
rect 177488 79348 177540 79354
rect 177488 79290 177540 79296
rect 177394 77616 177450 77625
rect 177394 77551 177450 77560
rect 177304 40724 177356 40730
rect 177304 40666 177356 40672
rect 177408 35222 177436 77551
rect 177500 75177 177528 79290
rect 177592 78577 177620 79863
rect 177684 78606 177712 79902
rect 177776 79354 177804 80174
rect 177868 79966 177896 80174
rect 177856 79960 177908 79966
rect 177856 79902 177908 79908
rect 177854 79792 177910 79801
rect 177854 79727 177910 79736
rect 177764 79348 177816 79354
rect 177764 79290 177816 79296
rect 177672 78600 177724 78606
rect 177578 78568 177634 78577
rect 177672 78542 177724 78548
rect 177578 78503 177634 78512
rect 177670 77888 177726 77897
rect 177670 77823 177726 77832
rect 177486 75168 177542 75177
rect 177486 75103 177542 75112
rect 177396 35216 177448 35222
rect 177396 35158 177448 35164
rect 177684 31074 177712 77823
rect 177764 76968 177816 76974
rect 177764 76910 177816 76916
rect 177776 75954 177804 76910
rect 177764 75948 177816 75954
rect 177764 75890 177816 75896
rect 177764 74928 177816 74934
rect 177764 74870 177816 74876
rect 177672 31068 177724 31074
rect 177672 31010 177724 31016
rect 177776 25566 177804 74870
rect 177764 25560 177816 25566
rect 177764 25502 177816 25508
rect 177868 22778 177896 79727
rect 177960 76974 177988 80566
rect 178052 79257 178080 80650
rect 178130 80608 178186 80617
rect 178130 80543 178186 80552
rect 178144 79422 178172 80543
rect 178420 80238 178448 80679
rect 182546 80679 182602 80688
rect 178592 80650 178644 80656
rect 178498 80336 178554 80345
rect 178498 80271 178554 80280
rect 178408 80232 178460 80238
rect 178408 80174 178460 80180
rect 178316 80164 178368 80170
rect 178316 80106 178368 80112
rect 178328 79422 178356 80106
rect 178132 79416 178184 79422
rect 178132 79358 178184 79364
rect 178316 79416 178368 79422
rect 178316 79358 178368 79364
rect 178038 79248 178094 79257
rect 178038 79183 178094 79192
rect 178222 78704 178278 78713
rect 178222 78639 178278 78648
rect 178038 78432 178094 78441
rect 178236 78418 178264 78639
rect 178314 78432 178370 78441
rect 178236 78390 178314 78418
rect 178038 78367 178094 78376
rect 178512 78402 178540 80271
rect 178604 80238 178632 80650
rect 178776 80368 178828 80374
rect 178776 80310 178828 80316
rect 178592 80232 178644 80238
rect 178592 80174 178644 80180
rect 178592 80028 178644 80034
rect 178592 79970 178644 79976
rect 178314 78367 178370 78376
rect 178500 78396 178552 78402
rect 178052 77450 178080 78367
rect 178500 78338 178552 78344
rect 178604 77489 178632 79970
rect 178682 79520 178738 79529
rect 178682 79455 178738 79464
rect 178590 77480 178646 77489
rect 178040 77444 178092 77450
rect 178590 77415 178646 77424
rect 178040 77386 178092 77392
rect 177948 76968 178000 76974
rect 177948 76910 178000 76916
rect 177948 76220 178000 76226
rect 177948 76162 178000 76168
rect 177856 22772 177908 22778
rect 177856 22714 177908 22720
rect 177960 18630 177988 76162
rect 177948 18624 178000 18630
rect 177948 18566 178000 18572
rect 178052 16574 178080 77386
rect 178052 16546 178632 16574
rect 176568 8968 176620 8974
rect 176568 8910 176620 8916
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 175924 3052 175976 3058
rect 175924 2994 175976 3000
rect 176672 480 176700 3334
rect 177856 3052 177908 3058
rect 177856 2994 177908 3000
rect 177868 480 177896 2994
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3670 178724 79455
rect 178788 78606 178816 80310
rect 182560 80238 182588 80679
rect 185214 80336 185270 80345
rect 185214 80271 185216 80280
rect 185268 80271 185270 80280
rect 185216 80242 185268 80248
rect 182548 80232 182600 80238
rect 182548 80174 182600 80180
rect 185228 80170 185256 80242
rect 185216 80164 185268 80170
rect 185216 80106 185268 80112
rect 182180 79484 182232 79490
rect 182180 79426 182232 79432
rect 178866 78704 178922 78713
rect 178866 78639 178922 78648
rect 178776 78600 178828 78606
rect 178776 78542 178828 78548
rect 178776 77784 178828 77790
rect 178776 77726 178828 77732
rect 178788 21486 178816 77726
rect 178880 77518 178908 78639
rect 179420 78260 179472 78266
rect 179420 78202 179472 78208
rect 178868 77512 178920 77518
rect 178868 77454 178920 77460
rect 178880 62898 178908 77454
rect 179432 77353 179460 78202
rect 181628 77920 181680 77926
rect 181628 77862 181680 77868
rect 180708 77852 180760 77858
rect 180708 77794 180760 77800
rect 180156 77648 180208 77654
rect 180156 77590 180208 77596
rect 179418 77344 179474 77353
rect 179418 77279 179474 77288
rect 179878 77208 179934 77217
rect 179878 77143 179934 77152
rect 179892 76022 179920 77143
rect 180064 76968 180116 76974
rect 180064 76910 180116 76916
rect 179880 76016 179932 76022
rect 179880 75958 179932 75964
rect 179420 69896 179472 69902
rect 179420 69838 179472 69844
rect 178868 62892 178920 62898
rect 178868 62834 178920 62840
rect 178776 21480 178828 21486
rect 178776 21422 178828 21428
rect 179432 16574 179460 69838
rect 179432 16546 180012 16574
rect 178684 3664 178736 3670
rect 178684 3606 178736 3612
rect 179984 3482 180012 16546
rect 180076 3602 180104 76910
rect 180168 4962 180196 77590
rect 180338 77344 180394 77353
rect 180338 77279 180394 77288
rect 180248 73704 180300 73710
rect 180248 73646 180300 73652
rect 180260 16574 180288 73646
rect 180352 68882 180380 77279
rect 180720 76362 180748 77794
rect 181350 77208 181406 77217
rect 181350 77143 181406 77152
rect 180708 76356 180760 76362
rect 180708 76298 180760 76304
rect 180340 68876 180392 68882
rect 180340 68818 180392 68824
rect 180720 27062 180748 76298
rect 181364 75954 181392 77143
rect 181444 76696 181496 76702
rect 181444 76638 181496 76644
rect 181352 75948 181404 75954
rect 181352 75890 181404 75896
rect 180800 75744 180852 75750
rect 180800 75686 180852 75692
rect 180708 27056 180760 27062
rect 180708 26998 180760 27004
rect 180812 16574 180840 75686
rect 180260 16546 180380 16574
rect 180812 16546 181024 16574
rect 180156 4956 180208 4962
rect 180156 4898 180208 4904
rect 180352 3602 180380 16546
rect 180064 3596 180116 3602
rect 180064 3538 180116 3544
rect 180340 3596 180392 3602
rect 180340 3538 180392 3544
rect 179984 3454 180288 3482
rect 180260 480 180288 3454
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 3942 181484 76638
rect 181534 71768 181590 71777
rect 181534 71703 181590 71712
rect 181444 3936 181496 3942
rect 181444 3878 181496 3884
rect 181548 3534 181576 71703
rect 181640 25770 181668 77862
rect 182192 71738 182220 79426
rect 182916 78464 182968 78470
rect 182916 78406 182968 78412
rect 182180 71732 182232 71738
rect 182180 71674 182232 71680
rect 182086 71496 182142 71505
rect 182086 71431 182142 71440
rect 182100 71097 182128 71431
rect 182086 71088 182142 71097
rect 182086 71023 182142 71032
rect 181628 25764 181680 25770
rect 181628 25706 181680 25712
rect 181536 3528 181588 3534
rect 181536 3470 181588 3476
rect 182100 3398 182128 71023
rect 182824 69692 182876 69698
rect 182824 69634 182876 69640
rect 182180 68876 182232 68882
rect 182180 68818 182232 68824
rect 182088 3392 182140 3398
rect 182088 3334 182140 3340
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 68818
rect 182836 2990 182864 69634
rect 182928 19990 182956 78406
rect 185032 75676 185084 75682
rect 185032 75618 185084 75624
rect 184204 71052 184256 71058
rect 184204 70994 184256 71000
rect 183560 65544 183612 65550
rect 183560 65486 183612 65492
rect 182916 19984 182968 19990
rect 182916 19926 182968 19932
rect 183572 16574 183600 65486
rect 183572 16546 183784 16574
rect 182824 2984 182876 2990
rect 182824 2926 182876 2932
rect 183756 480 183784 16546
rect 184216 4010 184244 70994
rect 185044 6914 185072 75618
rect 186608 64841 186636 199514
rect 186688 197804 186740 197810
rect 186688 197746 186740 197752
rect 186700 76566 186728 197746
rect 186792 80850 186820 200126
rect 186964 148708 187016 148714
rect 186964 148650 187016 148656
rect 186872 139392 186924 139398
rect 186872 139334 186924 139340
rect 186884 139233 186912 139334
rect 186870 139224 186926 139233
rect 186870 139159 186926 139168
rect 186870 139088 186926 139097
rect 186870 139023 186926 139032
rect 186780 80844 186832 80850
rect 186780 80786 186832 80792
rect 186688 76560 186740 76566
rect 186688 76502 186740 76508
rect 186594 64832 186650 64841
rect 186594 64767 186650 64776
rect 186608 64433 186636 64767
rect 186594 64424 186650 64433
rect 186594 64359 186650 64368
rect 186884 60625 186912 139023
rect 186976 71194 187004 148650
rect 187160 145625 187188 273226
rect 193588 265532 193640 265538
rect 193588 265474 193640 265480
rect 192024 265396 192076 265402
rect 192024 265338 192076 265344
rect 190828 263764 190880 263770
rect 190828 263706 190880 263712
rect 187884 263628 187936 263634
rect 187884 263570 187936 263576
rect 187700 262268 187752 262274
rect 187700 262210 187752 262216
rect 187332 259684 187384 259690
rect 187332 259626 187384 259632
rect 187240 259616 187292 259622
rect 187240 259558 187292 259564
rect 187146 145616 187202 145625
rect 187146 145551 187202 145560
rect 187056 143472 187108 143478
rect 187056 143414 187108 143420
rect 187068 73030 187096 143414
rect 187252 141982 187280 259558
rect 187240 141976 187292 141982
rect 187240 141918 187292 141924
rect 187344 141778 187372 259626
rect 187422 213888 187478 213897
rect 187422 213823 187478 213832
rect 187436 143478 187464 213823
rect 187516 200048 187568 200054
rect 187516 199990 187568 199996
rect 187528 199102 187556 199990
rect 187516 199096 187568 199102
rect 187516 199038 187568 199044
rect 187712 198966 187740 262210
rect 187700 198960 187752 198966
rect 187700 198902 187752 198908
rect 187700 197872 187752 197878
rect 187700 197814 187752 197820
rect 187424 143472 187476 143478
rect 187424 143414 187476 143420
rect 187332 141772 187384 141778
rect 187332 141714 187384 141720
rect 187240 140140 187292 140146
rect 187240 140082 187292 140088
rect 187148 139460 187200 139466
rect 187148 139402 187200 139408
rect 187056 73024 187108 73030
rect 187056 72966 187108 72972
rect 187160 71330 187188 139402
rect 187252 72350 187280 140082
rect 187332 140072 187384 140078
rect 187332 140014 187384 140020
rect 187344 76430 187372 140014
rect 187424 139528 187476 139534
rect 187424 139470 187476 139476
rect 187436 139097 187464 139470
rect 187422 139088 187478 139097
rect 187422 139023 187478 139032
rect 187424 80912 187476 80918
rect 187424 80854 187476 80860
rect 187436 80510 187464 80854
rect 187424 80504 187476 80510
rect 187424 80446 187476 80452
rect 187712 76634 187740 197814
rect 187792 196784 187844 196790
rect 187792 196726 187844 196732
rect 187700 76628 187752 76634
rect 187700 76570 187752 76576
rect 187332 76424 187384 76430
rect 187332 76366 187384 76372
rect 187608 73024 187660 73030
rect 187608 72966 187660 72972
rect 187620 72826 187648 72966
rect 187608 72820 187660 72826
rect 187608 72762 187660 72768
rect 187240 72344 187292 72350
rect 187240 72286 187292 72292
rect 187606 71768 187662 71777
rect 187606 71703 187662 71712
rect 187148 71324 187200 71330
rect 187148 71266 187200 71272
rect 186964 71188 187016 71194
rect 186964 71130 187016 71136
rect 187620 70514 187648 71703
rect 187608 70508 187660 70514
rect 187608 70450 187660 70456
rect 187700 64184 187752 64190
rect 187700 64126 187752 64132
rect 186870 60616 186926 60625
rect 186870 60551 186926 60560
rect 186320 60036 186372 60042
rect 186320 59978 186372 59984
rect 186332 16574 186360 59978
rect 187712 16574 187740 64126
rect 187804 61849 187832 196726
rect 187896 143614 187924 263570
rect 188528 263492 188580 263498
rect 188528 263434 188580 263440
rect 188540 262682 188568 263434
rect 189632 262880 189684 262886
rect 189632 262822 189684 262828
rect 187976 262676 188028 262682
rect 187976 262618 188028 262624
rect 188528 262676 188580 262682
rect 188528 262618 188580 262624
rect 187988 262313 188016 262618
rect 187974 262304 188030 262313
rect 187974 262239 188030 262248
rect 188344 261452 188396 261458
rect 188344 261394 188396 261400
rect 188068 260568 188120 260574
rect 188068 260510 188120 260516
rect 187976 260024 188028 260030
rect 187976 259966 188028 259972
rect 187884 143608 187936 143614
rect 187884 143550 187936 143556
rect 187884 143472 187936 143478
rect 187988 143449 188016 259966
rect 188080 143834 188108 260510
rect 188252 259820 188304 259826
rect 188252 259762 188304 259768
rect 188160 195152 188212 195158
rect 188160 195094 188212 195100
rect 188172 143954 188200 195094
rect 188264 146266 188292 259762
rect 188356 193186 188384 261394
rect 189356 260228 189408 260234
rect 189356 260170 189408 260176
rect 189080 197736 189132 197742
rect 189080 197678 189132 197684
rect 188712 193588 188764 193594
rect 188712 193530 188764 193536
rect 188344 193180 188396 193186
rect 188344 193122 188396 193128
rect 188620 178084 188672 178090
rect 188620 178026 188672 178032
rect 188526 146296 188582 146305
rect 188252 146260 188304 146266
rect 188526 146231 188582 146240
rect 188252 146202 188304 146208
rect 188344 146056 188396 146062
rect 188344 145998 188396 146004
rect 188160 143948 188212 143954
rect 188160 143890 188212 143896
rect 188080 143806 188292 143834
rect 188160 143676 188212 143682
rect 188160 143618 188212 143624
rect 188068 143608 188120 143614
rect 188068 143550 188120 143556
rect 187884 143414 187936 143420
rect 187974 143440 188030 143449
rect 187896 142186 187924 143414
rect 187974 143375 188030 143384
rect 188080 143041 188108 143550
rect 188066 143032 188122 143041
rect 188066 142967 188122 142976
rect 187884 142180 187936 142186
rect 187884 142122 187936 142128
rect 187790 61840 187846 61849
rect 187790 61775 187846 61784
rect 187790 59120 187846 59129
rect 187790 59055 187846 59064
rect 187804 58857 187832 59055
rect 187790 58848 187846 58857
rect 187790 58783 187846 58792
rect 187896 20670 187924 142122
rect 187976 141092 188028 141098
rect 187976 141034 188028 141040
rect 187988 139398 188016 141034
rect 188068 140004 188120 140010
rect 188068 139946 188120 139952
rect 187976 139392 188028 139398
rect 187976 139334 188028 139340
rect 187976 139256 188028 139262
rect 187976 139198 188028 139204
rect 187988 50697 188016 139198
rect 188080 52193 188108 139946
rect 188172 80782 188200 143618
rect 188264 142866 188292 143806
rect 188252 142860 188304 142866
rect 188252 142802 188304 142808
rect 188252 140616 188304 140622
rect 188252 140558 188304 140564
rect 188264 139466 188292 140558
rect 188252 139460 188304 139466
rect 188252 139402 188304 139408
rect 188250 139360 188306 139369
rect 188250 139295 188306 139304
rect 188160 80776 188212 80782
rect 188160 80718 188212 80724
rect 188264 64874 188292 139295
rect 188356 71262 188384 145998
rect 188436 143268 188488 143274
rect 188436 143210 188488 143216
rect 188448 142662 188476 143210
rect 188436 142656 188488 142662
rect 188436 142598 188488 142604
rect 188436 140956 188488 140962
rect 188436 140898 188488 140904
rect 188344 71256 188396 71262
rect 188344 71198 188396 71204
rect 188448 69630 188476 140898
rect 188540 75313 188568 146231
rect 188632 144294 188660 178026
rect 188620 144288 188672 144294
rect 188620 144230 188672 144236
rect 188620 140548 188672 140554
rect 188620 140490 188672 140496
rect 188632 139942 188660 140490
rect 188620 139936 188672 139942
rect 188620 139878 188672 139884
rect 188724 139777 188752 193530
rect 188710 139768 188766 139777
rect 188710 139703 188766 139712
rect 188620 80912 188672 80918
rect 188620 80854 188672 80860
rect 188632 80714 188660 80854
rect 188620 80708 188672 80714
rect 188620 80650 188672 80656
rect 188988 76968 189040 76974
rect 188988 76910 189040 76916
rect 188526 75304 188582 75313
rect 188526 75239 188582 75248
rect 188436 69624 188488 69630
rect 188436 69566 188488 69572
rect 189000 67634 189028 76910
rect 189092 72434 189120 197678
rect 189172 195220 189224 195226
rect 189172 195162 189224 195168
rect 189184 76974 189212 195162
rect 189262 194984 189318 194993
rect 189262 194919 189318 194928
rect 189276 80714 189304 194919
rect 189368 141642 189396 260170
rect 189540 260160 189592 260166
rect 189540 260102 189592 260108
rect 189448 260092 189500 260098
rect 189448 260034 189500 260040
rect 189460 142730 189488 260034
rect 189552 143342 189580 260102
rect 189644 145586 189672 262822
rect 190460 262336 190512 262342
rect 190460 262278 190512 262284
rect 189724 260976 189776 260982
rect 189724 260918 189776 260924
rect 189632 145580 189684 145586
rect 189632 145522 189684 145528
rect 189736 145382 189764 260918
rect 190366 199880 190422 199889
rect 190366 199815 190422 199824
rect 190380 192681 190408 199815
rect 190472 199442 190500 262278
rect 190552 259752 190604 259758
rect 190552 259694 190604 259700
rect 190564 200190 190592 259694
rect 190552 200184 190604 200190
rect 190552 200126 190604 200132
rect 190460 199436 190512 199442
rect 190460 199378 190512 199384
rect 190644 195968 190696 195974
rect 190644 195910 190696 195916
rect 190460 195560 190512 195566
rect 190460 195502 190512 195508
rect 190366 192672 190422 192681
rect 190366 192607 190422 192616
rect 189816 165640 189868 165646
rect 189816 165582 189868 165588
rect 189724 145376 189776 145382
rect 189724 145318 189776 145324
rect 189828 144226 189856 165582
rect 190092 145920 190144 145926
rect 190092 145862 190144 145868
rect 190000 145444 190052 145450
rect 190000 145386 190052 145392
rect 189816 144220 189868 144226
rect 189816 144162 189868 144168
rect 189540 143336 189592 143342
rect 189540 143278 189592 143284
rect 189448 142724 189500 142730
rect 189448 142666 189500 142672
rect 189356 141636 189408 141642
rect 189356 141578 189408 141584
rect 189540 141500 189592 141506
rect 189540 141442 189592 141448
rect 189356 140276 189408 140282
rect 189356 140218 189408 140224
rect 189264 80708 189316 80714
rect 189264 80650 189316 80656
rect 189172 76968 189224 76974
rect 189172 76910 189224 76916
rect 189092 72406 189304 72434
rect 189000 67606 189212 67634
rect 189078 67552 189134 67561
rect 189078 67487 189134 67496
rect 189092 67017 189120 67487
rect 189078 67008 189134 67017
rect 189078 66943 189134 66952
rect 188264 64846 188384 64874
rect 188356 58857 188384 64846
rect 189184 63209 189212 67606
rect 189276 67590 189304 72406
rect 189264 67584 189316 67590
rect 189264 67526 189316 67532
rect 189276 66978 189304 67526
rect 189264 66972 189316 66978
rect 189264 66914 189316 66920
rect 189170 63200 189226 63209
rect 189170 63135 189226 63144
rect 188342 58848 188398 58857
rect 188342 58783 188398 58792
rect 189368 53553 189396 140218
rect 189552 67561 189580 141442
rect 189908 140344 189960 140350
rect 189908 140286 189960 140292
rect 189816 140208 189868 140214
rect 189816 140150 189868 140156
rect 189828 72894 189856 140150
rect 189920 75138 189948 140286
rect 189908 75132 189960 75138
rect 189908 75074 189960 75080
rect 189816 72888 189868 72894
rect 189816 72830 189868 72836
rect 189538 67552 189594 67561
rect 189538 67487 189594 67496
rect 190012 60217 190040 145386
rect 190104 72418 190132 145862
rect 190184 145512 190236 145518
rect 190184 145454 190236 145460
rect 190196 73914 190224 145454
rect 190184 73908 190236 73914
rect 190184 73850 190236 73856
rect 190092 72412 190144 72418
rect 190092 72354 190144 72360
rect 190366 71768 190422 71777
rect 190366 71703 190422 71712
rect 190380 70446 190408 71703
rect 190368 70440 190420 70446
rect 190368 70382 190420 70388
rect 189998 60208 190054 60217
rect 189998 60143 190054 60152
rect 189354 53544 189410 53553
rect 189354 53479 189410 53488
rect 188066 52184 188122 52193
rect 188066 52119 188122 52128
rect 187974 50688 188030 50697
rect 187974 50623 188030 50632
rect 190472 45393 190500 195502
rect 190552 195424 190604 195430
rect 190552 195366 190604 195372
rect 190564 53825 190592 195366
rect 190656 57905 190684 195910
rect 190736 195900 190788 195906
rect 190736 195842 190788 195848
rect 190748 61713 190776 195842
rect 190840 141710 190868 263706
rect 190920 263696 190972 263702
rect 190920 263638 190972 263644
rect 190932 144770 190960 263638
rect 191012 262608 191064 262614
rect 191012 262550 191064 262556
rect 190920 144764 190972 144770
rect 190920 144706 190972 144712
rect 191024 144362 191052 262550
rect 191288 261248 191340 261254
rect 191288 261190 191340 261196
rect 191104 260432 191156 260438
rect 191104 260374 191156 260380
rect 191012 144356 191064 144362
rect 191012 144298 191064 144304
rect 191116 143070 191144 260374
rect 191196 259888 191248 259894
rect 191196 259830 191248 259836
rect 191104 143064 191156 143070
rect 191104 143006 191156 143012
rect 191208 142934 191236 259830
rect 191300 146198 191328 261190
rect 191840 195764 191892 195770
rect 191840 195706 191892 195712
rect 191288 146192 191340 146198
rect 191288 146134 191340 146140
rect 191380 145716 191432 145722
rect 191380 145658 191432 145664
rect 191196 142928 191248 142934
rect 191196 142870 191248 142876
rect 190920 142792 190972 142798
rect 190920 142734 190972 142740
rect 190828 141704 190880 141710
rect 190828 141646 190880 141652
rect 190828 140480 190880 140486
rect 190828 140422 190880 140428
rect 190734 61704 190790 61713
rect 190734 61639 190790 61648
rect 190642 57896 190698 57905
rect 190642 57831 190698 57840
rect 190550 53816 190606 53825
rect 190550 53751 190606 53760
rect 190840 53145 190868 140422
rect 190932 80054 190960 142734
rect 191286 140312 191342 140321
rect 191286 140247 191342 140256
rect 191102 139360 191158 139369
rect 191102 139295 191158 139304
rect 190932 80026 191052 80054
rect 191024 73098 191052 80026
rect 191116 77042 191144 139295
rect 191194 138680 191250 138689
rect 191194 138615 191250 138624
rect 191208 79150 191236 138615
rect 191300 81161 191328 140247
rect 191286 81152 191342 81161
rect 191286 81087 191342 81096
rect 191196 79144 191248 79150
rect 191196 79086 191248 79092
rect 191392 78878 191420 145658
rect 191380 78872 191432 78878
rect 191380 78814 191432 78820
rect 191104 77036 191156 77042
rect 191104 76978 191156 76984
rect 191012 73092 191064 73098
rect 191012 73034 191064 73040
rect 191024 72894 191052 73034
rect 191012 72888 191064 72894
rect 191012 72830 191064 72836
rect 191852 58721 191880 195706
rect 191932 195356 191984 195362
rect 191932 195298 191984 195304
rect 191944 60489 191972 195298
rect 192036 144702 192064 265338
rect 193128 263424 193180 263430
rect 193128 263366 193180 263372
rect 192392 262812 192444 262818
rect 192392 262754 192444 262760
rect 192208 262744 192260 262750
rect 192208 262686 192260 262692
rect 192116 262472 192168 262478
rect 192116 262414 192168 262420
rect 192024 144696 192076 144702
rect 192024 144638 192076 144644
rect 192128 141914 192156 262414
rect 192116 141908 192168 141914
rect 192116 141850 192168 141856
rect 192220 141574 192248 262686
rect 192300 262540 192352 262546
rect 192300 262482 192352 262488
rect 192312 262313 192340 262482
rect 192298 262304 192354 262313
rect 192298 262239 192354 262248
rect 192300 260500 192352 260506
rect 192300 260442 192352 260448
rect 192312 142118 192340 260442
rect 192404 144566 192432 262754
rect 193140 262546 193168 263366
rect 193128 262540 193180 262546
rect 193128 262482 193180 262488
rect 193312 200320 193364 200326
rect 193312 200262 193364 200268
rect 193220 197260 193272 197266
rect 193220 197202 193272 197208
rect 192576 195832 192628 195838
rect 192576 195774 192628 195780
rect 192484 193044 192536 193050
rect 192484 192986 192536 192992
rect 192392 144560 192444 144566
rect 192392 144502 192444 144508
rect 192300 142112 192352 142118
rect 192300 142054 192352 142060
rect 192208 141568 192260 141574
rect 192208 141510 192260 141516
rect 192024 140752 192076 140758
rect 192024 140694 192076 140700
rect 192036 66230 192064 140694
rect 192300 139936 192352 139942
rect 192300 139878 192352 139884
rect 192114 76936 192170 76945
rect 192114 76871 192170 76880
rect 192128 76537 192156 76871
rect 192114 76528 192170 76537
rect 192114 76463 192170 76472
rect 192116 71732 192168 71738
rect 192116 71674 192168 71680
rect 192128 71058 192156 71674
rect 192312 71466 192340 139878
rect 192496 75070 192524 192986
rect 192588 78266 192616 195774
rect 193126 146160 193182 146169
rect 193126 146095 193182 146104
rect 192944 145648 192996 145654
rect 193140 145625 193168 146095
rect 192944 145590 192996 145596
rect 193126 145616 193182 145625
rect 192760 144900 192812 144906
rect 192760 144842 192812 144848
rect 192666 138000 192722 138009
rect 192666 137935 192722 137944
rect 192576 78260 192628 78266
rect 192576 78202 192628 78208
rect 192588 77722 192616 78202
rect 192576 77716 192628 77722
rect 192576 77658 192628 77664
rect 192680 77294 192708 137935
rect 192588 77266 192708 77294
rect 192484 75064 192536 75070
rect 192484 75006 192536 75012
rect 192300 71460 192352 71466
rect 192300 71402 192352 71408
rect 192116 71052 192168 71058
rect 192116 70994 192168 71000
rect 192588 70106 192616 77266
rect 192576 70100 192628 70106
rect 192576 70042 192628 70048
rect 192772 70038 192800 144842
rect 192852 144492 192904 144498
rect 192852 144434 192904 144440
rect 192864 71058 192892 144434
rect 192956 76537 192984 145590
rect 193126 145551 193182 145560
rect 192942 76528 192998 76537
rect 192942 76463 192998 76472
rect 192852 71052 192904 71058
rect 192852 70994 192904 71000
rect 192760 70032 192812 70038
rect 192760 69974 192812 69980
rect 192772 69698 192800 69974
rect 192760 69692 192812 69698
rect 192760 69634 192812 69640
rect 192482 68232 192538 68241
rect 192482 68167 192538 68176
rect 192024 66224 192076 66230
rect 192024 66166 192076 66172
rect 191930 60480 191986 60489
rect 191930 60415 191986 60424
rect 191838 58712 191894 58721
rect 191838 58647 191894 58656
rect 190826 53136 190882 53145
rect 190826 53071 190882 53080
rect 190458 45384 190514 45393
rect 190458 45319 190514 45328
rect 191840 36916 191892 36922
rect 191840 36858 191892 36864
rect 187884 20664 187936 20670
rect 187884 20606 187936 20612
rect 191852 16574 191880 36858
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 191852 16546 192064 16574
rect 184952 6886 185072 6914
rect 184204 4004 184256 4010
rect 184204 3946 184256 3952
rect 184952 480 184980 6886
rect 186136 3528 186188 3534
rect 186136 3470 186188 3476
rect 186148 480 186176 3470
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 190828 3936 190880 3942
rect 190828 3878 190880 3884
rect 189724 2984 189776 2990
rect 189724 2926 189776 2932
rect 189736 480 189764 2926
rect 190840 480 190868 3878
rect 192036 480 192064 16546
rect 192496 3262 192524 68167
rect 193128 66224 193180 66230
rect 193128 66166 193180 66172
rect 193140 65550 193168 66166
rect 193128 65544 193180 65550
rect 193128 65486 193180 65492
rect 193126 60480 193182 60489
rect 193126 60415 193182 60424
rect 193140 60081 193168 60415
rect 193126 60072 193182 60081
rect 193126 60007 193182 60016
rect 193232 48113 193260 197202
rect 193324 57866 193352 200262
rect 193496 200252 193548 200258
rect 193496 200194 193548 200200
rect 193404 196648 193456 196654
rect 193404 196590 193456 196596
rect 193312 57860 193364 57866
rect 193312 57802 193364 57808
rect 193416 56506 193444 196590
rect 193508 63510 193536 200194
rect 193600 144838 193628 265474
rect 193772 265464 193824 265470
rect 193772 265406 193824 265412
rect 193680 262404 193732 262410
rect 193680 262346 193732 262352
rect 193588 144832 193640 144838
rect 193588 144774 193640 144780
rect 193692 143478 193720 262346
rect 193784 146742 193812 265406
rect 197820 265328 197872 265334
rect 197820 265270 197872 265276
rect 194968 265260 195020 265266
rect 194968 265202 195020 265208
rect 194048 198620 194100 198626
rect 194048 198562 194100 198568
rect 193864 197940 193916 197946
rect 193864 197882 193916 197888
rect 193772 146736 193824 146742
rect 193772 146678 193824 146684
rect 193876 146305 193904 197882
rect 193956 147280 194008 147286
rect 193956 147222 194008 147228
rect 193862 146296 193918 146305
rect 193862 146231 193918 146240
rect 193680 143472 193732 143478
rect 193680 143414 193732 143420
rect 193864 140412 193916 140418
rect 193864 140354 193916 140360
rect 193588 77104 193640 77110
rect 193588 77046 193640 77052
rect 193600 76702 193628 77046
rect 193588 76696 193640 76702
rect 193588 76638 193640 76644
rect 193876 74390 193904 140354
rect 193968 80889 193996 147222
rect 194060 146169 194088 198562
rect 194692 197056 194744 197062
rect 194692 196998 194744 197004
rect 194600 195628 194652 195634
rect 194600 195570 194652 195576
rect 194324 147484 194376 147490
rect 194324 147426 194376 147432
rect 194046 146160 194102 146169
rect 194046 146095 194102 146104
rect 194140 145988 194192 145994
rect 194140 145930 194192 145936
rect 194048 140004 194100 140010
rect 194048 139946 194100 139952
rect 193954 80880 194010 80889
rect 193954 80815 194010 80824
rect 194060 76702 194088 139946
rect 194048 76696 194100 76702
rect 194048 76638 194100 76644
rect 193864 74384 193916 74390
rect 193864 74326 193916 74332
rect 194152 70174 194180 145930
rect 194232 145852 194284 145858
rect 194232 145794 194284 145800
rect 194140 70168 194192 70174
rect 194140 70110 194192 70116
rect 193862 67280 193918 67289
rect 193862 67215 193918 67224
rect 193496 63504 193548 63510
rect 193496 63446 193548 63452
rect 193508 62830 193536 63446
rect 193496 62824 193548 62830
rect 193496 62766 193548 62772
rect 193404 56500 193456 56506
rect 193404 56442 193456 56448
rect 193310 55856 193366 55865
rect 193310 55791 193366 55800
rect 193218 48104 193274 48113
rect 193218 48039 193274 48048
rect 193324 16574 193352 55791
rect 193324 16546 193812 16574
rect 193784 3482 193812 16546
rect 193876 3942 193904 67215
rect 194046 66192 194102 66201
rect 194046 66127 194048 66136
rect 194100 66127 194102 66136
rect 194048 66098 194100 66104
rect 194244 60654 194272 145794
rect 194336 79422 194364 147426
rect 194324 79416 194376 79422
rect 194324 79358 194376 79364
rect 194508 66156 194560 66162
rect 194508 66098 194560 66104
rect 194520 64938 194548 66098
rect 194508 64932 194560 64938
rect 194508 64874 194560 64880
rect 194232 60648 194284 60654
rect 194232 60590 194284 60596
rect 194508 60648 194560 60654
rect 194508 60590 194560 60596
rect 194520 60042 194548 60590
rect 194508 60036 194560 60042
rect 194508 59978 194560 59984
rect 194508 57860 194560 57866
rect 194508 57802 194560 57808
rect 194520 57322 194548 57802
rect 194508 57316 194560 57322
rect 194508 57258 194560 57264
rect 194508 56500 194560 56506
rect 194508 56442 194560 56448
rect 194520 55962 194548 56442
rect 194508 55956 194560 55962
rect 194508 55898 194560 55904
rect 194612 52329 194640 195570
rect 194704 55185 194732 196998
rect 194876 196920 194928 196926
rect 194876 196862 194928 196868
rect 194784 195288 194836 195294
rect 194784 195230 194836 195236
rect 194796 59265 194824 195230
rect 194888 64870 194916 196862
rect 194980 144634 195008 265202
rect 195152 265192 195204 265198
rect 195152 265134 195204 265140
rect 195060 264988 195112 264994
rect 195060 264930 195112 264936
rect 195072 146033 195100 264930
rect 195164 146810 195192 265134
rect 196256 265124 196308 265130
rect 196256 265066 196308 265072
rect 195244 259548 195296 259554
rect 195244 259490 195296 259496
rect 195152 146804 195204 146810
rect 195152 146746 195204 146752
rect 195058 146024 195114 146033
rect 195058 145959 195114 145968
rect 195152 145784 195204 145790
rect 195152 145726 195204 145732
rect 194968 144628 195020 144634
rect 194968 144570 195020 144576
rect 195060 143404 195112 143410
rect 195060 143346 195112 143352
rect 195072 69578 195100 143346
rect 195164 80054 195192 145726
rect 195256 143342 195284 259490
rect 195520 199844 195572 199850
rect 195520 199786 195572 199792
rect 195532 179353 195560 199786
rect 195980 198688 196032 198694
rect 195978 198656 195980 198665
rect 196032 198656 196034 198665
rect 195978 198591 196034 198600
rect 196072 195696 196124 195702
rect 196072 195638 196124 195644
rect 195980 192772 196032 192778
rect 195980 192714 196032 192720
rect 195518 179344 195574 179353
rect 195518 179279 195574 179288
rect 195520 148776 195572 148782
rect 195520 148718 195572 148724
rect 195336 147416 195388 147422
rect 195336 147358 195388 147364
rect 195244 143336 195296 143342
rect 195244 143278 195296 143284
rect 195164 80026 195284 80054
rect 195072 69550 195192 69578
rect 195164 67522 195192 69550
rect 195256 68950 195284 80026
rect 195348 76673 195376 147358
rect 195428 147212 195480 147218
rect 195428 147154 195480 147160
rect 195440 78946 195468 147154
rect 195428 78940 195480 78946
rect 195428 78882 195480 78888
rect 195334 76664 195390 76673
rect 195334 76599 195390 76608
rect 195532 72214 195560 148718
rect 195520 72208 195572 72214
rect 195520 72150 195572 72156
rect 195244 68944 195296 68950
rect 195244 68886 195296 68892
rect 195256 68474 195284 68886
rect 195244 68468 195296 68474
rect 195244 68410 195296 68416
rect 195152 67516 195204 67522
rect 195152 67458 195204 67464
rect 195164 66910 195192 67458
rect 195152 66904 195204 66910
rect 195152 66846 195204 66852
rect 194876 64864 194928 64870
rect 194876 64806 194928 64812
rect 194888 64258 194916 64806
rect 194876 64252 194928 64258
rect 194876 64194 194928 64200
rect 194782 59256 194838 59265
rect 194782 59191 194838 59200
rect 195058 59256 195114 59265
rect 195058 59191 195114 59200
rect 195072 58585 195100 59191
rect 195058 58576 195114 58585
rect 195058 58511 195114 58520
rect 194690 55176 194746 55185
rect 194690 55111 194746 55120
rect 194598 52320 194654 52329
rect 194598 52255 194654 52264
rect 194612 52057 194640 52255
rect 194598 52048 194654 52057
rect 194598 51983 194654 51992
rect 195992 50833 196020 192714
rect 196084 53689 196112 195638
rect 196164 195492 196216 195498
rect 196164 195434 196216 195440
rect 196176 56545 196204 195434
rect 196268 139874 196296 265066
rect 196716 261180 196768 261186
rect 196716 261122 196768 261128
rect 196532 261112 196584 261118
rect 196532 261054 196584 261060
rect 196440 261044 196492 261050
rect 196440 260986 196492 260992
rect 196348 196852 196400 196858
rect 196348 196794 196400 196800
rect 196256 139868 196308 139874
rect 196256 139810 196308 139816
rect 196256 78940 196308 78946
rect 196256 78882 196308 78888
rect 196268 78538 196296 78882
rect 196256 78532 196308 78538
rect 196256 78474 196308 78480
rect 196360 75818 196388 196794
rect 196452 143206 196480 260986
rect 196544 147626 196572 261054
rect 196624 198348 196676 198354
rect 196624 198290 196676 198296
rect 196532 147620 196584 147626
rect 196532 147562 196584 147568
rect 196532 147348 196584 147354
rect 196532 147290 196584 147296
rect 196440 143200 196492 143206
rect 196440 143142 196492 143148
rect 196440 141840 196492 141846
rect 196440 141782 196492 141788
rect 196348 75812 196400 75818
rect 196348 75754 196400 75760
rect 196452 71398 196480 141782
rect 196544 78742 196572 147290
rect 196636 78946 196664 198290
rect 196728 148374 196756 261122
rect 197360 200524 197412 200530
rect 197360 200466 197412 200472
rect 196992 148504 197044 148510
rect 196992 148446 197044 148452
rect 196716 148368 196768 148374
rect 196716 148310 196768 148316
rect 196716 147076 196768 147082
rect 196716 147018 196768 147024
rect 196624 78940 196676 78946
rect 196624 78882 196676 78888
rect 196728 78810 196756 147018
rect 196806 139088 196862 139097
rect 196806 139023 196862 139032
rect 196820 93854 196848 139023
rect 196820 93826 196940 93854
rect 196806 80064 196862 80073
rect 196806 79999 196862 80008
rect 196820 79354 196848 79999
rect 196808 79348 196860 79354
rect 196808 79290 196860 79296
rect 196820 78810 196848 79290
rect 196716 78804 196768 78810
rect 196716 78746 196768 78752
rect 196808 78804 196860 78810
rect 196808 78746 196860 78752
rect 196532 78736 196584 78742
rect 196532 78678 196584 78684
rect 196912 78554 196940 93826
rect 196728 78526 196940 78554
rect 196728 77246 196756 78526
rect 196716 77240 196768 77246
rect 196716 77182 196768 77188
rect 196728 76634 196756 77182
rect 196716 76628 196768 76634
rect 196716 76570 196768 76576
rect 197004 71534 197032 148446
rect 196992 71528 197044 71534
rect 196992 71470 197044 71476
rect 196440 71392 196492 71398
rect 196440 71334 196492 71340
rect 196624 69828 196676 69834
rect 196624 69770 196676 69776
rect 196254 68912 196310 68921
rect 196254 68847 196256 68856
rect 196308 68847 196310 68856
rect 196256 68818 196308 68824
rect 196268 67658 196296 68818
rect 196256 67652 196308 67658
rect 196256 67594 196308 67600
rect 196162 56536 196218 56545
rect 196162 56471 196218 56480
rect 196176 56001 196204 56471
rect 196162 55992 196218 56001
rect 196162 55927 196218 55936
rect 196070 53680 196126 53689
rect 196070 53615 196126 53624
rect 196084 53281 196112 53615
rect 196070 53272 196126 53281
rect 196070 53207 196126 53216
rect 195978 50824 196034 50833
rect 195978 50759 196034 50768
rect 196438 50824 196494 50833
rect 196438 50759 196494 50768
rect 196452 50561 196480 50759
rect 196438 50552 196494 50561
rect 196438 50487 196494 50496
rect 194506 48104 194562 48113
rect 194506 48039 194562 48048
rect 194520 47841 194548 48039
rect 194506 47832 194562 47841
rect 194506 47767 194562 47776
rect 194600 32700 194652 32706
rect 194600 32642 194652 32648
rect 194612 16574 194640 32642
rect 196636 16574 196664 69770
rect 197372 49473 197400 200466
rect 197728 198416 197780 198422
rect 197728 198358 197780 198364
rect 197452 197124 197504 197130
rect 197452 197066 197504 197072
rect 197464 62218 197492 197066
rect 197544 196988 197596 196994
rect 197544 196930 197596 196936
rect 197452 62212 197504 62218
rect 197452 62154 197504 62160
rect 197452 62076 197504 62082
rect 197452 62018 197504 62024
rect 197464 61470 197492 62018
rect 197452 61464 197504 61470
rect 197452 61406 197504 61412
rect 197452 60716 197504 60722
rect 197452 60658 197504 60664
rect 197464 60110 197492 60658
rect 197452 60104 197504 60110
rect 197452 60046 197504 60052
rect 197452 57248 197504 57254
rect 197452 57190 197504 57196
rect 197358 49464 197414 49473
rect 197358 49399 197414 49408
rect 197464 16574 197492 57190
rect 197556 52465 197584 196930
rect 197636 196716 197688 196722
rect 197636 196658 197688 196664
rect 197648 62082 197676 196658
rect 197740 64705 197768 198358
rect 197832 146130 197860 265270
rect 197912 265056 197964 265062
rect 197912 264998 197964 265004
rect 197924 146878 197952 264998
rect 218072 263430 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 278089 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700670 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 234618 278080 234674 278089
rect 234618 278015 234674 278024
rect 218060 263424 218112 263430
rect 218060 263366 218112 263372
rect 282932 262886 282960 702406
rect 299492 276729 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700466 332548 703520
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 299478 276720 299534 276729
rect 299478 276655 299534 276664
rect 347792 263498 347820 702406
rect 364352 273970 364380 702406
rect 397472 699718 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 429856 699718 429884 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 396736 284889 396764 699654
rect 396722 284880 396778 284889
rect 396722 284815 396778 284824
rect 428476 275330 428504 699654
rect 462332 287706 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 287700 462372 287706
rect 462320 287642 462372 287648
rect 428464 275324 428516 275330
rect 428464 275266 428516 275272
rect 364340 273964 364392 273970
rect 364340 273906 364392 273912
rect 347780 263492 347832 263498
rect 347780 263434 347832 263440
rect 282920 262880 282972 262886
rect 477512 262857 477540 702406
rect 489184 700392 489236 700398
rect 489184 700334 489236 700340
rect 489196 283626 489224 700334
rect 489184 283620 489236 283626
rect 489184 283562 489236 283568
rect 494072 271182 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 527824 700392 527876 700398
rect 527824 700334 527876 700340
rect 498844 670744 498896 670750
rect 498844 670686 498896 670692
rect 494060 271176 494112 271182
rect 494060 271118 494112 271124
rect 498856 268394 498884 670686
rect 527836 269822 527864 700334
rect 543476 700330 543504 703520
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 527824 269816 527876 269822
rect 527824 269758 527876 269764
rect 498844 268388 498896 268394
rect 498844 268330 498896 268336
rect 580276 263566 580304 365055
rect 580264 263560 580316 263566
rect 580264 263502 580316 263508
rect 580356 263016 580408 263022
rect 580356 262958 580408 262964
rect 282920 262822 282972 262828
rect 477498 262848 477554 262857
rect 477498 262783 477554 262792
rect 198096 261384 198148 261390
rect 198096 261326 198148 261332
rect 198004 260908 198056 260914
rect 198004 260850 198056 260856
rect 197912 146872 197964 146878
rect 197912 146814 197964 146820
rect 197820 146124 197872 146130
rect 197820 146066 197872 146072
rect 198016 143138 198044 260850
rect 198108 147558 198136 261326
rect 471244 261316 471296 261322
rect 471244 261258 471296 261264
rect 471256 206990 471284 261258
rect 472624 260364 472676 260370
rect 472624 260306 472676 260312
rect 472636 245614 472664 260306
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 472624 245608 472676 245614
rect 580172 245608 580224 245614
rect 472624 245550 472676 245556
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580368 219065 580396 262958
rect 580448 262948 580500 262954
rect 580448 262890 580500 262896
rect 580460 232393 580488 262890
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 471244 206984 471296 206990
rect 471244 206926 471296 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 198832 200456 198884 200462
rect 198832 200398 198884 200404
rect 198740 199096 198792 199102
rect 198740 199038 198792 199044
rect 198188 198280 198240 198286
rect 198188 198222 198240 198228
rect 198200 147801 198228 198222
rect 198280 148572 198332 148578
rect 198280 148514 198332 148520
rect 198186 147792 198242 147801
rect 198186 147727 198242 147736
rect 198096 147552 198148 147558
rect 198096 147494 198148 147500
rect 198096 147008 198148 147014
rect 198096 146950 198148 146956
rect 198004 143132 198056 143138
rect 198004 143074 198056 143080
rect 198004 141432 198056 141438
rect 198004 141374 198056 141380
rect 197820 77172 197872 77178
rect 197820 77114 197872 77120
rect 197832 76566 197860 77114
rect 197820 76560 197872 76566
rect 197820 76502 197872 76508
rect 198016 71670 198044 141374
rect 198108 79218 198136 146950
rect 198186 138952 198242 138961
rect 198186 138887 198242 138896
rect 198096 79212 198148 79218
rect 198096 79154 198148 79160
rect 198200 77178 198228 138887
rect 198188 77172 198240 77178
rect 198188 77114 198240 77120
rect 198004 71664 198056 71670
rect 198004 71606 198056 71612
rect 198292 70242 198320 148514
rect 198372 147144 198424 147150
rect 198372 147086 198424 147092
rect 198384 75002 198412 147086
rect 198752 146305 198780 199038
rect 198738 146296 198794 146305
rect 198738 146231 198794 146240
rect 198740 78872 198792 78878
rect 198740 78814 198792 78820
rect 198752 78441 198780 78814
rect 198738 78432 198794 78441
rect 198738 78367 198794 78376
rect 198740 75608 198792 75614
rect 198740 75550 198792 75556
rect 198372 74996 198424 75002
rect 198372 74938 198424 74944
rect 198280 70236 198332 70242
rect 198280 70178 198332 70184
rect 197726 64696 197782 64705
rect 197726 64631 197782 64640
rect 197740 64297 197768 64631
rect 197726 64288 197782 64297
rect 197726 64223 197782 64232
rect 197728 62212 197780 62218
rect 197728 62154 197780 62160
rect 197636 62076 197688 62082
rect 197636 62018 197688 62024
rect 197740 60722 197768 62154
rect 197728 60716 197780 60722
rect 197728 60658 197780 60664
rect 197542 52456 197598 52465
rect 197542 52391 197598 52400
rect 198002 52456 198058 52465
rect 198002 52391 198058 52400
rect 198016 51785 198044 52391
rect 198002 51776 198058 51785
rect 198002 51711 198058 51720
rect 198462 49464 198518 49473
rect 198462 49399 198518 49408
rect 198476 49201 198504 49399
rect 198462 49192 198518 49201
rect 198462 49127 198518 49136
rect 194612 16546 195192 16574
rect 196636 16546 196940 16574
rect 197464 16546 197952 16574
rect 193864 3936 193916 3942
rect 193864 3878 193916 3884
rect 193784 3454 194456 3482
rect 192484 3256 192536 3262
rect 192484 3198 192536 3204
rect 193220 3256 193272 3262
rect 193220 3198 193272 3204
rect 193232 480 193260 3198
rect 194428 480 194456 3454
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196912 3942 196940 16546
rect 196808 3936 196860 3942
rect 196808 3878 196860 3884
rect 196900 3936 196952 3942
rect 196900 3878 196952 3884
rect 196820 480 196848 3878
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 75550
rect 198844 55049 198872 200398
rect 201498 200288 201554 200297
rect 201498 200223 201554 200232
rect 199568 199776 199620 199782
rect 199568 199718 199620 199724
rect 199108 198484 199160 198490
rect 199108 198426 199160 198432
rect 199016 197328 199068 197334
rect 199016 197270 199068 197276
rect 198922 196616 198978 196625
rect 198922 196551 198978 196560
rect 198936 57361 198964 196551
rect 199028 63345 199056 197270
rect 199120 79286 199148 198426
rect 199580 198218 199608 199718
rect 201040 199164 201092 199170
rect 201040 199106 201092 199112
rect 200212 199028 200264 199034
rect 200212 198970 200264 198976
rect 199568 198212 199620 198218
rect 199568 198154 199620 198160
rect 199384 198008 199436 198014
rect 199384 197950 199436 197956
rect 199200 152652 199252 152658
rect 199200 152594 199252 152600
rect 199108 79280 199160 79286
rect 199108 79222 199160 79228
rect 199108 78736 199160 78742
rect 199108 78678 199160 78684
rect 199120 77489 199148 78678
rect 199106 77480 199162 77489
rect 199106 77415 199162 77424
rect 199108 69012 199160 69018
rect 199108 68954 199160 68960
rect 199120 68406 199148 68954
rect 199108 68400 199160 68406
rect 199108 68342 199160 68348
rect 199014 63336 199070 63345
rect 199014 63271 199070 63280
rect 199212 62778 199240 152594
rect 199292 152584 199344 152590
rect 199292 152526 199344 152532
rect 199304 71602 199332 152526
rect 199396 78878 199424 197950
rect 199660 197192 199712 197198
rect 199660 197134 199712 197140
rect 199476 148436 199528 148442
rect 199476 148378 199528 148384
rect 199384 78872 199436 78878
rect 199384 78814 199436 78820
rect 199488 73166 199516 148378
rect 199566 145616 199622 145625
rect 199566 145551 199622 145560
rect 199580 78742 199608 145551
rect 199568 78736 199620 78742
rect 199568 78678 199620 78684
rect 199476 73160 199528 73166
rect 199476 73102 199528 73108
rect 199292 71596 199344 71602
rect 199292 71538 199344 71544
rect 199566 70408 199622 70417
rect 199566 70343 199622 70352
rect 199580 69970 199608 70343
rect 199568 69964 199620 69970
rect 199568 69906 199620 69912
rect 199580 69086 199608 69906
rect 199568 69080 199620 69086
rect 199568 69022 199620 69028
rect 199672 69018 199700 197134
rect 200118 138816 200174 138825
rect 200118 138751 200174 138760
rect 200132 71210 200160 138751
rect 200040 71182 200160 71210
rect 200040 70922 200068 71182
rect 200120 71052 200172 71058
rect 200120 70994 200172 71000
rect 200028 70916 200080 70922
rect 200028 70858 200080 70864
rect 199660 69012 199712 69018
rect 199660 68954 199712 68960
rect 199382 63336 199438 63345
rect 199382 63271 199438 63280
rect 199396 63073 199424 63271
rect 199382 63064 199438 63073
rect 199382 62999 199438 63008
rect 199028 62750 199240 62778
rect 199028 62014 199056 62750
rect 199016 62008 199068 62014
rect 199016 61950 199068 61956
rect 199028 61402 199056 61950
rect 199016 61396 199068 61402
rect 199016 61338 199068 61344
rect 198922 57352 198978 57361
rect 198922 57287 198978 57296
rect 198830 55040 198886 55049
rect 198830 54975 198886 54984
rect 198844 54505 198872 54975
rect 198830 54496 198886 54505
rect 198830 54431 198886 54440
rect 200132 16574 200160 70994
rect 200224 50969 200252 198970
rect 200948 198824 201000 198830
rect 200948 198766 201000 198772
rect 200580 198756 200632 198762
rect 200580 198698 200632 198704
rect 200396 198144 200448 198150
rect 200396 198086 200448 198092
rect 200304 192568 200356 192574
rect 200304 192510 200356 192516
rect 200210 50960 200266 50969
rect 200210 50895 200266 50904
rect 200316 48249 200344 192510
rect 200408 59945 200436 198086
rect 200486 195256 200542 195265
rect 200486 195191 200542 195200
rect 200500 62121 200528 195191
rect 200592 71641 200620 198698
rect 200672 198076 200724 198082
rect 200672 198018 200724 198024
rect 200684 78305 200712 198018
rect 200764 192500 200816 192506
rect 200764 192442 200816 192448
rect 200670 78296 200726 78305
rect 200670 78231 200726 78240
rect 200776 76362 200804 192442
rect 200856 152516 200908 152522
rect 200856 152458 200908 152464
rect 200764 76356 200816 76362
rect 200764 76298 200816 76304
rect 200868 74526 200896 152458
rect 200960 138145 200988 198766
rect 200946 138136 201002 138145
rect 200946 138071 201002 138080
rect 200856 74520 200908 74526
rect 200856 74462 200908 74468
rect 200578 71632 200634 71641
rect 200578 71567 200634 71576
rect 201052 68785 201080 199106
rect 201406 150376 201462 150385
rect 201406 150311 201408 150320
rect 201460 150311 201462 150320
rect 201408 150282 201460 150288
rect 201406 71632 201462 71641
rect 201406 71567 201462 71576
rect 201420 71097 201448 71567
rect 201406 71088 201462 71097
rect 201406 71023 201462 71032
rect 201038 68776 201094 68785
rect 201038 68711 201094 68720
rect 201406 68776 201462 68785
rect 201406 68711 201462 68720
rect 201420 68241 201448 68711
rect 201406 68232 201462 68241
rect 201406 68167 201462 68176
rect 200854 67552 200910 67561
rect 200854 67487 200910 67496
rect 200868 67454 200896 67487
rect 200856 67448 200908 67454
rect 200856 67390 200908 67396
rect 201408 67448 201460 67454
rect 201408 67390 201460 67396
rect 201420 66298 201448 67390
rect 201408 66292 201460 66298
rect 201408 66234 201460 66240
rect 200486 62112 200542 62121
rect 200486 62047 200542 62056
rect 201406 62112 201462 62121
rect 201406 62047 201462 62056
rect 201420 61577 201448 62047
rect 201406 61568 201462 61577
rect 201406 61503 201462 61512
rect 200394 59936 200450 59945
rect 200394 59871 200450 59880
rect 200670 56536 200726 56545
rect 200670 56471 200726 56480
rect 200684 56438 200712 56471
rect 200672 56432 200724 56438
rect 200672 56374 200724 56380
rect 201408 56432 201460 56438
rect 201408 56374 201460 56380
rect 201420 55282 201448 56374
rect 201408 55276 201460 55282
rect 201408 55218 201460 55224
rect 201512 52426 201540 200223
rect 201958 200152 202014 200161
rect 201958 200087 202014 200096
rect 201868 198892 201920 198898
rect 201868 198834 201920 198840
rect 201592 194268 201644 194274
rect 201592 194210 201644 194216
rect 201500 52420 201552 52426
rect 201500 52362 201552 52368
rect 201406 50960 201462 50969
rect 201406 50895 201462 50904
rect 201420 50425 201448 50895
rect 201406 50416 201462 50425
rect 201406 50351 201462 50360
rect 201500 49156 201552 49162
rect 201500 49098 201552 49104
rect 200302 48240 200358 48249
rect 200302 48175 200358 48184
rect 201406 48240 201462 48249
rect 201406 48175 201462 48184
rect 201420 47705 201448 48175
rect 201406 47696 201462 47705
rect 201406 47631 201462 47640
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 49098
rect 201604 45529 201632 194210
rect 201776 192976 201828 192982
rect 201776 192918 201828 192924
rect 201684 192636 201736 192642
rect 201684 192578 201736 192584
rect 201696 46889 201724 192578
rect 201788 49609 201816 192918
rect 201880 56574 201908 198834
rect 201972 59362 202000 200087
rect 203064 199368 203116 199374
rect 203064 199310 203116 199316
rect 202970 195392 203026 195401
rect 202970 195327 203026 195336
rect 202052 194064 202104 194070
rect 202052 194006 202104 194012
rect 202064 74458 202092 194006
rect 202880 192704 202932 192710
rect 202880 192646 202932 192652
rect 202328 155236 202380 155242
rect 202328 155178 202380 155184
rect 202142 152416 202198 152425
rect 202142 152351 202198 152360
rect 202052 74452 202104 74458
rect 202052 74394 202104 74400
rect 202064 73914 202092 74394
rect 202052 73908 202104 73914
rect 202052 73850 202104 73856
rect 201960 59356 202012 59362
rect 201960 59298 202012 59304
rect 201868 56568 201920 56574
rect 201868 56510 201920 56516
rect 202156 55214 202184 152351
rect 202236 150272 202288 150278
rect 202236 150214 202288 150220
rect 202248 70378 202276 150214
rect 202340 75886 202368 155178
rect 202788 150408 202840 150414
rect 202786 150376 202788 150385
rect 202840 150376 202842 150385
rect 202786 150311 202842 150320
rect 202328 75880 202380 75886
rect 202328 75822 202380 75828
rect 202236 70372 202288 70378
rect 202236 70314 202288 70320
rect 202788 59356 202840 59362
rect 202788 59298 202840 59304
rect 202800 58750 202828 59298
rect 202788 58744 202840 58750
rect 202788 58686 202840 58692
rect 202788 56568 202840 56574
rect 202788 56510 202840 56516
rect 202800 55894 202828 56510
rect 202788 55888 202840 55894
rect 202788 55830 202840 55836
rect 202156 55186 202368 55214
rect 201774 49600 201830 49609
rect 201774 49535 201830 49544
rect 201682 46880 201738 46889
rect 201682 46815 201738 46824
rect 201590 45520 201646 45529
rect 201590 45455 201646 45464
rect 201604 45121 201632 45455
rect 201590 45112 201646 45121
rect 201590 45047 201646 45056
rect 201592 44940 201644 44946
rect 201592 44882 201644 44888
rect 201604 16574 201632 44882
rect 202340 44169 202368 55186
rect 202788 52420 202840 52426
rect 202788 52362 202840 52368
rect 202800 51814 202828 52362
rect 202788 51808 202840 51814
rect 202788 51750 202840 51756
rect 202786 49600 202842 49609
rect 202786 49535 202842 49544
rect 202800 49065 202828 49535
rect 202786 49056 202842 49065
rect 202786 48991 202842 49000
rect 202786 46880 202842 46889
rect 202786 46815 202842 46824
rect 202800 46209 202828 46815
rect 202786 46200 202842 46209
rect 202786 46135 202842 46144
rect 202326 44160 202382 44169
rect 202326 44095 202382 44104
rect 202340 43625 202368 44095
rect 202892 44033 202920 192646
rect 202984 49337 203012 195327
rect 203076 55214 203104 199310
rect 204720 198212 204772 198218
rect 204720 198154 204772 198160
rect 203154 196752 203210 196761
rect 203154 196687 203210 196696
rect 203168 56409 203196 196687
rect 203340 194200 203392 194206
rect 203340 194142 203392 194148
rect 203248 194132 203300 194138
rect 203248 194074 203300 194080
rect 203260 64802 203288 194074
rect 203352 78402 203380 194142
rect 204352 193112 204404 193118
rect 204352 193054 204404 193060
rect 203432 155372 203484 155378
rect 203432 155314 203484 155320
rect 203340 78396 203392 78402
rect 203340 78338 203392 78344
rect 203248 64796 203300 64802
rect 203248 64738 203300 64744
rect 203260 64190 203288 64738
rect 203248 64184 203300 64190
rect 203248 64126 203300 64132
rect 203444 57934 203472 155314
rect 203524 155304 203576 155310
rect 203524 155246 203576 155252
rect 203536 70310 203564 155246
rect 203708 150068 203760 150074
rect 203708 150010 203760 150016
rect 203616 150000 203668 150006
rect 203616 149942 203668 149948
rect 203628 76809 203656 149942
rect 203720 79082 203748 150010
rect 203708 79076 203760 79082
rect 203708 79018 203760 79024
rect 204364 77081 204392 193054
rect 204442 192672 204498 192681
rect 204442 192607 204498 192616
rect 204456 78169 204484 192607
rect 204536 150204 204588 150210
rect 204536 150146 204588 150152
rect 204442 78160 204498 78169
rect 204442 78095 204498 78104
rect 204350 77072 204406 77081
rect 204350 77007 204406 77016
rect 203614 76800 203670 76809
rect 203614 76735 203670 76744
rect 203616 74316 203668 74322
rect 203616 74258 203668 74264
rect 203524 70304 203576 70310
rect 203524 70246 203576 70252
rect 203432 57928 203484 57934
rect 203432 57870 203484 57876
rect 203154 56400 203210 56409
rect 203154 56335 203210 56344
rect 203064 55208 203116 55214
rect 203064 55150 203116 55156
rect 203076 54534 203104 55150
rect 203064 54528 203116 54534
rect 203064 54470 203116 54476
rect 202970 49328 203026 49337
rect 202970 49263 203026 49272
rect 202878 44024 202934 44033
rect 202878 43959 202934 43968
rect 202326 43616 202382 43625
rect 202326 43551 202382 43560
rect 202892 43489 202920 43959
rect 202878 43480 202934 43489
rect 202878 43415 202934 43424
rect 201604 16546 202736 16574
rect 202708 480 202736 16546
rect 203628 4078 203656 74258
rect 204168 57928 204220 57934
rect 204168 57870 204220 57876
rect 204180 57254 204208 57870
rect 204168 57248 204220 57254
rect 204168 57190 204220 57196
rect 204166 56400 204222 56409
rect 204166 56335 204222 56344
rect 204180 55865 204208 56335
rect 204166 55856 204222 55865
rect 204166 55791 204222 55800
rect 204260 53168 204312 53174
rect 204260 53110 204312 53116
rect 204166 49328 204222 49337
rect 204166 49263 204222 49272
rect 204180 48929 204208 49263
rect 204166 48920 204222 48929
rect 204166 48855 204222 48864
rect 204272 16574 204300 53110
rect 204548 44849 204576 150146
rect 204628 150136 204680 150142
rect 204628 150078 204680 150084
rect 204640 73778 204668 150078
rect 204628 73772 204680 73778
rect 204628 73714 204680 73720
rect 204732 50289 204760 198154
rect 205824 193996 205876 194002
rect 205824 193938 205876 193944
rect 205732 193928 205784 193934
rect 205732 193870 205784 193876
rect 205638 192536 205694 192545
rect 205638 192471 205694 192480
rect 204718 50280 204774 50289
rect 204718 50215 204774 50224
rect 205652 44985 205680 192471
rect 205744 63481 205772 193870
rect 205836 74497 205864 193938
rect 206100 193860 206152 193866
rect 206100 193802 206152 193808
rect 205916 192908 205968 192914
rect 205916 192850 205968 192856
rect 205822 74488 205878 74497
rect 205822 74423 205878 74432
rect 205836 73817 205864 74423
rect 205822 73808 205878 73817
rect 205822 73743 205878 73752
rect 205928 72282 205956 192850
rect 206008 192840 206060 192846
rect 206008 192782 206060 192788
rect 206020 75857 206048 192782
rect 206112 80918 206140 193802
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 206192 149932 206244 149938
rect 206192 149874 206244 149880
rect 206100 80912 206152 80918
rect 206100 80854 206152 80860
rect 206006 75848 206062 75857
rect 206006 75783 206062 75792
rect 206204 75721 206232 149874
rect 206284 149864 206336 149870
rect 206284 149806 206336 149812
rect 206296 78849 206324 149806
rect 206376 149796 206428 149802
rect 206376 149738 206428 149744
rect 206388 79014 206416 149738
rect 206468 146940 206520 146946
rect 206468 146882 206520 146888
rect 206480 80753 206508 146882
rect 580262 146432 580318 146441
rect 580262 146367 580318 146376
rect 464344 140888 464396 140894
rect 464344 140830 464396 140836
rect 327722 139632 327778 139641
rect 327722 139567 327778 139576
rect 234620 80912 234672 80918
rect 234620 80854 234672 80860
rect 206466 80744 206522 80753
rect 206466 80679 206522 80688
rect 206376 79008 206428 79014
rect 206376 78950 206428 78956
rect 206282 78840 206338 78849
rect 206282 78775 206338 78784
rect 211804 76900 211856 76906
rect 211804 76842 211856 76848
rect 206190 75712 206246 75721
rect 206190 75647 206246 75656
rect 205916 72276 205968 72282
rect 205916 72218 205968 72224
rect 207020 65680 207072 65686
rect 207020 65622 207072 65628
rect 205730 63472 205786 63481
rect 205730 63407 205786 63416
rect 205638 44976 205694 44985
rect 205638 44911 205694 44920
rect 204534 44840 204590 44849
rect 204534 44775 204590 44784
rect 205640 36848 205692 36854
rect 205640 36790 205692 36796
rect 205652 16574 205680 36790
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 203616 4072 203668 4078
rect 203616 4014 203668 4020
rect 203892 3936 203944 3942
rect 203892 3878 203944 3884
rect 203904 480 203932 3878
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 65622
rect 209872 58812 209924 58818
rect 209872 58754 209924 58760
rect 208398 46336 208454 46345
rect 208398 46271 208454 46280
rect 208412 16574 208440 46271
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209884 6914 209912 58754
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210976 4004 211028 4010
rect 210976 3946 211028 3952
rect 210988 480 211016 3946
rect 211816 3942 211844 76842
rect 224224 76832 224276 76838
rect 224224 76774 224276 76780
rect 216680 75540 216732 75546
rect 216680 75482 216732 75488
rect 213918 67144 213974 67153
rect 213918 67079 213974 67088
rect 213932 16574 213960 67079
rect 215300 51876 215352 51882
rect 215300 51818 215352 51824
rect 213932 16546 214512 16574
rect 213366 7576 213422 7585
rect 213366 7511 213422 7520
rect 211804 3936 211856 3942
rect 211804 3878 211856 3884
rect 212172 3868 212224 3874
rect 212172 3810 212224 3816
rect 212184 480 212212 3810
rect 213380 480 213408 7511
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 51818
rect 216692 16574 216720 75482
rect 223580 75472 223632 75478
rect 223580 75414 223632 75420
rect 218058 71360 218114 71369
rect 218058 71295 218114 71304
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 71295
rect 220818 68368 220874 68377
rect 220818 68303 220874 68312
rect 218152 49088 218204 49094
rect 218152 49030 218204 49036
rect 218164 16574 218192 49030
rect 219440 23044 219492 23050
rect 219440 22986 219492 22992
rect 219452 16574 219480 22986
rect 220832 16574 220860 68303
rect 222200 47728 222252 47734
rect 222200 47670 222252 47676
rect 222212 16574 222240 47670
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 75414
rect 224236 4010 224264 76774
rect 224960 64320 225012 64326
rect 224960 64262 225012 64268
rect 224972 16574 225000 64262
rect 227720 62892 227772 62898
rect 227720 62834 227772 62840
rect 226340 18896 226392 18902
rect 226340 18838 226392 18844
rect 224972 16546 225184 16574
rect 224224 4004 224276 4010
rect 224224 3946 224276 3952
rect 225156 480 225184 16546
rect 226352 480 226380 18838
rect 227732 16574 227760 62834
rect 231858 56128 231914 56137
rect 231858 56063 231914 56072
rect 229098 42120 229154 42129
rect 229098 42055 229154 42064
rect 229112 16574 229140 42055
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 227536 9240 227588 9246
rect 227536 9182 227588 9188
rect 227548 480 227576 9182
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231032 3936 231084 3942
rect 231032 3878 231084 3884
rect 231044 480 231072 3878
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 56063
rect 233240 43580 233292 43586
rect 233240 43522 233292 43528
rect 233252 16574 233280 43522
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 80854
rect 252560 80844 252612 80850
rect 252560 80786 252612 80792
rect 238760 80232 238812 80238
rect 238760 80174 238812 80180
rect 237380 74248 237432 74254
rect 237380 74190 237432 74196
rect 236000 57384 236052 57390
rect 236000 57326 236052 57332
rect 236012 16574 236040 57326
rect 237392 16574 237420 74190
rect 238772 16574 238800 80174
rect 247684 74180 247736 74186
rect 247684 74122 247736 74128
rect 242164 72956 242216 72962
rect 242164 72898 242216 72904
rect 241520 17536 241572 17542
rect 241520 17478 241572 17484
rect 241532 16574 241560 17478
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234620 10532 234672 10538
rect 234620 10474 234672 10480
rect 234632 480 234660 10474
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240508 3868 240560 3874
rect 240508 3810 240560 3816
rect 240520 480 240548 3810
rect 241716 480 241744 16546
rect 242176 3874 242204 72898
rect 242900 67040 242952 67046
rect 242900 66982 242952 66988
rect 242164 3868 242216 3874
rect 242164 3810 242216 3816
rect 242912 480 242940 66982
rect 245658 61976 245714 61985
rect 245658 61911 245714 61920
rect 242990 29608 243046 29617
rect 242990 29543 243046 29552
rect 243004 16574 243032 29543
rect 245672 16574 245700 61911
rect 243004 16546 244136 16574
rect 245672 16546 245976 16574
rect 244108 480 244136 16546
rect 245200 12028 245252 12034
rect 245200 11970 245252 11976
rect 245212 480 245240 11970
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247696 4078 247724 74122
rect 249798 58984 249854 58993
rect 249798 58919 249854 58928
rect 249812 16574 249840 58919
rect 251180 39636 251232 39642
rect 251180 39578 251232 39584
rect 249812 16546 250024 16574
rect 247684 4072 247736 4078
rect 247684 4014 247736 4020
rect 248788 4072 248840 4078
rect 248788 4014 248840 4020
rect 247592 4004 247644 4010
rect 247592 3946 247644 3952
rect 247604 480 247632 3946
rect 248800 480 248828 4014
rect 249996 480 250024 16546
rect 251192 480 251220 39578
rect 252572 16574 252600 80786
rect 270500 80776 270552 80782
rect 270500 80718 270552 80724
rect 255964 78328 256016 78334
rect 255964 78270 256016 78276
rect 255976 73982 256004 78270
rect 264242 77888 264298 77897
rect 264242 77823 264298 77832
rect 260840 76764 260892 76770
rect 260840 76706 260892 76712
rect 255320 73976 255372 73982
rect 255320 73918 255372 73924
rect 255964 73976 256016 73982
rect 255964 73918 256016 73924
rect 253940 54664 253992 54670
rect 253940 54606 253992 54612
rect 253952 16574 253980 54606
rect 255332 16574 255360 73918
rect 256698 64424 256754 64433
rect 256698 64359 256754 64368
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 16108 252428 16114
rect 252376 16050 252428 16056
rect 252388 480 252416 16050
rect 253492 480 253520 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 64359
rect 259458 63336 259514 63345
rect 259458 63271 259514 63280
rect 258080 28552 258132 28558
rect 258080 28494 258132 28500
rect 258092 16574 258120 28494
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 259472 3398 259500 63271
rect 260852 16574 260880 76706
rect 264256 73846 264284 77823
rect 261484 73840 261536 73846
rect 261484 73782 261536 73788
rect 264244 73840 264296 73846
rect 264244 73782 264296 73788
rect 269118 73808 269174 73817
rect 260852 16546 261432 16574
rect 259552 5092 259604 5098
rect 259552 5034 259604 5040
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 259564 2530 259592 5034
rect 261404 3482 261432 16546
rect 261496 3942 261524 73782
rect 269118 73743 269174 73752
rect 263598 60344 263654 60353
rect 263598 60279 263654 60288
rect 263612 16574 263640 60279
rect 267740 47660 267792 47666
rect 267740 47602 267792 47608
rect 266360 35420 266412 35426
rect 266360 35362 266412 35368
rect 266372 16574 266400 35362
rect 263612 16546 264192 16574
rect 266372 16546 266584 16574
rect 261484 3936 261536 3942
rect 261484 3878 261536 3884
rect 262956 3936 263008 3942
rect 262956 3878 263008 3884
rect 261404 3454 261800 3482
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 259472 2502 259592 2530
rect 259472 480 259500 2502
rect 260668 480 260696 3334
rect 261772 480 261800 3454
rect 262968 480 262996 3878
rect 264164 480 264192 16546
rect 264978 13016 265034 13025
rect 264978 12951 265034 12960
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 12951
rect 266556 480 266584 16546
rect 267752 480 267780 47602
rect 267832 38208 267884 38214
rect 267832 38150 267884 38156
rect 267844 16574 267872 38150
rect 269132 16574 269160 73743
rect 270512 16574 270540 80718
rect 288440 80708 288492 80714
rect 288440 80650 288492 80656
rect 287704 78396 287756 78402
rect 287704 78338 287756 78344
rect 284300 74112 284352 74118
rect 284300 74054 284352 74060
rect 274640 65612 274692 65618
rect 274640 65554 274692 65560
rect 273260 44872 273312 44878
rect 273260 44814 273312 44820
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 14748 272484 14754
rect 272432 14690 272484 14696
rect 272444 480 272472 14690
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 44814
rect 274652 16574 274680 65554
rect 277398 61840 277454 61849
rect 277398 61775 277454 61784
rect 276020 40996 276072 41002
rect 276020 40938 276072 40944
rect 276032 16574 276060 40938
rect 277412 16574 277440 61775
rect 281538 58848 281594 58857
rect 281538 58783 281594 58792
rect 278780 32632 278832 32638
rect 278780 32574 278832 32580
rect 278792 16574 278820 32574
rect 280160 20256 280212 20262
rect 280160 20198 280212 20204
rect 280172 16574 280200 20198
rect 274652 16546 274864 16574
rect 276032 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 274836 480 274864 16546
rect 276020 6384 276072 6390
rect 276020 6326 276072 6332
rect 276032 480 276060 6326
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 58783
rect 282918 26888 282974 26897
rect 282918 26823 282974 26832
rect 282932 16574 282960 26823
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 480 284340 74054
rect 285680 46368 285732 46374
rect 285680 46310 285732 46316
rect 284392 24404 284444 24410
rect 284392 24346 284444 24352
rect 284404 16574 284432 24346
rect 285692 16574 285720 46310
rect 287716 20126 287744 78338
rect 287060 20120 287112 20126
rect 287060 20062 287112 20068
rect 287704 20120 287756 20126
rect 287704 20062 287756 20068
rect 287072 16574 287100 20062
rect 288452 16574 288480 80650
rect 302240 80164 302292 80170
rect 302240 80106 302292 80112
rect 289820 76016 289872 76022
rect 289820 75958 289872 75964
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 75958
rect 296720 75948 296772 75954
rect 296720 75890 296772 75896
rect 295340 66972 295392 66978
rect 295340 66914 295392 66920
rect 292578 63200 292634 63209
rect 292578 63135 292634 63144
rect 291200 20188 291252 20194
rect 291200 20130 291252 20136
rect 291212 16574 291240 20130
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 63135
rect 293960 50380 294012 50386
rect 293960 50322 294012 50328
rect 292672 42288 292724 42294
rect 292672 42230 292724 42236
rect 292684 16574 292712 42230
rect 293972 16574 294000 50322
rect 295352 16574 295380 66914
rect 296732 16574 296760 75890
rect 301504 72888 301556 72894
rect 301504 72830 301556 72836
rect 299478 60208 299534 60217
rect 299478 60143 299534 60152
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 298468 3868 298520 3874
rect 298468 3810 298520 3816
rect 298480 480 298508 3810
rect 299492 3482 299520 60143
rect 299572 34060 299624 34066
rect 299572 34002 299624 34008
rect 299584 3874 299612 34002
rect 300860 18828 300912 18834
rect 300860 18770 300912 18776
rect 300872 6914 300900 18770
rect 301516 16574 301544 72830
rect 302252 16574 302280 80106
rect 306378 79792 306434 79801
rect 306378 79727 306434 79736
rect 305000 72820 305052 72826
rect 305000 72762 305052 72768
rect 303620 36780 303672 36786
rect 303620 36722 303672 36728
rect 303632 16574 303660 36722
rect 305012 16574 305040 72762
rect 301516 16546 301636 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 300872 6886 301544 6914
rect 299572 3868 299624 3874
rect 299572 3810 299624 3816
rect 300768 3868 300820 3874
rect 300768 3810 300820 3816
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3810
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 6886
rect 301608 4146 301636 16546
rect 301596 4140 301648 4146
rect 301596 4082 301648 4088
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 79727
rect 324320 78260 324372 78266
rect 324320 78202 324372 78208
rect 311164 72752 311216 72758
rect 311164 72694 311216 72700
rect 309138 61704 309194 61713
rect 309138 61639 309194 61648
rect 307852 42220 307904 42226
rect 307852 42162 307904 42168
rect 307864 16574 307892 42162
rect 309152 16574 309180 61639
rect 310520 25832 310572 25838
rect 310520 25774 310572 25780
rect 310532 16574 310560 25774
rect 307864 16546 307984 16574
rect 309152 16546 309824 16574
rect 310532 16546 311112 16574
rect 307956 480 307984 16546
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 309060 480 309088 4082
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311084 3482 311112 16546
rect 311176 3874 311204 72694
rect 318800 72684 318852 72690
rect 318800 72626 318852 72632
rect 313278 57488 313334 57497
rect 313278 57423 313334 57432
rect 313292 16574 313320 57423
rect 315302 45248 315358 45257
rect 315302 45183 315358 45192
rect 313292 16546 313872 16574
rect 311164 3868 311216 3874
rect 311164 3810 311216 3816
rect 312636 3868 312688 3874
rect 312636 3810 312688 3816
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 312648 480 312676 3810
rect 313844 480 313872 16546
rect 314660 14680 314712 14686
rect 314660 14622 314712 14628
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 14622
rect 315316 4146 315344 45183
rect 317420 31340 317472 31346
rect 317420 31282 317472 31288
rect 317432 16574 317460 31282
rect 318812 16574 318840 72626
rect 320178 53544 320234 53553
rect 320178 53479 320234 53488
rect 320192 16574 320220 53479
rect 322940 40928 322992 40934
rect 322940 40870 322992 40876
rect 321560 35352 321612 35358
rect 321560 35294 321612 35300
rect 321572 16574 321600 35294
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316224 7812 316276 7818
rect 316224 7754 316276 7760
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316236 480 316264 7754
rect 317328 4140 317380 4146
rect 317328 4082 317380 4088
rect 317340 480 317368 4082
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 40870
rect 324332 3210 324360 78202
rect 327736 73166 327764 139567
rect 464356 86970 464384 140830
rect 485044 140820 485096 140826
rect 485044 140762 485096 140768
rect 464344 86964 464396 86970
rect 464344 86906 464396 86912
rect 382278 80200 382334 80209
rect 382278 80135 382334 80144
rect 380900 80096 380952 80102
rect 380900 80038 380952 80044
rect 337384 78192 337436 78198
rect 337384 78134 337436 78140
rect 327724 73160 327776 73166
rect 327724 73102 327776 73108
rect 324964 72616 325016 72622
rect 324964 72558 325016 72564
rect 324412 13252 324464 13258
rect 324412 13194 324464 13200
rect 324424 3398 324452 13194
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 324976 3330 325004 72558
rect 332600 72548 332652 72554
rect 332600 72490 332652 72496
rect 331218 58712 331274 58721
rect 331218 58647 331274 58656
rect 328460 24336 328512 24342
rect 328460 24278 328512 24284
rect 328472 16574 328500 24278
rect 329104 21684 329156 21690
rect 329104 21626 329156 21632
rect 328472 16546 328776 16574
rect 328000 3800 328052 3806
rect 328000 3742 328052 3748
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324964 3324 325016 3330
rect 324964 3266 325016 3272
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 326804 3324 326856 3330
rect 326804 3266 326856 3272
rect 326816 480 326844 3266
rect 328012 480 328040 3742
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 329116 3398 329144 21626
rect 329104 3392 329156 3398
rect 329104 3334 329156 3340
rect 330392 3392 330444 3398
rect 330392 3334 330444 3340
rect 330404 480 330432 3334
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 58647
rect 332612 3398 332640 72490
rect 333980 54596 334032 54602
rect 333980 54538 334032 54544
rect 332692 29844 332744 29850
rect 332692 29786 332744 29792
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 29786
rect 333992 16574 334020 54538
rect 337396 21622 337424 78134
rect 353300 76696 353352 76702
rect 353300 76638 353352 76644
rect 347780 74044 347832 74050
rect 347780 73986 347832 73992
rect 346400 65544 346452 65550
rect 346400 65486 346452 65492
rect 340880 62824 340932 62830
rect 340880 62766 340932 62772
rect 338118 60072 338174 60081
rect 338118 60007 338174 60016
rect 336740 21616 336792 21622
rect 336740 21558 336792 21564
rect 337384 21616 337436 21622
rect 337384 21558 337436 21564
rect 336752 16574 336780 21558
rect 338132 16574 338160 60007
rect 339500 28484 339552 28490
rect 339500 28426 339552 28432
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336278 6216 336334 6225
rect 336278 6151 336334 6160
rect 336292 480 336320 6151
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 28426
rect 340892 1834 340920 62766
rect 345020 57316 345072 57322
rect 345020 57258 345072 57264
rect 340972 33992 341024 33998
rect 340972 33934 341024 33940
rect 340880 1828 340932 1834
rect 340880 1770 340932 1776
rect 340984 480 341012 33934
rect 342904 21548 342956 21554
rect 342904 21490 342956 21496
rect 342916 16574 342944 21490
rect 345032 16574 345060 57258
rect 346412 16574 346440 65486
rect 347792 16574 347820 73986
rect 349160 55956 349212 55962
rect 349160 55898 349212 55904
rect 342916 16546 343036 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 342904 11960 342956 11966
rect 342904 11902 342956 11908
rect 342168 1828 342220 1834
rect 342168 1770 342220 1776
rect 342180 480 342208 1770
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 11902
rect 343008 3398 343036 16546
rect 342996 3392 343048 3398
rect 342996 3334 343048 3340
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 344572 480 344600 3334
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3210 349200 55898
rect 351918 53408 351974 53417
rect 351918 53343 351974 53352
rect 350540 31272 350592 31278
rect 350540 31214 350592 31220
rect 350552 16574 350580 31214
rect 351932 16574 351960 53343
rect 353312 16574 353340 76638
rect 374000 76628 374052 76634
rect 374000 76570 374052 76576
rect 354680 69760 354732 69766
rect 354680 69702 354732 69708
rect 354692 16574 354720 69702
rect 367100 68468 367152 68474
rect 367100 68410 367152 68416
rect 358820 64252 358872 64258
rect 358820 64194 358872 64200
rect 356058 50688 356114 50697
rect 356058 50623 356114 50632
rect 356072 16574 356100 50623
rect 357532 39568 357584 39574
rect 357532 39510 357584 39516
rect 356704 32564 356756 32570
rect 356704 32506 356756 32512
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 349252 10464 349304 10470
rect 349252 10406 349304 10412
rect 349264 3398 349292 10406
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 356716 3398 356744 32506
rect 357544 3806 357572 39510
rect 358832 16574 358860 64194
rect 362958 58576 363014 58585
rect 362958 58511 363014 58520
rect 361580 43512 361632 43518
rect 361580 43454 361632 43460
rect 361592 16574 361620 43454
rect 362972 16574 363000 58511
rect 364982 54632 365038 54641
rect 364982 54567 365038 54576
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 357532 3800 357584 3806
rect 357532 3742 357584 3748
rect 358728 3800 358780 3806
rect 358728 3742 358780 3748
rect 356704 3392 356756 3398
rect 356704 3334 356756 3340
rect 357532 3392 357584 3398
rect 357532 3334 357584 3340
rect 357544 480 357572 3334
rect 358740 480 358768 3742
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 16040 361172 16046
rect 361120 15982 361172 15988
rect 361132 480 361160 15982
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 15972 364668 15978
rect 364616 15914 364668 15920
rect 364628 480 364656 15914
rect 364996 3398 365024 54567
rect 365812 22976 365864 22982
rect 365812 22918 365864 22924
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 22918
rect 367112 16574 367140 68410
rect 369858 52048 369914 52057
rect 369858 51983 369914 51992
rect 368480 38140 368532 38146
rect 368480 38082 368532 38088
rect 368492 16574 368520 38082
rect 369872 16574 369900 51983
rect 372620 20052 372672 20058
rect 372620 19994 372672 20000
rect 372632 16574 372660 19994
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371700 9172 371752 9178
rect 371700 9114 371752 9120
rect 371712 480 371740 9114
rect 372908 480 372936 16546
rect 374012 3398 374040 76570
rect 375380 72480 375432 72486
rect 375380 72422 375432 72428
rect 374090 51912 374146 51921
rect 374090 51847 374146 51856
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 51847
rect 375392 16574 375420 72422
rect 378784 29776 378836 29782
rect 378784 29718 378836 29724
rect 375392 16546 376064 16574
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377680 3732 377732 3738
rect 377680 3674 377732 3680
rect 377692 480 377720 3674
rect 378796 3398 378824 29718
rect 380912 16574 380940 80038
rect 380912 16546 381216 16574
rect 378876 7744 378928 7750
rect 378876 7686 378928 7692
rect 378784 3392 378836 3398
rect 378784 3334 378836 3340
rect 378888 480 378916 7686
rect 379980 3392 380032 3398
rect 379980 3334 380032 3340
rect 379992 480 380020 3334
rect 381188 480 381216 16546
rect 382292 3330 382320 80135
rect 483020 78940 483072 78946
rect 483020 78882 483072 78888
rect 393320 78124 393372 78130
rect 393320 78066 393372 78072
rect 391940 76560 391992 76566
rect 389178 76528 389234 76537
rect 391940 76502 391992 76508
rect 389178 76463 389234 76472
rect 382922 55992 382978 56001
rect 382922 55927 382978 55936
rect 382372 5024 382424 5030
rect 382372 4966 382424 4972
rect 382280 3324 382332 3330
rect 382280 3266 382332 3272
rect 382384 480 382412 4966
rect 382936 3398 382964 55927
rect 387798 53272 387854 53281
rect 387798 53207 387854 53216
rect 385040 33924 385092 33930
rect 385040 33866 385092 33872
rect 385052 16574 385080 33866
rect 385052 16546 386000 16574
rect 382924 3392 382976 3398
rect 382924 3334 382976 3340
rect 384764 3392 384816 3398
rect 384764 3334 384816 3340
rect 383568 3324 383620 3330
rect 383568 3266 383620 3272
rect 383580 480 383608 3266
rect 384776 480 384804 3334
rect 385972 480 386000 16546
rect 387156 9104 387208 9110
rect 387156 9046 387208 9052
rect 387168 480 387196 9046
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 53207
rect 389192 16574 389220 76463
rect 390558 50552 390614 50561
rect 390558 50487 390614 50496
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 2514 390600 50487
rect 391952 16574 391980 76502
rect 393332 16574 393360 78066
rect 400864 78056 400916 78062
rect 400864 77998 400916 78004
rect 400220 77988 400272 77994
rect 400220 77930 400272 77936
rect 394700 61464 394752 61470
rect 394700 61406 394752 61412
rect 394712 16574 394740 61406
rect 398840 60104 398892 60110
rect 398840 60046 398892 60052
rect 396080 60036 396132 60042
rect 396080 59978 396132 59984
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 390652 11892 390704 11898
rect 390652 11834 390704 11840
rect 390560 2508 390612 2514
rect 390560 2450 390612 2456
rect 390664 480 390692 11834
rect 391848 2508 391900 2514
rect 391848 2450 391900 2456
rect 391860 480 391888 2450
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 59978
rect 397460 28416 397512 28422
rect 397460 28358 397512 28364
rect 397472 16574 397500 28358
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3210 398880 60046
rect 398932 14612 398984 14618
rect 398932 14554 398984 14560
rect 398944 3398 398972 14554
rect 400232 6914 400260 77930
rect 400876 15978 400904 77998
rect 454684 75336 454736 75342
rect 454684 75278 454736 75284
rect 475382 75304 475438 75313
rect 446404 73908 446456 73914
rect 446404 73850 446456 73856
rect 430580 69692 430632 69698
rect 430580 69634 430632 69640
rect 412640 68400 412692 68406
rect 412640 68342 412692 68348
rect 402980 66904 403032 66910
rect 402980 66846 403032 66852
rect 400954 51776 401010 51785
rect 400954 51711 401010 51720
rect 400864 15972 400916 15978
rect 400864 15914 400916 15920
rect 400232 6886 400904 6914
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 6886
rect 400968 3262 400996 51711
rect 402992 16574 403020 66846
rect 405738 49192 405794 49201
rect 405738 49127 405794 49136
rect 405752 16574 405780 49127
rect 408498 47832 408554 47841
rect 408498 47767 408554 47776
rect 408512 16574 408540 47767
rect 409880 27124 409932 27130
rect 409880 27066 409932 27072
rect 409892 16574 409920 27066
rect 402992 16546 403664 16574
rect 405752 16546 406056 16574
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 400956 3256 401008 3262
rect 400956 3198 401008 3204
rect 402520 3256 402572 3262
rect 402520 3198 402572 3204
rect 402532 480 402560 3198
rect 403636 480 403664 16546
rect 404360 14544 404412 14550
rect 404360 14486 404412 14492
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 14486
rect 406028 480 406056 16546
rect 407212 13184 407264 13190
rect 407212 13126 407264 13132
rect 407224 480 407252 13126
rect 408408 3664 408460 3670
rect 408408 3606 408460 3612
rect 408420 480 408448 3606
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411904 6316 411956 6322
rect 411904 6258 411956 6264
rect 411916 480 411944 6258
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 68342
rect 423678 67008 423734 67017
rect 423678 66943 423734 66952
rect 414662 63064 414718 63073
rect 414662 62999 414718 63008
rect 414296 6248 414348 6254
rect 414296 6190 414348 6196
rect 414308 480 414336 6190
rect 414676 3398 414704 62999
rect 418802 57352 418858 57361
rect 418802 57287 418858 57296
rect 418160 46300 418212 46306
rect 418160 46242 418212 46248
rect 416780 22908 416832 22914
rect 416780 22850 416832 22856
rect 415492 21480 415544 21486
rect 415492 21422 415544 21428
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 21422
rect 416792 16574 416820 22850
rect 418172 16574 418200 46242
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3398 418844 57287
rect 420920 31204 420972 31210
rect 420920 31146 420972 31152
rect 418804 3392 418856 3398
rect 418804 3334 418856 3340
rect 420184 3392 420236 3398
rect 420184 3334 420236 3340
rect 420196 480 420224 3334
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 31146
rect 422576 4956 422628 4962
rect 422576 4898 422628 4904
rect 422588 480 422616 4898
rect 423692 2922 423720 66943
rect 423770 54496 423826 54505
rect 423770 54431 423826 54440
rect 423680 2916 423732 2922
rect 423680 2858 423732 2864
rect 423784 480 423812 54431
rect 426440 43444 426492 43450
rect 426440 43386 426492 43392
rect 425060 17468 425112 17474
rect 425060 17410 425112 17416
rect 425072 16574 425100 17410
rect 426452 16574 426480 43386
rect 427820 40860 427872 40866
rect 427820 40802 427872 40808
rect 427832 16574 427860 40802
rect 429200 27056 429252 27062
rect 429200 26998 429252 27004
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 424968 2916 425020 2922
rect 424968 2858 425020 2864
rect 424980 480 425008 2858
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 26998
rect 430592 16574 430620 69634
rect 440238 61568 440294 61577
rect 440238 61503 440294 61512
rect 433338 53136 433394 53145
rect 433338 53071 433394 53080
rect 431960 32496 432012 32502
rect 431960 32438 432012 32444
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 3398 432000 32438
rect 433352 16574 433380 53071
rect 437478 50416 437534 50425
rect 437478 50351 437534 50360
rect 436100 25764 436152 25770
rect 436100 25706 436152 25712
rect 436112 16574 436140 25706
rect 433352 16546 434024 16574
rect 436112 16546 436784 16574
rect 432052 15904 432104 15910
rect 432052 15846 432104 15852
rect 431960 3392 432012 3398
rect 431960 3334 432012 3340
rect 432064 480 432092 15846
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 435088 11824 435140 11830
rect 435088 11766 435140 11772
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 11766
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 50351
rect 439136 10396 439188 10402
rect 439136 10338 439188 10344
rect 439148 480 439176 10338
rect 440252 2650 440280 61503
rect 444378 47696 444434 47705
rect 444378 47631 444434 47640
rect 440332 21412 440384 21418
rect 440332 21354 440384 21360
rect 440240 2644 440292 2650
rect 440240 2586 440292 2592
rect 440344 480 440372 21354
rect 443000 19984 443052 19990
rect 443000 19926 443052 19932
rect 441620 17400 441672 17406
rect 441620 17342 441672 17348
rect 441632 16574 441660 17342
rect 443012 16574 443040 19926
rect 444392 16574 444420 47631
rect 445760 17332 445812 17338
rect 445760 17274 445812 17280
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 441528 2644 441580 2650
rect 441528 2586 441580 2592
rect 441540 480 441568 2586
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 17274
rect 446416 3398 446444 73850
rect 453304 68332 453356 68338
rect 453304 68274 453356 68280
rect 448520 58744 448572 58750
rect 448520 58686 448572 58692
rect 446404 3392 446456 3398
rect 446404 3334 446456 3340
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 447428 480 447456 3334
rect 448532 3210 448560 58686
rect 450544 55888 450596 55894
rect 450544 55830 450596 55836
rect 448610 43616 448666 43625
rect 448610 43551 448666 43560
rect 448624 3398 448652 43551
rect 449900 24268 449952 24274
rect 449900 24210 449952 24216
rect 449912 16574 449940 24210
rect 449912 16546 450492 16574
rect 450464 3482 450492 16546
rect 450556 4146 450584 55830
rect 452660 29708 452712 29714
rect 452660 29650 452712 29656
rect 452672 6914 452700 29650
rect 453316 16574 453344 68274
rect 453316 16546 453436 16574
rect 452672 6886 453344 6914
rect 450544 4140 450596 4146
rect 450544 4082 450596 4088
rect 451004 4140 451056 4146
rect 451004 4082 451056 4088
rect 450464 3454 450952 3482
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 3454
rect 451016 3330 451044 4082
rect 451004 3324 451056 3330
rect 451004 3266 451056 3272
rect 452108 3324 452160 3330
rect 452108 3266 452160 3272
rect 452120 480 452148 3266
rect 453316 480 453344 6886
rect 453408 3398 453436 16546
rect 454696 3670 454724 75278
rect 475382 75239 475438 75248
rect 456800 73976 456852 73982
rect 456800 73918 456852 73924
rect 455418 49056 455474 49065
rect 455418 48991 455474 49000
rect 455432 16574 455460 48991
rect 455432 16546 455736 16574
rect 454684 3664 454736 3670
rect 454684 3606 454736 3612
rect 453396 3392 453448 3398
rect 453396 3334 453448 3340
rect 454500 3392 454552 3398
rect 454500 3334 454552 3340
rect 454512 480 454540 3334
rect 455708 480 455736 16546
rect 456812 3398 456840 73918
rect 472624 64184 472676 64190
rect 472624 64126 472676 64132
rect 459560 61396 459612 61402
rect 459560 61338 459612 61344
rect 458178 45112 458234 45121
rect 458178 45047 458234 45056
rect 458192 16574 458220 45047
rect 459572 16574 459600 61338
rect 468484 54528 468536 54534
rect 468484 54470 468536 54476
rect 464344 51808 464396 51814
rect 464344 51750 464396 51756
rect 463700 46232 463752 46238
rect 462318 46200 462374 46209
rect 463700 46174 463752 46180
rect 462318 46135 462374 46144
rect 460940 33856 460992 33862
rect 460940 33798 460992 33804
rect 460952 16574 460980 33798
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 456892 9036 456944 9042
rect 456892 8978 456944 8984
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 8978
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 46135
rect 463712 16574 463740 46174
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 464356 3058 464384 51750
rect 466458 48920 466514 48929
rect 466458 48855 466514 48864
rect 465172 20120 465224 20126
rect 465172 20062 465224 20068
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 20062
rect 466472 16574 466500 48855
rect 466472 16546 467512 16574
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 16546
rect 468496 3602 468524 54470
rect 470600 28348 470652 28354
rect 470600 28290 470652 28296
rect 468300 3596 468352 3602
rect 468300 3538 468352 3544
rect 468484 3596 468536 3602
rect 468484 3538 468536 3544
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468312 354 468340 3538
rect 469876 480 469904 3538
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 28290
rect 471980 21616 472032 21622
rect 471980 21558 472032 21564
rect 471992 16574 472020 21558
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 472636 3602 472664 64126
rect 473452 57248 473504 57254
rect 473452 57190 473504 57196
rect 473464 16574 473492 57190
rect 474740 31136 474792 31142
rect 474740 31078 474792 31084
rect 474752 16574 474780 31078
rect 473464 16546 474136 16574
rect 474752 16546 475332 16574
rect 472624 3596 472676 3602
rect 472624 3538 472676 3544
rect 473452 3596 473504 3602
rect 473452 3538 473504 3544
rect 473464 480 473492 3538
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475304 3482 475332 16546
rect 475396 3602 475424 75239
rect 480260 70508 480312 70514
rect 480260 70450 480312 70456
rect 476118 43480 476174 43489
rect 476118 43415 476174 43424
rect 476132 16574 476160 43415
rect 477500 39500 477552 39506
rect 477500 39442 477552 39448
rect 477512 16574 477540 39442
rect 480272 16574 480300 70450
rect 481638 55856 481694 55865
rect 481638 55791 481694 55800
rect 481652 16574 481680 55791
rect 483032 16574 483060 78882
rect 484400 39432 484452 39438
rect 484400 39374 484452 39380
rect 484412 16574 484440 39374
rect 485056 20670 485084 140762
rect 576122 139496 576178 139505
rect 576122 139431 576178 139440
rect 525800 79348 525852 79354
rect 525800 79290 525852 79296
rect 500960 78872 501012 78878
rect 500960 78814 501012 78820
rect 494058 71224 494114 71233
rect 494058 71159 494114 71168
rect 489920 58676 489972 58682
rect 489920 58618 489972 58624
rect 486424 49020 486476 49026
rect 486424 48962 486476 48968
rect 485044 20664 485096 20670
rect 485044 20606 485096 20612
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 481652 16546 481772 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 475384 3596 475436 3602
rect 475384 3538 475436 3544
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 478880 15972 478932 15978
rect 478880 15914 478932 15920
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 15914
rect 480548 480 480576 16546
rect 481744 480 481772 16546
rect 482836 7676 482888 7682
rect 482836 7618 482888 7624
rect 482848 480 482876 7618
rect 484044 480 484072 16546
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486332 4888 486384 4894
rect 486332 4830 486384 4836
rect 486344 2530 486372 4830
rect 486436 3398 486464 48962
rect 488540 38072 488592 38078
rect 488540 38014 488592 38020
rect 488552 16574 488580 38014
rect 488552 16546 488856 16574
rect 486424 3392 486476 3398
rect 486424 3334 486476 3340
rect 487620 3392 487672 3398
rect 487620 3334 487672 3340
rect 486344 2502 486464 2530
rect 486436 480 486464 2502
rect 487632 480 487660 3334
rect 488828 480 488856 16546
rect 489932 480 489960 58618
rect 490012 36712 490064 36718
rect 490012 36654 490064 36660
rect 490024 16574 490052 36654
rect 491300 35284 491352 35290
rect 491300 35226 491352 35232
rect 491312 16574 491340 35226
rect 492680 17264 492732 17270
rect 492680 17206 492732 17212
rect 492692 16574 492720 17206
rect 494072 16574 494100 71159
rect 498198 69592 498254 69601
rect 498198 69527 498254 69536
rect 496082 66872 496138 66881
rect 496082 66807 496138 66816
rect 495440 33788 495492 33794
rect 495440 33730 495492 33736
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 33730
rect 496096 3466 496124 66807
rect 496084 3460 496136 3466
rect 496084 3402 496136 3408
rect 497096 3460 497148 3466
rect 497096 3402 497148 3408
rect 497108 480 497136 3402
rect 498212 480 498240 69527
rect 498292 42152 498344 42158
rect 498292 42094 498344 42100
rect 498304 16574 498332 42094
rect 500972 16574 501000 78814
rect 523132 78804 523184 78810
rect 523132 78746 523184 78752
rect 504364 75404 504416 75410
rect 504364 75346 504416 75352
rect 502340 36644 502392 36650
rect 502340 36586 502392 36592
rect 502352 16574 502380 36586
rect 498304 16546 498976 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500592 3664 500644 3670
rect 500592 3606 500644 3612
rect 500604 480 500632 3606
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 503720 14476 503772 14482
rect 503720 14418 503772 14424
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 14418
rect 504376 3534 504404 75346
rect 511264 75268 511316 75274
rect 511264 75210 511316 75216
rect 507858 65512 507914 65521
rect 507858 65447 507914 65456
rect 506572 29640 506624 29646
rect 506572 29582 506624 29588
rect 506584 6914 506612 29582
rect 507872 16574 507900 65447
rect 509240 28280 509292 28286
rect 509240 28222 509292 28228
rect 509252 16574 509280 28222
rect 511276 16574 511304 75210
rect 521660 75200 521712 75206
rect 521660 75142 521712 75148
rect 518900 73840 518952 73846
rect 518900 73782 518952 73788
rect 511998 64288 512054 64297
rect 511998 64223 512054 64232
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 511276 16546 511396 16574
rect 506492 6886 506612 6914
rect 504364 3528 504416 3534
rect 504364 3470 504416 3476
rect 505376 3392 505428 3398
rect 505376 3334 505428 3340
rect 505388 480 505416 3334
rect 506492 480 506520 6886
rect 507676 3528 507728 3534
rect 507676 3470 507728 3476
rect 507688 480 507716 3470
rect 508884 480 508912 16546
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511264 13116 511316 13122
rect 511264 13058 511316 13064
rect 511276 480 511304 13058
rect 511368 3194 511396 16546
rect 511356 3188 511408 3194
rect 511356 3130 511408 3136
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 64223
rect 514022 62928 514078 62937
rect 514022 62863 514078 62872
rect 513380 26988 513432 26994
rect 513380 26930 513432 26936
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 26930
rect 514036 3058 514064 62863
rect 516140 40792 516192 40798
rect 516140 40734 516192 40740
rect 516152 16574 516180 40734
rect 518912 16574 518940 73782
rect 520922 47560 520978 47569
rect 520922 47495 520978 47504
rect 520280 25696 520332 25702
rect 520280 25638 520332 25644
rect 516152 16546 517192 16574
rect 518912 16546 519584 16574
rect 514760 3188 514812 3194
rect 514760 3130 514812 3136
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 514772 480 514800 3130
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 515968 480 515996 2994
rect 517164 480 517192 16546
rect 518348 3596 518400 3602
rect 518348 3538 518400 3544
rect 518360 480 518388 3538
rect 519556 480 519584 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 25638
rect 520936 3262 520964 47495
rect 520924 3256 520976 3262
rect 520924 3198 520976 3204
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 75142
rect 523144 6914 523172 78746
rect 525062 59936 525118 59945
rect 525062 59871 525118 59880
rect 523052 6886 523172 6914
rect 523052 480 523080 6886
rect 525076 3602 525104 59871
rect 525812 16574 525840 79290
rect 536840 78736 536892 78742
rect 536840 78678 536892 78684
rect 531320 70440 531372 70446
rect 531320 70382 531372 70388
rect 529940 64932 529992 64938
rect 529940 64874 529992 64880
rect 527824 38004 527876 38010
rect 527824 37946 527876 37952
rect 527180 24200 527232 24206
rect 527180 24142 527232 24148
rect 525812 16546 526208 16574
rect 525432 6180 525484 6186
rect 525432 6122 525484 6128
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 524236 3256 524288 3262
rect 524236 3198 524288 3204
rect 524248 480 524276 3198
rect 525444 480 525472 6122
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527192 6914 527220 24142
rect 527836 16574 527864 37946
rect 529204 18760 529256 18766
rect 529204 18702 529256 18708
rect 527836 16546 527956 16574
rect 527192 6886 527864 6914
rect 527836 480 527864 6886
rect 527928 4146 527956 16546
rect 527916 4140 527968 4146
rect 527916 4082 527968 4088
rect 529020 4140 529072 4146
rect 529020 4082 529072 4088
rect 529032 480 529060 4082
rect 529216 3534 529244 18702
rect 529204 3528 529256 3534
rect 529204 3470 529256 3476
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 529952 354 529980 64874
rect 531332 480 531360 70382
rect 534080 39364 534132 39370
rect 534080 39306 534132 39312
rect 531412 32428 531464 32434
rect 531412 32370 531464 32376
rect 531424 16574 531452 32370
rect 534092 16574 534120 39306
rect 535460 26920 535512 26926
rect 535460 26862 535512 26868
rect 535472 16574 535500 26862
rect 536852 16574 536880 78678
rect 549258 75168 549314 75177
rect 549258 75103 549314 75112
rect 543738 71088 543794 71097
rect 543738 71023 543794 71032
rect 539690 68232 539746 68241
rect 539690 68167 539746 68176
rect 538864 42084 538916 42090
rect 538864 42026 538916 42032
rect 538220 22840 538272 22846
rect 538220 22782 538272 22788
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3596 533764 3602
rect 533712 3538 533764 3544
rect 533724 480 533752 3538
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 22782
rect 538876 3602 538904 42026
rect 539704 16574 539732 68167
rect 542360 47592 542412 47598
rect 542360 47534 542412 47540
rect 542372 16574 542400 47534
rect 543752 16574 543780 71023
rect 547878 64152 547934 64161
rect 547878 64087 547934 64096
rect 545762 57216 545818 57225
rect 545762 57151 545818 57160
rect 539704 16546 540376 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 538864 3596 538916 3602
rect 538864 3538 538916 3544
rect 539600 3596 539652 3602
rect 539600 3538 539652 3544
rect 539612 480 539640 3538
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541992 4820 542044 4826
rect 541992 4762 542044 4768
rect 542004 480 542032 4762
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 7608 545540 7614
rect 545488 7550 545540 7556
rect 545500 480 545528 7550
rect 545776 3602 545804 57151
rect 546500 25628 546552 25634
rect 546500 25570 546552 25576
rect 545764 3596 545816 3602
rect 545764 3538 545816 3544
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 25570
rect 547892 480 547920 64087
rect 549272 16574 549300 75103
rect 561680 69080 561732 69086
rect 561680 69022 561732 69028
rect 557540 66292 557592 66298
rect 557540 66234 557592 66240
rect 556160 53100 556212 53106
rect 556160 53042 556212 53048
rect 553398 44976 553454 44985
rect 553398 44911 553454 44920
rect 552020 37936 552072 37942
rect 552020 37878 552072 37884
rect 552032 16574 552060 37878
rect 553412 16574 553440 44911
rect 554780 40724 554832 40730
rect 554780 40666 554832 40672
rect 549272 16546 550312 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 548616 11756 548668 11762
rect 548616 11698 548668 11704
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 11698
rect 550284 480 550312 16546
rect 551468 3596 551520 3602
rect 551468 3538 551520 3544
rect 551480 480 551508 3538
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 40666
rect 556172 16574 556200 53042
rect 557552 16574 557580 66234
rect 560944 55276 560996 55282
rect 560944 55218 560996 55224
rect 558920 36576 558972 36582
rect 558920 36518 558972 36524
rect 558932 16574 558960 36518
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 556160 8968 556212 8974
rect 556160 8910 556212 8916
rect 556172 480 556200 8910
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 560956 3534 560984 55218
rect 561692 16574 561720 69022
rect 574744 67652 574796 67658
rect 574744 67594 574796 67600
rect 567842 62792 567898 62801
rect 567842 62727 567898 62736
rect 563702 61432 563758 61441
rect 563702 61367 563758 61376
rect 561692 16546 562088 16574
rect 560852 3528 560904 3534
rect 560852 3470 560904 3476
rect 560944 3528 560996 3534
rect 560944 3470 560996 3476
rect 560864 480 560892 3470
rect 562060 480 562088 16546
rect 563060 10328 563112 10334
rect 563060 10270 563112 10276
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 10270
rect 563716 3058 563744 61367
rect 565818 44840 565874 44849
rect 565818 44775 565874 44784
rect 564532 24132 564584 24138
rect 564532 24074 564584 24080
rect 564544 6914 564572 24074
rect 565832 16574 565860 44775
rect 567200 18692 567252 18698
rect 567200 18634 567252 18640
rect 567212 16574 567240 18634
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 564452 6886 564572 6914
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 564452 480 564480 6886
rect 565636 3052 565688 3058
rect 565636 2994 565688 3000
rect 565648 480 565676 2994
rect 566844 480 566872 16546
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3534 567884 62727
rect 569958 50280 570014 50289
rect 569958 50215 570014 50224
rect 569972 16574 570000 50215
rect 571984 31068 572036 31074
rect 571984 31010 572036 31016
rect 571340 25560 571392 25566
rect 571340 25502 571392 25508
rect 569972 16546 570368 16574
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 569132 3528 569184 3534
rect 569132 3470 569184 3476
rect 569144 480 569172 3470
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 25502
rect 571996 3058 572024 31010
rect 574100 18624 574152 18630
rect 574100 18566 574152 18572
rect 574112 16574 574140 18566
rect 574112 16546 574692 16574
rect 572720 3596 572772 3602
rect 572720 3538 572772 3544
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 3538
rect 574664 3482 574692 16546
rect 574756 3602 574784 67594
rect 576136 6866 576164 139431
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580276 99521 580304 146367
rect 580368 143546 580396 152623
rect 580356 143540 580408 143546
rect 580356 143482 580408 143488
rect 580262 99512 580318 99521
rect 580262 99447 580318 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580262 79384 580318 79393
rect 580262 79319 580318 79328
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580276 59673 580304 79319
rect 581090 78568 581146 78577
rect 581090 78503 581146 78512
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 578240 51740 578292 51746
rect 578240 51682 578292 51688
rect 576216 35216 576268 35222
rect 576216 35158 576268 35164
rect 576124 6860 576176 6866
rect 576124 6802 576176 6808
rect 576228 4146 576256 35158
rect 578252 16574 578280 51682
rect 580264 22772 580316 22778
rect 580264 22714 580316 22720
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 578252 16546 578648 16574
rect 576216 4140 576268 4146
rect 576216 4082 576268 4088
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 576308 3596 576360 3602
rect 576308 3538 576360 3544
rect 574664 3454 575152 3482
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 3454
rect 576320 480 576348 3538
rect 577424 480 577452 4082
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 580276 3534 580304 22714
rect 581104 16574 581132 78503
rect 581104 16546 581776 16574
rect 580264 3528 580316 3534
rect 580264 3470 580316 3476
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581012 480 581040 3470
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 2778 371340 2834 371376
rect 2778 371320 2780 371340
rect 2780 371320 2832 371340
rect 2832 371320 2834 371340
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3054 267144 3110 267200
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 358420 3570 358456
rect 3514 358400 3516 358420
rect 3516 358400 3568 358420
rect 3568 358400 3570 358420
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 2778 214920 2834 214976
rect 3514 254088 3570 254144
rect 3514 241032 3570 241088
rect 3422 201864 3478 201920
rect 104806 201048 104862 201104
rect 3422 188808 3478 188864
rect 3422 162832 3478 162888
rect 3422 149776 3478 149832
rect 3146 110608 3202 110664
rect 3514 136720 3570 136776
rect 3514 84632 3570 84688
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 3422 45464 3478 45520
rect 3422 19352 3478 19408
rect 7562 75112 7618 75168
rect 3422 6432 3478 6488
rect 8942 68176 8998 68232
rect 11058 66816 11114 66872
rect 77298 81504 77354 81560
rect 14462 73752 14518 73808
rect 17222 36488 17278 36544
rect 22742 75248 22798 75304
rect 26238 73888 26294 73944
rect 25502 57160 25558 57216
rect 24858 33768 24914 33824
rect 27710 51720 27766 51776
rect 40038 66952 40094 67008
rect 39302 48864 39358 48920
rect 44178 47504 44234 47560
rect 49698 58520 49754 58576
rect 56598 46144 56654 46200
rect 93858 67088 93914 67144
rect 92478 64096 92534 64152
rect 100482 148280 100538 148336
rect 100666 193840 100722 193896
rect 100758 57840 100814 57896
rect 101678 57840 101734 57896
rect 100758 57160 100814 57216
rect 100758 52400 100814 52456
rect 101770 52400 101826 52456
rect 100758 51720 100814 51776
rect 100758 49544 100814 49600
rect 101954 49544 102010 49600
rect 100758 48864 100814 48920
rect 102138 67360 102194 67416
rect 102138 66952 102194 67008
rect 102138 53080 102194 53136
rect 100758 48184 100814 48240
rect 102046 48184 102102 48240
rect 100758 47504 100814 47560
rect 102230 46824 102286 46880
rect 102690 46824 102746 46880
rect 102230 46144 102286 46200
rect 103058 73888 103114 73944
rect 103242 192480 103298 192536
rect 103150 67360 103206 67416
rect 104438 196832 104494 196888
rect 104162 77152 104218 77208
rect 104622 194112 104678 194168
rect 107290 200368 107346 200424
rect 105542 71848 105598 71904
rect 104806 59200 104862 59256
rect 104070 58520 104126 58576
rect 104806 58520 104862 58576
rect 106186 192616 106242 192672
rect 106094 72664 106150 72720
rect 106094 71848 106150 71904
rect 107106 196560 107162 196616
rect 107382 200096 107438 200152
rect 107106 75656 107162 75712
rect 108210 196968 108266 197024
rect 108486 196696 108542 196752
rect 108486 75384 108542 75440
rect 107566 53760 107622 53816
rect 107566 53080 107622 53136
rect 108670 73752 108726 73808
rect 108946 199144 109002 199200
rect 109774 76608 109830 76664
rect 109866 71712 109922 71768
rect 108762 67088 108818 67144
rect 110142 67496 110198 67552
rect 110418 66952 110474 67008
rect 112442 195336 112498 195392
rect 111798 76880 111854 76936
rect 110878 64776 110934 64832
rect 110878 64096 110934 64152
rect 112350 76880 112406 76936
rect 112442 71168 112498 71224
rect 112810 75792 112866 75848
rect 113086 74432 113142 74488
rect 113454 146920 113510 146976
rect 114374 75520 114430 75576
rect 115202 192752 115258 192808
rect 114926 67088 114982 67144
rect 115754 77016 115810 77072
rect 116306 151000 116362 151056
rect 115846 72936 115902 72992
rect 116214 71576 116270 71632
rect 116398 79736 116454 79792
rect 116858 145696 116914 145752
rect 117962 261160 118018 261216
rect 117962 260888 118018 260944
rect 117686 195880 117742 195936
rect 117686 151136 117742 151192
rect 117134 74976 117190 75032
rect 118054 74024 118110 74080
rect 118882 138080 118938 138136
rect 119802 138896 119858 138952
rect 118514 72528 118570 72584
rect 119986 144744 120042 144800
rect 119894 76744 119950 76800
rect 120722 143384 120778 143440
rect 121182 259528 121238 259584
rect 121274 199688 121330 199744
rect 120538 80144 120594 80200
rect 120814 138760 120870 138816
rect 120722 73888 120778 73944
rect 129830 263200 129886 263256
rect 121734 143248 121790 143304
rect 122194 139032 122250 139088
rect 121918 71440 121974 71496
rect 121826 71304 121882 71360
rect 124862 260480 124918 260536
rect 127622 261160 127678 261216
rect 127622 260888 127678 260944
rect 133970 261024 134026 261080
rect 135902 265104 135958 265160
rect 137466 260888 137522 260944
rect 138754 264968 138810 265024
rect 138662 262928 138718 262984
rect 140318 262792 140374 262848
rect 142158 262384 142214 262440
rect 142250 260072 142306 260128
rect 142894 262384 142950 262440
rect 144182 262520 144238 262576
rect 143630 260208 143686 260264
rect 143400 260072 143456 260128
rect 144504 260208 144560 260264
rect 146206 263880 146262 263936
rect 145562 263744 145618 263800
rect 144918 259936 144974 259992
rect 146942 262656 146998 262712
rect 147678 260208 147734 260264
rect 148598 263608 148654 263664
rect 148368 260208 148424 260264
rect 148138 259664 148194 259720
rect 149058 260208 149114 260264
rect 150438 284280 150494 284336
rect 150530 263064 150586 263120
rect 150024 260208 150080 260264
rect 153382 275984 153438 276040
rect 156050 277480 156106 277536
rect 155958 260208 156014 260264
rect 156648 260208 156704 260264
rect 149242 259800 149298 259856
rect 158718 260888 158774 260944
rect 160834 265240 160890 265296
rect 160098 260208 160154 260264
rect 162214 265104 162270 265160
rect 162030 262656 162086 262712
rect 161064 260208 161120 260264
rect 161478 260208 161534 260264
rect 163410 263064 163466 263120
rect 163410 262384 163466 262440
rect 162720 260208 162776 260264
rect 162858 259936 162914 259992
rect 163594 263064 163650 263120
rect 164882 264968 164938 265024
rect 165158 264968 165214 265024
rect 164974 262520 165030 262576
rect 167550 265376 167606 265432
rect 161202 259800 161258 259856
rect 156878 259664 156934 259720
rect 123298 259528 123354 259584
rect 123942 259528 123998 259584
rect 155222 259528 155278 259584
rect 181350 260072 181406 260128
rect 181350 259664 181406 259720
rect 185674 259528 185730 259584
rect 122838 259392 122894 259448
rect 122562 209616 122618 209672
rect 122562 205536 122618 205592
rect 122562 201048 122618 201104
rect 124034 200640 124090 200696
rect 122378 140256 122434 140312
rect 122378 132504 122434 132560
rect 122378 132368 122434 132424
rect 122378 122848 122434 122904
rect 122378 122712 122434 122768
rect 122378 113192 122434 113248
rect 122378 113056 122434 113112
rect 122378 103536 122434 103592
rect 122378 103400 122434 103456
rect 122378 93880 122434 93936
rect 122378 93744 122434 93800
rect 122378 84224 122434 84280
rect 122378 84088 122434 84144
rect 122562 196016 122618 196072
rect 122562 190440 122618 190496
rect 122562 190304 122618 190360
rect 122562 180784 122618 180840
rect 122378 74568 122434 74624
rect 122838 148960 122894 149016
rect 124126 200504 124182 200560
rect 132038 200504 132094 200560
rect 126610 200368 126666 200424
rect 131946 200368 132002 200424
rect 124034 140936 124090 140992
rect 128910 200232 128966 200288
rect 126610 199416 126666 199472
rect 125230 148552 125286 148608
rect 125414 140800 125470 140856
rect 125230 140256 125286 140312
rect 125046 139848 125102 139904
rect 125598 141616 125654 141672
rect 128818 199552 128874 199608
rect 126978 146376 127034 146432
rect 126794 143384 126850 143440
rect 126794 142160 126850 142216
rect 126702 140256 126758 140312
rect 127346 141072 127402 141128
rect 130198 200096 130254 200152
rect 129646 199008 129702 199064
rect 129186 197240 129242 197296
rect 128910 140120 128966 140176
rect 129186 139984 129242 140040
rect 130198 198872 130254 198928
rect 131578 200096 131634 200152
rect 131946 199960 132002 200016
rect 131486 198736 131542 198792
rect 130474 197104 130530 197160
rect 130290 146240 130346 146296
rect 129830 146104 129886 146160
rect 129922 145968 129978 146024
rect 132038 195200 132094 195256
rect 131118 145832 131174 145888
rect 132820 199824 132876 199880
rect 133372 199824 133428 199880
rect 132774 197376 132830 197432
rect 133142 199280 133198 199336
rect 133142 199028 133198 199064
rect 133142 199008 133144 199028
rect 133144 199008 133196 199028
rect 133196 199008 133198 199028
rect 133050 194112 133106 194168
rect 132314 188400 132370 188456
rect 133602 198464 133658 198520
rect 134292 199824 134348 199880
rect 134844 199824 134900 199880
rect 134614 196832 134670 196888
rect 135580 199824 135636 199880
rect 135166 197376 135222 197432
rect 135350 199416 135406 199472
rect 133970 189080 134026 189136
rect 136224 199824 136280 199880
rect 136776 199858 136832 199914
rect 135994 196152 136050 196208
rect 136178 198872 136234 198928
rect 136178 196288 136234 196344
rect 136270 196016 136326 196072
rect 135626 188400 135682 188456
rect 136546 199416 136602 199472
rect 137144 199824 137200 199880
rect 137512 199824 137568 199880
rect 136638 199144 136694 199200
rect 136454 194928 136510 194984
rect 136914 199144 136970 199200
rect 136822 198872 136878 198928
rect 136730 192480 136786 192536
rect 137374 199416 137430 199472
rect 137190 194928 137246 194984
rect 137006 188400 137062 188456
rect 135442 187040 135498 187096
rect 137282 192616 137338 192672
rect 137282 187992 137338 188048
rect 137190 187584 137246 187640
rect 133050 148280 133106 148336
rect 137880 199858 137936 199914
rect 138156 199824 138212 199880
rect 137926 199008 137982 199064
rect 137834 196968 137890 197024
rect 138202 199416 138258 199472
rect 138018 195880 138074 195936
rect 137650 188400 137706 188456
rect 137466 186224 137522 186280
rect 138202 196560 138258 196616
rect 138478 196696 138534 196752
rect 138386 194928 138442 194984
rect 138662 198736 138718 198792
rect 138570 194792 138626 194848
rect 138846 199416 138902 199472
rect 139306 199280 139362 199336
rect 139214 199008 139270 199064
rect 139214 198328 139270 198384
rect 139214 197648 139270 197704
rect 139214 196016 139270 196072
rect 139122 194928 139178 194984
rect 138938 188536 138994 188592
rect 138846 188400 138902 188456
rect 139674 199144 139730 199200
rect 140042 199008 140098 199064
rect 140042 197376 140098 197432
rect 140318 199280 140374 199336
rect 140318 199144 140374 199200
rect 140226 199008 140282 199064
rect 140226 198872 140282 198928
rect 139766 188536 139822 188592
rect 140594 199280 140650 199336
rect 140410 188400 140466 188456
rect 140870 144608 140926 144664
rect 138662 143928 138718 143984
rect 139398 143792 139454 143848
rect 142112 199858 142168 199914
rect 142480 199858 142536 199914
rect 142066 191120 142122 191176
rect 142434 199552 142490 199608
rect 142342 195336 142398 195392
rect 142250 192752 142306 192808
rect 142158 190984 142214 191040
rect 141698 190304 141754 190360
rect 142066 180784 142122 180840
rect 142066 180648 142122 180704
rect 141422 141480 141478 141536
rect 142066 171128 142122 171184
rect 142066 170992 142122 171048
rect 142066 161472 142122 161528
rect 142066 161336 142122 161392
rect 142066 151816 142122 151872
rect 142066 151680 142122 151736
rect 143492 199858 143548 199914
rect 144136 199858 144192 199914
rect 144320 199858 144376 199914
rect 144504 199858 144560 199914
rect 143906 195064 143962 195120
rect 144182 199552 144238 199608
rect 144550 199688 144606 199744
rect 144872 199824 144928 199880
rect 144458 188264 144514 188320
rect 145516 199858 145572 199914
rect 145470 199688 145526 199744
rect 145884 199824 145940 199880
rect 145378 198192 145434 198248
rect 145286 197648 145342 197704
rect 145746 199416 145802 199472
rect 145470 193976 145526 194032
rect 144642 183776 144698 183832
rect 142526 144472 142582 144528
rect 142066 142296 142122 142352
rect 141606 141208 141662 141264
rect 144182 144336 144238 144392
rect 143078 143248 143134 143304
rect 143630 141616 143686 141672
rect 145010 142976 145066 143032
rect 146206 199008 146262 199064
rect 146114 191120 146170 191176
rect 146482 197920 146538 197976
rect 146574 197512 146630 197568
rect 146942 195608 146998 195664
rect 147218 191120 147274 191176
rect 145746 148552 145802 148608
rect 147586 199688 147642 199744
rect 148000 199858 148056 199914
rect 148644 199858 148700 199914
rect 147770 197648 147826 197704
rect 146298 145696 146354 145752
rect 145838 144200 145894 144256
rect 146390 143112 146446 143168
rect 147586 146920 147642 146976
rect 148046 195472 148102 195528
rect 149656 199824 149712 199880
rect 148874 198736 148930 198792
rect 149058 196016 149114 196072
rect 147678 145560 147734 145616
rect 148046 142840 148102 142896
rect 149334 198736 149390 198792
rect 150024 199824 150080 199880
rect 150484 199858 150540 199914
rect 150070 199724 150072 199744
rect 150072 199724 150124 199744
rect 150124 199724 150126 199744
rect 149242 195744 149298 195800
rect 149702 195472 149758 195528
rect 150070 199688 150126 199724
rect 149978 195472 150034 195528
rect 149978 188400 150034 188456
rect 151128 199824 151184 199880
rect 151496 199858 151552 199914
rect 150806 199552 150862 199608
rect 150714 195200 150770 195256
rect 150346 195064 150402 195120
rect 150346 191120 150402 191176
rect 150346 149640 150402 149696
rect 149702 142704 149758 142760
rect 150438 141344 150494 141400
rect 152324 199824 152380 199880
rect 151542 195880 151598 195936
rect 152094 199552 152150 199608
rect 152600 199824 152656 199880
rect 152278 194112 152334 194168
rect 152094 191528 152150 191584
rect 152462 199144 152518 199200
rect 151082 144064 151138 144120
rect 153980 199824 154036 199880
rect 154348 199858 154404 199914
rect 152554 188808 152610 188864
rect 152738 187312 152794 187368
rect 153290 197240 153346 197296
rect 153566 197240 153622 197296
rect 154026 199552 154082 199608
rect 153750 199280 153806 199336
rect 153658 195200 153714 195256
rect 153382 148416 153438 148472
rect 153290 145560 153346 145616
rect 154808 199858 154864 199914
rect 155268 199858 155324 199914
rect 154394 195472 154450 195528
rect 154302 195200 154358 195256
rect 154670 199416 154726 199472
rect 154670 197104 154726 197160
rect 155314 199688 155370 199744
rect 155498 199688 155554 199744
rect 156004 199824 156060 199880
rect 156372 199824 156428 199880
rect 156832 199858 156888 199914
rect 155774 199688 155830 199744
rect 154946 189896 155002 189952
rect 155682 199416 155738 199472
rect 154946 149776 155002 149832
rect 154762 147192 154818 147248
rect 154486 144336 154542 144392
rect 155130 142840 155186 142896
rect 156326 199688 156382 199744
rect 155958 198736 156014 198792
rect 156142 198736 156198 198792
rect 155866 195880 155922 195936
rect 156878 199280 156934 199336
rect 156786 198328 156842 198384
rect 156602 197376 156658 197432
rect 157154 199416 157210 199472
rect 157154 199300 157210 199336
rect 157154 199280 157156 199300
rect 157156 199280 157208 199300
rect 157208 199280 157210 199300
rect 157752 199824 157808 199880
rect 157430 198056 157486 198112
rect 156050 147328 156106 147384
rect 156970 142704 157026 142760
rect 157614 150320 157670 150376
rect 157430 150184 157486 150240
rect 157246 149912 157302 149968
rect 158304 199858 158360 199914
rect 158258 199688 158314 199744
rect 159040 199824 159096 199880
rect 157982 193976 158038 194032
rect 158534 191120 158590 191176
rect 157798 149504 157854 149560
rect 158994 198464 159050 198520
rect 158902 189216 158958 189272
rect 159086 190984 159142 191040
rect 159684 199824 159740 199880
rect 159362 199416 159418 199472
rect 159362 184048 159418 184104
rect 160098 199688 160154 199744
rect 160374 199688 160430 199744
rect 160282 195880 160338 195936
rect 160190 191256 160246 191312
rect 160650 194928 160706 194984
rect 160466 191392 160522 191448
rect 158074 144064 158130 144120
rect 157338 142024 157394 142080
rect 157154 141344 157210 141400
rect 157062 140120 157118 140176
rect 159454 144200 159510 144256
rect 158534 139984 158590 140040
rect 161064 199824 161120 199880
rect 160742 191120 160798 191176
rect 161202 199436 161258 199472
rect 161202 199416 161204 199436
rect 161204 199416 161256 199436
rect 161256 199416 161258 199436
rect 161386 190984 161442 191040
rect 161846 195064 161902 195120
rect 160650 145696 160706 145752
rect 160006 142976 160062 143032
rect 161938 187040 161994 187096
rect 162306 198328 162362 198384
rect 163088 199824 163144 199880
rect 163042 199688 163098 199744
rect 162674 191120 162730 191176
rect 162950 199416 163006 199472
rect 163042 195880 163098 195936
rect 162950 195336 163006 195392
rect 163272 199688 163328 199744
rect 163226 199416 163282 199472
rect 162490 187448 162546 187504
rect 162306 145832 162362 145888
rect 162214 144472 162270 144528
rect 161938 143112 161994 143168
rect 163732 199824 163788 199880
rect 163594 198192 163650 198248
rect 164008 199824 164064 199880
rect 163962 199688 164018 199744
rect 164376 199824 164432 199880
rect 164836 199824 164892 199880
rect 165204 199824 165260 199880
rect 165848 199858 165904 199914
rect 164054 195200 164110 195256
rect 164974 196560 165030 196616
rect 163870 187312 163926 187368
rect 163594 143248 163650 143304
rect 164146 141480 164202 141536
rect 164698 195200 164754 195256
rect 164514 194928 164570 194984
rect 164974 188536 165030 188592
rect 165618 199688 165674 199744
rect 165434 185816 165490 185872
rect 165250 182552 165306 182608
rect 164422 145968 164478 146024
rect 165250 143384 165306 143440
rect 166400 199858 166456 199914
rect 166354 199688 166410 199744
rect 166676 199858 166732 199914
rect 166952 199824 167008 199880
rect 166538 197240 166594 197296
rect 166814 199708 166870 199744
rect 166814 199688 166816 199708
rect 166816 199688 166868 199708
rect 166868 199688 166870 199708
rect 167090 199688 167146 199744
rect 167090 198056 167146 198112
rect 167090 197648 167146 197704
rect 166906 191120 166962 191176
rect 165986 190032 166042 190088
rect 165894 152496 165950 152552
rect 167366 195472 167422 195528
rect 168240 199824 168296 199880
rect 167642 198600 167698 198656
rect 167918 195336 167974 195392
rect 168608 199824 168664 199880
rect 168378 195472 168434 195528
rect 168286 152360 168342 152416
rect 169068 199858 169124 199914
rect 169528 199824 169584 199880
rect 169988 199824 170044 199880
rect 168746 195336 168802 195392
rect 169574 199416 169630 199472
rect 169758 199452 169760 199472
rect 169760 199452 169812 199472
rect 169812 199452 169814 199472
rect 169758 199416 169814 199452
rect 169666 198464 169722 198520
rect 169758 198056 169814 198112
rect 169574 196696 169630 196752
rect 169850 196968 169906 197024
rect 169298 191120 169354 191176
rect 168746 185816 168802 185872
rect 170126 199416 170182 199472
rect 170448 199824 170504 199880
rect 171000 199824 171056 199880
rect 168470 154400 168526 154456
rect 168010 144744 168066 144800
rect 166354 144608 166410 144664
rect 165526 143928 165582 143984
rect 169758 140392 169814 140448
rect 170402 199416 170458 199472
rect 170402 189216 170458 189272
rect 170770 199688 170826 199744
rect 170770 199452 170772 199472
rect 170772 199452 170824 199472
rect 170824 199452 170826 199472
rect 170770 199416 170826 199452
rect 170862 198328 170918 198384
rect 170678 195472 170734 195528
rect 171368 199858 171424 199914
rect 171046 199724 171048 199744
rect 171048 199724 171100 199744
rect 171100 199724 171102 199744
rect 171046 199688 171102 199724
rect 171644 199824 171700 199880
rect 171506 198600 171562 198656
rect 169942 140256 169998 140312
rect 172288 199824 172344 199880
rect 172334 199688 172390 199744
rect 171874 198056 171930 198112
rect 171782 196832 171838 196888
rect 172242 199416 172298 199472
rect 172426 199416 172482 199472
rect 172058 191120 172114 191176
rect 172794 199416 172850 199472
rect 173760 199824 173816 199880
rect 173162 191256 173218 191312
rect 172978 191120 173034 191176
rect 174312 199858 174368 199914
rect 173806 199436 173862 199472
rect 173806 199416 173808 199436
rect 173808 199416 173860 199436
rect 173860 199416 173862 199436
rect 175140 199824 175196 199880
rect 173714 190984 173770 191040
rect 172610 147056 172666 147112
rect 174266 150048 174322 150104
rect 174634 196424 174690 196480
rect 174910 198056 174966 198112
rect 175416 199824 175472 199880
rect 175462 199688 175518 199744
rect 175002 195472 175058 195528
rect 175278 195608 175334 195664
rect 175462 192480 175518 192536
rect 175876 199824 175932 199880
rect 176336 199824 176392 199880
rect 175922 199724 175924 199744
rect 175924 199724 175976 199744
rect 175976 199724 175978 199744
rect 175922 199688 175978 199724
rect 175646 194792 175702 194848
rect 175462 187720 175518 187776
rect 176290 199688 176346 199744
rect 176888 199824 176944 199880
rect 177072 199824 177128 199880
rect 176290 196968 176346 197024
rect 176474 191120 176530 191176
rect 176198 188400 176254 188456
rect 176750 198056 176806 198112
rect 176750 197512 176806 197568
rect 176658 187992 176714 188048
rect 174082 146240 174138 146296
rect 173898 146104 173954 146160
rect 176658 141616 176714 141672
rect 177486 188400 177542 188456
rect 178222 200368 178278 200424
rect 178866 200096 178922 200152
rect 177302 188264 177358 188320
rect 178314 195064 178370 195120
rect 176750 141208 176806 141264
rect 179050 140120 179106 140176
rect 124494 139304 124550 139360
rect 125506 139304 125562 139360
rect 125966 139304 126022 139360
rect 126150 139304 126206 139360
rect 127622 139304 127678 139360
rect 130014 139304 130070 139360
rect 131026 139304 131082 139360
rect 132222 139304 132278 139360
rect 149610 139304 149666 139360
rect 150990 139304 151046 139360
rect 155222 139304 155278 139360
rect 155774 139304 155830 139360
rect 159546 139304 159602 139360
rect 159822 139304 159878 139360
rect 165342 139304 165398 139360
rect 178866 139304 178922 139360
rect 181442 198212 181498 198248
rect 181442 198192 181444 198212
rect 181444 198192 181496 198212
rect 181496 198192 181498 198212
rect 180154 139712 180210 139768
rect 183006 197104 183062 197160
rect 182270 140528 182326 140584
rect 181626 139984 181682 140040
rect 183466 139984 183522 140040
rect 186410 194792 186466 194848
rect 184018 139576 184074 139632
rect 184662 139576 184718 139632
rect 183834 139440 183890 139496
rect 184386 139440 184442 139496
rect 180154 139304 180210 139360
rect 184570 139440 184626 139496
rect 185858 140120 185914 140176
rect 186226 140120 186282 140176
rect 186226 139712 186282 139768
rect 177762 80688 177818 80744
rect 131854 80416 131910 80472
rect 124126 80280 124182 80336
rect 124034 78376 124090 78432
rect 124034 74296 124090 74352
rect 124126 72800 124182 72856
rect 130842 79464 130898 79520
rect 177946 80708 178002 80744
rect 177946 80688 177948 80708
rect 177948 80688 178000 80708
rect 178000 80688 178002 80708
rect 178406 80688 178462 80744
rect 132130 80416 132186 80472
rect 131762 79872 131818 79928
rect 131026 78648 131082 78704
rect 131118 76608 131174 76664
rect 131578 76608 131634 76664
rect 132222 79600 132278 79656
rect 132222 79464 132278 79520
rect 132222 78648 132278 78704
rect 132038 78512 132094 78568
rect 132820 79906 132876 79962
rect 133188 79906 133244 79962
rect 133556 79906 133612 79962
rect 133924 79872 133980 79928
rect 134292 79872 134348 79928
rect 133326 79620 133382 79656
rect 133326 79600 133328 79620
rect 133328 79600 133380 79620
rect 133380 79600 133382 79620
rect 133234 73752 133290 73808
rect 133602 79464 133658 79520
rect 133970 78512 134026 78568
rect 134246 79600 134302 79656
rect 134062 77696 134118 77752
rect 135212 79872 135268 79928
rect 134062 74160 134118 74216
rect 135166 79600 135222 79656
rect 135166 77696 135222 77752
rect 135074 75928 135130 75984
rect 136500 79872 136556 79928
rect 136776 79872 136832 79928
rect 137144 79906 137200 79962
rect 137328 79872 137384 79928
rect 135718 79600 135774 79656
rect 135534 79484 135590 79520
rect 135534 79464 135536 79484
rect 135536 79464 135588 79484
rect 135588 79464 135590 79484
rect 135442 77696 135498 77752
rect 135718 79484 135774 79520
rect 135718 79464 135720 79484
rect 135720 79464 135772 79484
rect 135772 79464 135774 79484
rect 135350 77560 135406 77616
rect 135350 76628 135406 76664
rect 135350 76608 135352 76628
rect 135352 76608 135404 76628
rect 135404 76608 135406 76628
rect 135902 79600 135958 79656
rect 135810 77424 135866 77480
rect 135994 78512 136050 78568
rect 136730 79600 136786 79656
rect 137006 79620 137062 79656
rect 137006 79600 137008 79620
rect 137008 79600 137060 79620
rect 137060 79600 137062 79620
rect 137006 79484 137062 79520
rect 137006 79464 137008 79484
rect 137008 79464 137060 79484
rect 137060 79464 137062 79484
rect 137374 79600 137430 79656
rect 137972 79872 138028 79928
rect 137650 79464 137706 79520
rect 138432 79906 138488 79962
rect 137834 77968 137890 78024
rect 138202 77832 138258 77888
rect 138110 77696 138166 77752
rect 138018 77152 138074 77208
rect 138524 79736 138580 79792
rect 138478 79636 138480 79656
rect 138480 79636 138532 79656
rect 138532 79636 138534 79656
rect 138478 79600 138534 79636
rect 138708 79906 138764 79962
rect 139260 79872 139316 79928
rect 139214 79600 139270 79656
rect 138662 78376 138718 78432
rect 138754 77832 138810 77888
rect 138754 77288 138810 77344
rect 139536 79736 139592 79792
rect 140088 79872 140144 79928
rect 139490 77696 139546 77752
rect 139582 77560 139638 77616
rect 140134 79736 140190 79792
rect 140364 79906 140420 79962
rect 140548 79906 140604 79962
rect 140042 79328 140098 79384
rect 140226 79600 140282 79656
rect 140594 79772 140596 79792
rect 140596 79772 140648 79792
rect 140648 79772 140650 79792
rect 140594 79736 140650 79772
rect 140502 79600 140558 79656
rect 140870 79328 140926 79384
rect 140778 78512 140834 78568
rect 142020 79872 142076 79928
rect 141744 79736 141800 79792
rect 141054 77696 141110 77752
rect 140962 77560 141018 77616
rect 141330 79328 141386 79384
rect 141238 76880 141294 76936
rect 141606 79364 141608 79384
rect 141608 79364 141660 79384
rect 141660 79364 141662 79384
rect 141606 79328 141662 79364
rect 142664 79906 142720 79962
rect 143032 79906 143088 79962
rect 142848 79736 142904 79792
rect 143768 79872 143824 79928
rect 142710 79600 142766 79656
rect 142066 70352 142122 70408
rect 142066 66952 142122 67008
rect 143170 79600 143226 79656
rect 143630 79736 143686 79792
rect 142710 75928 142766 75984
rect 142894 76608 142950 76664
rect 143170 75928 143226 75984
rect 143538 78648 143594 78704
rect 143814 79636 143816 79656
rect 143816 79636 143868 79656
rect 143868 79636 143870 79656
rect 143814 79600 143870 79636
rect 144504 79872 144560 79928
rect 144688 79872 144744 79928
rect 144412 79736 144468 79792
rect 144550 78512 144606 78568
rect 144642 74432 144698 74488
rect 145148 79872 145204 79928
rect 144826 79328 144882 79384
rect 145332 79736 145388 79792
rect 146160 79906 146216 79962
rect 145378 79600 145434 79656
rect 145286 79328 145342 79384
rect 145654 77288 145710 77344
rect 145746 76744 145802 76800
rect 146206 79736 146262 79792
rect 146206 79192 146262 79248
rect 146620 79838 146676 79894
rect 146022 76200 146078 76256
rect 146390 78512 146446 78568
rect 146896 79872 146952 79928
rect 147356 79906 147412 79962
rect 147632 79872 147688 79928
rect 147402 79736 147458 79792
rect 148000 79872 148056 79928
rect 148184 79838 148240 79894
rect 146758 79328 146814 79384
rect 146850 76608 146906 76664
rect 147862 79636 147864 79656
rect 147864 79636 147916 79656
rect 147916 79636 147918 79656
rect 147862 79600 147918 79636
rect 147494 79328 147550 79384
rect 146758 71712 146814 71768
rect 147218 79192 147274 79248
rect 147402 79192 147458 79248
rect 147310 78648 147366 78704
rect 148138 79600 148194 79656
rect 148046 79328 148102 79384
rect 148644 79872 148700 79928
rect 148506 77968 148562 78024
rect 148690 79328 148746 79384
rect 148690 79192 148746 79248
rect 148874 79772 148876 79792
rect 148876 79772 148928 79792
rect 148928 79772 148930 79792
rect 148874 79736 148930 79772
rect 148966 79192 149022 79248
rect 148598 77832 148654 77888
rect 149380 79906 149436 79962
rect 149426 79736 149482 79792
rect 150024 79906 150080 79962
rect 150208 79872 150264 79928
rect 150392 79906 150448 79962
rect 150576 79872 150632 79928
rect 149426 79192 149482 79248
rect 149334 76200 149390 76256
rect 149518 78104 149574 78160
rect 149610 76336 149666 76392
rect 149794 79600 149850 79656
rect 150070 79600 150126 79656
rect 150254 79464 150310 79520
rect 150438 79464 150494 79520
rect 150346 79192 150402 79248
rect 150622 79736 150678 79792
rect 150852 79906 150908 79962
rect 150898 79736 150954 79792
rect 151128 79872 151184 79928
rect 151312 79906 151368 79962
rect 150530 78376 150586 78432
rect 150530 77288 150586 77344
rect 151082 79328 151138 79384
rect 150990 77288 151046 77344
rect 151266 79736 151322 79792
rect 151358 79464 151414 79520
rect 151772 79872 151828 79928
rect 151680 79736 151736 79792
rect 151450 78512 151506 78568
rect 151726 79600 151782 79656
rect 151910 79056 151966 79112
rect 152232 79772 152234 79792
rect 152234 79772 152286 79792
rect 152286 79772 152288 79792
rect 152232 79736 152288 79772
rect 152600 79906 152656 79962
rect 152784 79838 152840 79894
rect 152462 79600 152518 79656
rect 152370 75928 152426 75984
rect 152922 79600 152978 79656
rect 152830 74568 152886 74624
rect 153612 79872 153668 79928
rect 153106 79464 153162 79520
rect 153014 79056 153070 79112
rect 153290 76744 153346 76800
rect 153474 79500 153476 79520
rect 153476 79500 153528 79520
rect 153528 79500 153530 79520
rect 153474 79464 153530 79500
rect 153382 74432 153438 74488
rect 153474 73072 153530 73128
rect 152462 63008 152518 63064
rect 153842 79600 153898 79656
rect 153934 79464 153990 79520
rect 154026 76608 154082 76664
rect 153566 69944 153622 70000
rect 154302 79736 154358 79792
rect 154210 78648 154266 78704
rect 154302 78104 154358 78160
rect 154210 73072 154266 73128
rect 154118 69944 154174 70000
rect 154716 79906 154772 79962
rect 155084 79906 155140 79962
rect 154900 79770 154956 79826
rect 155130 79736 155186 79792
rect 155268 79736 155324 79792
rect 155636 79872 155692 79928
rect 154486 79600 154542 79656
rect 154578 79464 154634 79520
rect 154394 77832 154450 77888
rect 154854 79600 154910 79656
rect 154762 79192 154818 79248
rect 155820 79872 155876 79928
rect 156096 79906 156152 79962
rect 156464 79906 156520 79962
rect 155590 79600 155646 79656
rect 155590 79328 155646 79384
rect 155866 79600 155922 79656
rect 155774 79192 155830 79248
rect 155682 74160 155738 74216
rect 156142 78920 156198 78976
rect 157016 79736 157072 79792
rect 157200 79872 157256 79928
rect 156602 79636 156604 79656
rect 156604 79636 156656 79656
rect 156656 79636 156658 79656
rect 156602 79600 156658 79636
rect 156510 79464 156566 79520
rect 156418 79056 156474 79112
rect 156970 79192 157026 79248
rect 156970 79056 157026 79112
rect 156878 78784 156934 78840
rect 156786 75792 156842 75848
rect 156878 75520 156934 75576
rect 156786 74024 156842 74080
rect 156602 70080 156658 70136
rect 157844 79872 157900 79928
rect 158580 79872 158636 79928
rect 158304 79736 158360 79792
rect 157522 79636 157524 79656
rect 157524 79636 157576 79656
rect 157576 79636 157578 79656
rect 157154 74976 157210 75032
rect 157522 79600 157578 79636
rect 157430 79464 157486 79520
rect 157614 79464 157670 79520
rect 157706 78784 157762 78840
rect 157982 79464 158038 79520
rect 158166 79600 158222 79656
rect 157890 79056 157946 79112
rect 158166 79328 158222 79384
rect 158074 78920 158130 78976
rect 158074 74296 158130 74352
rect 157982 72800 158038 72856
rect 157338 21256 157394 21312
rect 158442 79620 158498 79656
rect 158626 79636 158628 79656
rect 158628 79636 158680 79656
rect 158680 79636 158682 79656
rect 158442 79600 158444 79620
rect 158444 79600 158496 79620
rect 158496 79600 158498 79620
rect 158626 79600 158682 79636
rect 158718 79464 158774 79520
rect 158534 78512 158590 78568
rect 158534 78104 158590 78160
rect 158350 74296 158406 74352
rect 158350 73908 158406 73944
rect 158350 73888 158352 73908
rect 158352 73888 158404 73908
rect 158404 73888 158406 73908
rect 158442 72392 158498 72448
rect 158902 78920 158958 78976
rect 159776 79872 159832 79928
rect 159408 79736 159464 79792
rect 160512 79872 160568 79928
rect 159960 79736 160016 79792
rect 160190 79736 160246 79792
rect 159546 78412 159548 78432
rect 159548 78412 159600 78432
rect 159600 78412 159602 78432
rect 159546 78376 159602 78412
rect 159822 79500 159824 79520
rect 159824 79500 159876 79520
rect 159876 79500 159878 79520
rect 159822 79464 159878 79500
rect 159822 72936 159878 72992
rect 160006 75928 160062 75984
rect 160466 79736 160522 79792
rect 160788 79906 160844 79962
rect 161248 79906 161304 79962
rect 161064 79736 161120 79792
rect 160466 78240 160522 78296
rect 160374 75656 160430 75712
rect 160650 79600 160706 79656
rect 160742 79464 160798 79520
rect 160834 75928 160890 75984
rect 161110 79464 161166 79520
rect 160098 30912 160154 30968
rect 161432 79736 161488 79792
rect 161616 79872 161672 79928
rect 161202 78512 161258 78568
rect 161202 78240 161258 78296
rect 161386 79600 161442 79656
rect 161754 79600 161810 79656
rect 161984 79736 162040 79792
rect 162720 79906 162776 79962
rect 163088 79872 163144 79928
rect 163548 79872 163604 79928
rect 162214 79600 162270 79656
rect 162490 79600 162546 79656
rect 162398 79464 162454 79520
rect 162122 73072 162178 73128
rect 162122 72392 162178 72448
rect 162582 79328 162638 79384
rect 162490 77016 162546 77072
rect 162490 76880 162546 76936
rect 161294 8880 161350 8936
rect 162950 77696 163006 77752
rect 162858 77560 162914 77616
rect 162674 76880 162730 76936
rect 163318 79736 163374 79792
rect 163134 78920 163190 78976
rect 163916 79736 163972 79792
rect 163502 79484 163558 79520
rect 163502 79464 163504 79484
rect 163504 79464 163556 79484
rect 163556 79464 163558 79484
rect 163594 73616 163650 73672
rect 164192 79872 164248 79928
rect 163778 78512 163834 78568
rect 164054 79500 164056 79520
rect 164056 79500 164108 79520
rect 164108 79500 164110 79520
rect 164054 79464 164110 79500
rect 164146 77152 164202 77208
rect 164744 79736 164800 79792
rect 164928 79872 164984 79928
rect 165480 79872 165536 79928
rect 164606 79328 164662 79384
rect 164790 78104 164846 78160
rect 164974 78376 165030 78432
rect 165158 79192 165214 79248
rect 165250 78784 165306 78840
rect 165342 78376 165398 78432
rect 165250 77968 165306 78024
rect 165848 79872 165904 79928
rect 165434 73616 165490 73672
rect 166078 79736 166134 79792
rect 166584 79872 166640 79928
rect 166308 79736 166364 79792
rect 166952 79906 167008 79962
rect 166538 79192 166594 79248
rect 166446 77968 166502 78024
rect 166630 78784 166686 78840
rect 166906 75928 166962 75984
rect 167182 79328 167238 79384
rect 167182 76472 167238 76528
rect 167688 79872 167744 79928
rect 167458 79328 167514 79384
rect 167274 75656 167330 75712
rect 167734 79600 167790 79656
rect 167826 76064 167882 76120
rect 168148 79906 168204 79962
rect 168424 79872 168480 79928
rect 168010 75792 168066 75848
rect 168194 79600 168250 79656
rect 168194 79328 168250 79384
rect 168286 79192 168342 79248
rect 168470 79736 168526 79792
rect 168700 79906 168756 79962
rect 168378 75928 168434 75984
rect 169022 79620 169078 79656
rect 169022 79600 169024 79620
rect 169024 79600 169076 79620
rect 169076 79600 169078 79620
rect 169436 79872 169492 79928
rect 169804 79906 169860 79962
rect 169574 79736 169630 79792
rect 169390 79636 169392 79656
rect 169392 79636 169444 79656
rect 169444 79636 169446 79656
rect 169390 79600 169446 79636
rect 169390 79328 169446 79384
rect 169666 79600 169722 79656
rect 170080 79906 170136 79962
rect 170448 79872 170504 79928
rect 170126 79756 170182 79792
rect 170126 79736 170128 79756
rect 170128 79736 170180 79756
rect 170180 79736 170182 79756
rect 171000 79736 171056 79792
rect 171368 79872 171424 79928
rect 171552 79872 171608 79928
rect 169758 79056 169814 79112
rect 169942 79192 169998 79248
rect 169850 76472 169906 76528
rect 170402 79600 170458 79656
rect 170586 79328 170642 79384
rect 170494 78920 170550 78976
rect 170954 79192 171010 79248
rect 170770 76064 170826 76120
rect 171322 79600 171378 79656
rect 171322 78784 171378 78840
rect 171230 75928 171286 75984
rect 171138 71168 171194 71224
rect 172012 79736 172068 79792
rect 172380 79872 172436 79928
rect 171782 79620 171838 79656
rect 171782 79600 171784 79620
rect 171784 79600 171836 79620
rect 171836 79600 171838 79620
rect 171966 79192 172022 79248
rect 171690 79056 171746 79112
rect 171506 78648 171562 78704
rect 171966 78648 172022 78704
rect 172242 79328 172298 79384
rect 172058 75928 172114 75984
rect 172150 70216 172206 70272
rect 172334 77968 172390 78024
rect 172748 79906 172804 79962
rect 173760 79906 173816 79962
rect 173484 79736 173540 79792
rect 172610 79600 172666 79656
rect 172426 74296 172482 74352
rect 172426 73752 172482 73808
rect 172702 75792 172758 75848
rect 172978 79328 173034 79384
rect 173254 79328 173310 79384
rect 173070 75112 173126 75168
rect 173346 76608 173402 76664
rect 174128 79838 174184 79894
rect 174496 79906 174552 79962
rect 174680 79906 174736 79962
rect 174864 79872 174920 79928
rect 173898 79328 173954 79384
rect 173714 75384 173770 75440
rect 174082 79620 174138 79656
rect 174082 79600 174084 79620
rect 174084 79600 174136 79620
rect 174136 79600 174138 79620
rect 174082 76608 174138 76664
rect 174358 79600 174414 79656
rect 173990 75248 174046 75304
rect 174358 78648 174414 78704
rect 174542 79328 174598 79384
rect 175140 79872 175196 79928
rect 175094 79736 175150 79792
rect 174910 79600 174966 79656
rect 174450 68720 174506 68776
rect 174726 75248 174782 75304
rect 175186 79192 175242 79248
rect 175186 77016 175242 77072
rect 175186 76744 175242 76800
rect 175094 74296 175150 74352
rect 175968 79960 176024 79962
rect 175968 79908 175970 79960
rect 175970 79908 176022 79960
rect 176022 79908 176024 79960
rect 175968 79906 176024 79908
rect 176152 79872 176208 79928
rect 176014 79772 176016 79792
rect 176016 79772 176068 79792
rect 176068 79772 176070 79792
rect 176014 79736 176070 79772
rect 176198 79736 176254 79792
rect 176336 79736 176392 79792
rect 175646 79328 175702 79384
rect 175554 75656 175610 75712
rect 175462 75112 175518 75168
rect 175922 79328 175978 79384
rect 175830 77560 175886 77616
rect 175830 77288 175886 77344
rect 176106 79600 176162 79656
rect 176382 79620 176438 79656
rect 176382 79600 176384 79620
rect 176384 79600 176436 79620
rect 176436 79600 176438 79620
rect 176198 78784 176254 78840
rect 176198 77560 176254 77616
rect 176658 79600 176714 79656
rect 176566 77152 176622 77208
rect 176474 77016 176530 77072
rect 176566 75656 176622 75712
rect 175922 18536 175978 18592
rect 171966 3304 172022 3360
rect 176750 79192 176806 79248
rect 177348 79872 177404 79928
rect 177578 79872 177634 79928
rect 176842 77832 176898 77888
rect 176842 77016 176898 77072
rect 177026 78104 177082 78160
rect 177302 79192 177358 79248
rect 177210 71440 177266 71496
rect 177486 79736 177542 79792
rect 177394 77560 177450 77616
rect 177854 79736 177910 79792
rect 177578 78512 177634 78568
rect 177670 77832 177726 77888
rect 177486 75112 177542 75168
rect 178130 80552 178186 80608
rect 182546 80688 182602 80744
rect 178498 80280 178554 80336
rect 178038 79192 178094 79248
rect 178222 78648 178278 78704
rect 178038 78376 178094 78432
rect 178314 78376 178370 78432
rect 178682 79464 178738 79520
rect 178590 77424 178646 77480
rect 185214 80300 185270 80336
rect 185214 80280 185216 80300
rect 185216 80280 185268 80300
rect 185268 80280 185270 80300
rect 178866 78648 178922 78704
rect 179418 77288 179474 77344
rect 179878 77152 179934 77208
rect 180338 77288 180394 77344
rect 181350 77152 181406 77208
rect 181534 71712 181590 71768
rect 182086 71440 182142 71496
rect 182086 71032 182142 71088
rect 186870 139168 186926 139224
rect 186870 139032 186926 139088
rect 186594 64776 186650 64832
rect 186594 64368 186650 64424
rect 187146 145560 187202 145616
rect 187422 213832 187478 213888
rect 187422 139032 187478 139088
rect 187606 71712 187662 71768
rect 186870 60560 186926 60616
rect 187974 262248 188030 262304
rect 188526 146240 188582 146296
rect 187974 143384 188030 143440
rect 188066 142976 188122 143032
rect 187790 61784 187846 61840
rect 187790 59064 187846 59120
rect 187790 58792 187846 58848
rect 188250 139304 188306 139360
rect 188710 139712 188766 139768
rect 188526 75248 188582 75304
rect 189262 194928 189318 194984
rect 190366 199824 190422 199880
rect 190366 192616 190422 192672
rect 189078 67496 189134 67552
rect 189078 66952 189134 67008
rect 189170 63144 189226 63200
rect 188342 58792 188398 58848
rect 189538 67496 189594 67552
rect 190366 71712 190422 71768
rect 189998 60152 190054 60208
rect 189354 53488 189410 53544
rect 188066 52128 188122 52184
rect 187974 50632 188030 50688
rect 190734 61648 190790 61704
rect 190642 57840 190698 57896
rect 190550 53760 190606 53816
rect 191286 140256 191342 140312
rect 191102 139304 191158 139360
rect 191194 138624 191250 138680
rect 191286 81096 191342 81152
rect 192298 262248 192354 262304
rect 192114 76880 192170 76936
rect 192114 76472 192170 76528
rect 193126 146104 193182 146160
rect 192666 137944 192722 138000
rect 193126 145560 193182 145616
rect 192942 76472 192998 76528
rect 192482 68176 192538 68232
rect 191930 60424 191986 60480
rect 191838 58656 191894 58712
rect 190826 53080 190882 53136
rect 190458 45328 190514 45384
rect 193126 60424 193182 60480
rect 193126 60016 193182 60072
rect 193862 146240 193918 146296
rect 194046 146104 194102 146160
rect 193954 80824 194010 80880
rect 193862 67224 193918 67280
rect 193310 55800 193366 55856
rect 193218 48048 193274 48104
rect 194046 66156 194102 66192
rect 194046 66136 194048 66156
rect 194048 66136 194100 66156
rect 194100 66136 194102 66156
rect 195058 145968 195114 146024
rect 195978 198636 195980 198656
rect 195980 198636 196032 198656
rect 196032 198636 196034 198656
rect 195978 198600 196034 198636
rect 195518 179288 195574 179344
rect 195334 76608 195390 76664
rect 194782 59200 194838 59256
rect 195058 59200 195114 59256
rect 195058 58520 195114 58576
rect 194690 55120 194746 55176
rect 194598 52264 194654 52320
rect 194598 51992 194654 52048
rect 196806 139032 196862 139088
rect 196806 80008 196862 80064
rect 196254 68876 196310 68912
rect 196254 68856 196256 68876
rect 196256 68856 196308 68876
rect 196308 68856 196310 68876
rect 196162 56480 196218 56536
rect 196162 55936 196218 55992
rect 196070 53624 196126 53680
rect 196070 53216 196126 53272
rect 195978 50768 196034 50824
rect 196438 50768 196494 50824
rect 196438 50496 196494 50552
rect 194506 48048 194562 48104
rect 194506 47776 194562 47832
rect 197358 49408 197414 49464
rect 234618 278024 234674 278080
rect 299478 276664 299534 276720
rect 396722 284824 396778 284880
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580262 365064 580318 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 477498 262792 477554 262848
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580446 232328 580502 232384
rect 580354 219000 580410 219056
rect 579802 205672 579858 205728
rect 198186 147736 198242 147792
rect 198186 138896 198242 138952
rect 198738 146240 198794 146296
rect 198738 78376 198794 78432
rect 197726 64640 197782 64696
rect 197726 64232 197782 64288
rect 197542 52400 197598 52456
rect 198002 52400 198058 52456
rect 198002 51720 198058 51776
rect 198462 49408 198518 49464
rect 198462 49136 198518 49192
rect 201498 200232 201554 200288
rect 198922 196560 198978 196616
rect 199106 77424 199162 77480
rect 199014 63280 199070 63336
rect 199566 145560 199622 145616
rect 199566 70352 199622 70408
rect 200118 138760 200174 138816
rect 199382 63280 199438 63336
rect 199382 63008 199438 63064
rect 198922 57296 198978 57352
rect 198830 54984 198886 55040
rect 198830 54440 198886 54496
rect 200210 50904 200266 50960
rect 200486 195200 200542 195256
rect 200670 78240 200726 78296
rect 200946 138080 201002 138136
rect 200578 71576 200634 71632
rect 201406 150340 201462 150376
rect 201406 150320 201408 150340
rect 201408 150320 201460 150340
rect 201460 150320 201462 150340
rect 201406 71576 201462 71632
rect 201406 71032 201462 71088
rect 201038 68720 201094 68776
rect 201406 68720 201462 68776
rect 201406 68176 201462 68232
rect 200854 67496 200910 67552
rect 200486 62056 200542 62112
rect 201406 62056 201462 62112
rect 201406 61512 201462 61568
rect 200394 59880 200450 59936
rect 200670 56480 200726 56536
rect 201958 200096 202014 200152
rect 201406 50904 201462 50960
rect 201406 50360 201462 50416
rect 200302 48184 200358 48240
rect 201406 48184 201462 48240
rect 201406 47640 201462 47696
rect 202970 195336 203026 195392
rect 202142 152360 202198 152416
rect 202786 150356 202788 150376
rect 202788 150356 202840 150376
rect 202840 150356 202842 150376
rect 202786 150320 202842 150356
rect 201774 49544 201830 49600
rect 201682 46824 201738 46880
rect 201590 45464 201646 45520
rect 201590 45056 201646 45112
rect 202786 49544 202842 49600
rect 202786 49000 202842 49056
rect 202786 46824 202842 46880
rect 202786 46144 202842 46200
rect 202326 44104 202382 44160
rect 203154 196696 203210 196752
rect 204442 192616 204498 192672
rect 204442 78104 204498 78160
rect 204350 77016 204406 77072
rect 203614 76744 203670 76800
rect 203154 56344 203210 56400
rect 202970 49272 203026 49328
rect 202878 43968 202934 44024
rect 202326 43560 202382 43616
rect 202878 43424 202934 43480
rect 204166 56344 204222 56400
rect 204166 55800 204222 55856
rect 204166 49272 204222 49328
rect 204166 48864 204222 48920
rect 205638 192480 205694 192536
rect 204718 50224 204774 50280
rect 205822 74432 205878 74488
rect 205822 73752 205878 73808
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580354 152632 580410 152688
rect 206006 75792 206062 75848
rect 580262 146376 580318 146432
rect 327722 139576 327778 139632
rect 206466 80688 206522 80744
rect 206282 78784 206338 78840
rect 206190 75656 206246 75712
rect 205730 63416 205786 63472
rect 205638 44920 205694 44976
rect 204534 44784 204590 44840
rect 208398 46280 208454 46336
rect 213918 67088 213974 67144
rect 213366 7520 213422 7576
rect 218058 71304 218114 71360
rect 220818 68312 220874 68368
rect 231858 56072 231914 56128
rect 229098 42064 229154 42120
rect 245658 61920 245714 61976
rect 242990 29552 243046 29608
rect 249798 58928 249854 58984
rect 264242 77832 264298 77888
rect 256698 64368 256754 64424
rect 259458 63280 259514 63336
rect 269118 73752 269174 73808
rect 263598 60288 263654 60344
rect 264978 12960 265034 13016
rect 277398 61784 277454 61840
rect 281538 58792 281594 58848
rect 282918 26832 282974 26888
rect 292578 63144 292634 63200
rect 299478 60152 299534 60208
rect 306378 79736 306434 79792
rect 309138 61648 309194 61704
rect 313278 57432 313334 57488
rect 315302 45192 315358 45248
rect 320178 53488 320234 53544
rect 382278 80144 382334 80200
rect 331218 58656 331274 58712
rect 338118 60016 338174 60072
rect 336278 6160 336334 6216
rect 351918 53352 351974 53408
rect 356058 50632 356114 50688
rect 362958 58520 363014 58576
rect 364982 54576 365038 54632
rect 369858 51992 369914 52048
rect 374090 51856 374146 51912
rect 389178 76472 389234 76528
rect 382922 55936 382978 55992
rect 387798 53216 387854 53272
rect 390558 50496 390614 50552
rect 400954 51720 401010 51776
rect 405738 49136 405794 49192
rect 408498 47776 408554 47832
rect 423678 66952 423734 67008
rect 414662 63008 414718 63064
rect 418802 57296 418858 57352
rect 423770 54440 423826 54496
rect 440238 61512 440294 61568
rect 433338 53080 433394 53136
rect 437478 50360 437534 50416
rect 444378 47640 444434 47696
rect 448610 43560 448666 43616
rect 475382 75248 475438 75304
rect 455418 49000 455474 49056
rect 458178 45056 458234 45112
rect 462318 46144 462374 46200
rect 466458 48864 466514 48920
rect 476118 43424 476174 43480
rect 481638 55800 481694 55856
rect 576122 139440 576178 139496
rect 494058 71168 494114 71224
rect 498198 69536 498254 69592
rect 496082 66816 496138 66872
rect 507858 65456 507914 65512
rect 511998 64232 512054 64288
rect 514022 62872 514078 62928
rect 520922 47504 520978 47560
rect 525062 59880 525118 59936
rect 549258 75112 549314 75168
rect 543738 71032 543794 71088
rect 539690 68176 539746 68232
rect 547878 64096 547934 64152
rect 545762 57160 545818 57216
rect 553398 44920 553454 44976
rect 567842 62736 567898 62792
rect 563702 61376 563758 61432
rect 565818 44784 565874 44840
rect 569958 50224 570014 50280
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580262 99456 580318 99512
rect 580170 86128 580226 86184
rect 580262 79328 580318 79384
rect 579986 72936 580042 72992
rect 581090 78512 581146 78568
rect 580262 59608 580318 59664
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect 396717 284882 396783 284885
rect 190410 284880 396783 284882
rect 190410 284824 396722 284880
rect 396778 284824 396783 284880
rect 190410 284822 396783 284824
rect 150433 284338 150499 284341
rect 187366 284338 187372 284340
rect 150433 284336 187372 284338
rect 150433 284280 150438 284336
rect 150494 284280 187372 284336
rect 150433 284278 187372 284280
rect 150433 284275 150499 284278
rect 187366 284276 187372 284278
rect 187436 284338 187442 284340
rect 190410 284338 190470 284822
rect 396717 284819 396783 284822
rect 187436 284278 190470 284338
rect 187436 284276 187442 284278
rect -960 279972 480 280212
rect 189022 278020 189028 278084
rect 189092 278082 189098 278084
rect 234613 278082 234679 278085
rect 189092 278080 234679 278082
rect 189092 278024 234618 278080
rect 234674 278024 234679 278080
rect 189092 278022 234679 278024
rect 189092 278020 189098 278022
rect 234613 278019 234679 278022
rect 156045 277538 156111 277541
rect 189022 277538 189028 277540
rect 156045 277536 189028 277538
rect 156045 277480 156050 277536
rect 156106 277480 189028 277536
rect 156045 277478 189028 277480
rect 156045 277475 156111 277478
rect 189022 277476 189028 277478
rect 189092 277476 189098 277540
rect 299473 276722 299539 276725
rect 190410 276720 299539 276722
rect 190410 276664 299478 276720
rect 299534 276664 299539 276720
rect 190410 276662 299539 276664
rect 153377 276042 153443 276045
rect 187734 276042 187740 276044
rect 153377 276040 187740 276042
rect 153377 275984 153382 276040
rect 153438 275984 187740 276040
rect 153377 275982 187740 275984
rect 153377 275979 153443 275982
rect 187734 275980 187740 275982
rect 187804 276042 187810 276044
rect 190410 276042 190470 276662
rect 299473 276659 299539 276662
rect 187804 275982 190470 276042
rect 187804 275980 187810 275982
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 167545 265434 167611 265437
rect 196198 265434 196204 265436
rect 167545 265432 196204 265434
rect 167545 265376 167550 265432
rect 167606 265376 196204 265432
rect 167545 265374 196204 265376
rect 167545 265371 167611 265374
rect 196198 265372 196204 265374
rect 196268 265372 196274 265436
rect 160829 265298 160895 265301
rect 193254 265298 193260 265300
rect 160829 265296 193260 265298
rect 160829 265240 160834 265296
rect 160890 265240 193260 265296
rect 160829 265238 193260 265240
rect 160829 265235 160895 265238
rect 193254 265236 193260 265238
rect 193324 265236 193330 265300
rect 112846 265100 112852 265164
rect 112916 265162 112922 265164
rect 135897 265162 135963 265165
rect 112916 265160 135963 265162
rect 112916 265104 135902 265160
rect 135958 265104 135963 265160
rect 112916 265102 135963 265104
rect 112916 265100 112922 265102
rect 135897 265099 135963 265102
rect 162209 265162 162275 265165
rect 194726 265162 194732 265164
rect 162209 265160 194732 265162
rect 162209 265104 162214 265160
rect 162270 265104 194732 265160
rect 162209 265102 194732 265104
rect 162209 265099 162275 265102
rect 194726 265100 194732 265102
rect 194796 265100 194802 265164
rect 113030 264964 113036 265028
rect 113100 265026 113106 265028
rect 138749 265026 138815 265029
rect 113100 265024 138815 265026
rect 113100 264968 138754 265024
rect 138810 264968 138815 265024
rect 113100 264966 138815 264968
rect 113100 264964 113106 264966
rect 138749 264963 138815 264966
rect 164877 265026 164943 265029
rect 165153 265026 165219 265029
rect 197486 265026 197492 265028
rect 164877 265024 197492 265026
rect 164877 264968 164882 265024
rect 164938 264968 165158 265024
rect 165214 264968 197492 265024
rect 164877 264966 197492 264968
rect 164877 264963 164943 264966
rect 165153 264963 165219 264966
rect 197486 264964 197492 264966
rect 197556 264964 197562 265028
rect 122598 263876 122604 263940
rect 122668 263938 122674 263940
rect 146201 263938 146267 263941
rect 122668 263936 146267 263938
rect 122668 263880 146206 263936
rect 146262 263880 146267 263936
rect 122668 263878 146267 263880
rect 122668 263876 122674 263878
rect 146201 263875 146267 263878
rect 115790 263740 115796 263804
rect 115860 263802 115866 263804
rect 145557 263802 145623 263805
rect 115860 263800 145623 263802
rect 115860 263744 145562 263800
rect 145618 263744 145623 263800
rect 115860 263742 145623 263744
rect 115860 263740 115866 263742
rect 145557 263739 145623 263742
rect 118366 263604 118372 263668
rect 118436 263666 118442 263668
rect 148593 263666 148659 263669
rect 118436 263664 148659 263666
rect 118436 263608 148598 263664
rect 148654 263608 148659 263664
rect 118436 263606 148659 263608
rect 118436 263604 118442 263606
rect 148593 263603 148659 263606
rect 116894 263196 116900 263260
rect 116964 263258 116970 263260
rect 129825 263258 129891 263261
rect 116964 263256 129891 263258
rect 116964 263200 129830 263256
rect 129886 263200 129891 263256
rect 116964 263198 129891 263200
rect 116964 263196 116970 263198
rect 129825 263195 129891 263198
rect 119838 263060 119844 263124
rect 119908 263122 119914 263124
rect 150525 263122 150591 263125
rect 163405 263122 163471 263125
rect 163589 263122 163655 263125
rect 119908 263120 151830 263122
rect 119908 263064 150530 263120
rect 150586 263064 151830 263120
rect 119908 263062 151830 263064
rect 119908 263060 119914 263062
rect 150525 263059 150591 263062
rect 113766 262924 113772 262988
rect 113836 262986 113842 262988
rect 138657 262986 138723 262989
rect 113836 262984 138723 262986
rect 113836 262928 138662 262984
rect 138718 262928 138723 262984
rect 113836 262926 138723 262928
rect 113836 262924 113842 262926
rect 138657 262923 138723 262926
rect 113950 262788 113956 262852
rect 114020 262850 114026 262852
rect 140313 262850 140379 262853
rect 114020 262848 140379 262850
rect 114020 262792 140318 262848
rect 140374 262792 140379 262848
rect 114020 262790 140379 262792
rect 151770 262850 151830 263062
rect 163405 263120 163655 263122
rect 163405 263064 163410 263120
rect 163466 263064 163594 263120
rect 163650 263064 163655 263120
rect 163405 263062 163655 263064
rect 163405 263059 163471 263062
rect 163589 263059 163655 263062
rect 477493 262850 477559 262853
rect 151770 262848 477559 262850
rect 151770 262792 477498 262848
rect 477554 262792 477559 262848
rect 151770 262790 477559 262792
rect 114020 262788 114026 262790
rect 140313 262787 140379 262790
rect 477493 262787 477559 262790
rect 118182 262652 118188 262716
rect 118252 262714 118258 262716
rect 146937 262714 147003 262717
rect 118252 262712 147003 262714
rect 118252 262656 146942 262712
rect 146998 262656 147003 262712
rect 118252 262654 147003 262656
rect 118252 262652 118258 262654
rect 146937 262651 147003 262654
rect 162025 262714 162091 262717
rect 193438 262714 193444 262716
rect 162025 262712 193444 262714
rect 162025 262656 162030 262712
rect 162086 262656 193444 262712
rect 162025 262654 193444 262656
rect 162025 262651 162091 262654
rect 193438 262652 193444 262654
rect 193508 262652 193514 262716
rect 115422 262516 115428 262580
rect 115492 262578 115498 262580
rect 144177 262578 144243 262581
rect 115492 262576 144243 262578
rect 115492 262520 144182 262576
rect 144238 262520 144243 262576
rect 115492 262518 144243 262520
rect 115492 262516 115498 262518
rect 144177 262515 144243 262518
rect 164969 262578 165035 262581
rect 192150 262578 192156 262580
rect 164969 262576 192156 262578
rect 164969 262520 164974 262576
rect 165030 262520 192156 262576
rect 164969 262518 192156 262520
rect 164969 262515 165035 262518
rect 192150 262516 192156 262518
rect 192220 262516 192226 262580
rect 114134 262380 114140 262444
rect 114204 262442 114210 262444
rect 142153 262442 142219 262445
rect 142889 262442 142955 262445
rect 114204 262440 142955 262442
rect 114204 262384 142158 262440
rect 142214 262384 142894 262440
rect 142950 262384 142955 262440
rect 114204 262382 142955 262384
rect 114204 262380 114210 262382
rect 142153 262379 142219 262382
rect 142889 262379 142955 262382
rect 163405 262442 163471 262445
rect 191966 262442 191972 262444
rect 163405 262440 191972 262442
rect 163405 262384 163410 262440
rect 163466 262384 191972 262440
rect 163405 262382 191972 262384
rect 163405 262379 163471 262382
rect 191966 262380 191972 262382
rect 192036 262380 192042 262444
rect 187969 262308 188035 262309
rect 187918 262306 187924 262308
rect 187878 262246 187924 262306
rect 187988 262304 188035 262308
rect 188030 262248 188035 262304
rect 187918 262244 187924 262246
rect 187988 262244 188035 262248
rect 187969 262243 188035 262244
rect 192293 262308 192359 262309
rect 192293 262304 192340 262308
rect 192404 262306 192410 262308
rect 192293 262248 192298 262304
rect 192293 262244 192340 262248
rect 192404 262246 192450 262306
rect 192404 262244 192410 262246
rect 192293 262243 192359 262244
rect 117957 261218 118023 261221
rect 127617 261218 127683 261221
rect 117957 261216 127683 261218
rect 117957 261160 117962 261216
rect 118018 261160 127622 261216
rect 127678 261160 127683 261216
rect 117957 261158 127683 261160
rect 117957 261155 118023 261158
rect 127617 261155 127683 261158
rect 111558 261020 111564 261084
rect 111628 261082 111634 261084
rect 133965 261082 134031 261085
rect 111628 261080 134031 261082
rect 111628 261024 133970 261080
rect 134026 261024 134031 261080
rect 111628 261022 134031 261024
rect 111628 261020 111634 261022
rect 133965 261019 134031 261022
rect 111374 260884 111380 260948
rect 111444 260946 111450 260948
rect 117957 260946 118023 260949
rect 111444 260944 118023 260946
rect 111444 260888 117962 260944
rect 118018 260888 118023 260944
rect 111444 260886 118023 260888
rect 111444 260884 111450 260886
rect 117957 260883 118023 260886
rect 127617 260946 127683 260949
rect 137461 260946 137527 260949
rect 127617 260944 137527 260946
rect 127617 260888 127622 260944
rect 127678 260888 137466 260944
rect 137522 260888 137527 260944
rect 127617 260886 137527 260888
rect 127617 260883 127683 260886
rect 137461 260883 137527 260886
rect 158713 260946 158779 260949
rect 193622 260946 193628 260948
rect 158713 260944 193628 260946
rect 158713 260888 158718 260944
rect 158774 260888 193628 260944
rect 158713 260886 193628 260888
rect 158713 260883 158779 260886
rect 193622 260884 193628 260886
rect 193692 260884 193698 260948
rect 115606 260476 115612 260540
rect 115676 260538 115682 260540
rect 124857 260538 124923 260541
rect 115676 260536 124923 260538
rect 115676 260480 124862 260536
rect 124918 260480 124923 260536
rect 115676 260478 124923 260480
rect 115676 260476 115682 260478
rect 124857 260475 124923 260478
rect 117078 260340 117084 260404
rect 117148 260402 117154 260404
rect 117148 260342 148610 260402
rect 117148 260340 117154 260342
rect 120942 260204 120948 260268
rect 121012 260266 121018 260268
rect 143625 260266 143691 260269
rect 144499 260266 144565 260269
rect 121012 260264 144565 260266
rect 121012 260208 143630 260264
rect 143686 260208 144504 260264
rect 144560 260208 144565 260264
rect 121012 260206 144565 260208
rect 121012 260204 121018 260206
rect 143625 260203 143691 260206
rect 144499 260203 144565 260206
rect 147673 260266 147739 260269
rect 148363 260266 148429 260269
rect 147673 260264 148429 260266
rect 147673 260208 147678 260264
rect 147734 260208 148368 260264
rect 148424 260208 148429 260264
rect 147673 260206 148429 260208
rect 148550 260266 148610 260342
rect 149053 260266 149119 260269
rect 150019 260266 150085 260269
rect 148550 260264 150085 260266
rect 148550 260208 149058 260264
rect 149114 260208 150024 260264
rect 150080 260208 150085 260264
rect 148550 260206 150085 260208
rect 147673 260203 147739 260206
rect 148363 260203 148429 260206
rect 149053 260203 149119 260206
rect 150019 260203 150085 260206
rect 155953 260266 156019 260269
rect 156643 260266 156709 260269
rect 155953 260264 156709 260266
rect 155953 260208 155958 260264
rect 156014 260208 156648 260264
rect 156704 260208 156709 260264
rect 155953 260206 156709 260208
rect 155953 260203 156019 260206
rect 156643 260203 156709 260206
rect 160093 260266 160159 260269
rect 161059 260266 161125 260269
rect 160093 260264 161125 260266
rect 160093 260208 160098 260264
rect 160154 260208 161064 260264
rect 161120 260208 161125 260264
rect 160093 260206 161125 260208
rect 160093 260203 160159 260206
rect 161059 260203 161125 260206
rect 161473 260266 161539 260269
rect 162715 260266 162781 260269
rect 161473 260264 162781 260266
rect 161473 260208 161478 260264
rect 161534 260208 162720 260264
rect 162776 260208 162781 260264
rect 161473 260206 162781 260208
rect 161473 260203 161539 260206
rect 162715 260203 162781 260206
rect 118550 260068 118556 260132
rect 118620 260130 118626 260132
rect 142245 260130 142311 260133
rect 143395 260130 143461 260133
rect 118620 260128 143461 260130
rect 118620 260072 142250 260128
rect 142306 260072 143400 260128
rect 143456 260072 143461 260128
rect 118620 260070 143461 260072
rect 118620 260068 118626 260070
rect 142245 260067 142311 260070
rect 143395 260067 143461 260070
rect 181345 260130 181411 260133
rect 189390 260130 189396 260132
rect 181345 260128 189396 260130
rect 181345 260072 181350 260128
rect 181406 260072 189396 260128
rect 181345 260070 189396 260072
rect 181345 260067 181411 260070
rect 189390 260068 189396 260070
rect 189460 260068 189466 260132
rect 119654 259932 119660 259996
rect 119724 259994 119730 259996
rect 144913 259994 144979 259997
rect 119724 259992 144979 259994
rect 119724 259936 144918 259992
rect 144974 259936 144979 259992
rect 119724 259934 144979 259936
rect 119724 259932 119730 259934
rect 144913 259931 144979 259934
rect 162853 259994 162919 259997
rect 188102 259994 188108 259996
rect 162853 259992 188108 259994
rect 162853 259936 162858 259992
rect 162914 259936 188108 259992
rect 162853 259934 188108 259936
rect 162853 259931 162919 259934
rect 188102 259932 188108 259934
rect 188172 259932 188178 259996
rect 122230 259796 122236 259860
rect 122300 259858 122306 259860
rect 149237 259858 149303 259861
rect 122300 259856 149303 259858
rect 122300 259800 149242 259856
rect 149298 259800 149303 259856
rect 122300 259798 149303 259800
rect 122300 259796 122306 259798
rect 149237 259795 149303 259798
rect 161197 259858 161263 259861
rect 188286 259858 188292 259860
rect 161197 259856 188292 259858
rect 161197 259800 161202 259856
rect 161258 259800 188292 259856
rect 161197 259798 188292 259800
rect 161197 259795 161263 259798
rect 188286 259796 188292 259798
rect 188356 259796 188362 259860
rect 116710 259660 116716 259724
rect 116780 259722 116786 259724
rect 148133 259722 148199 259725
rect 116780 259720 148199 259722
rect 116780 259664 148138 259720
rect 148194 259664 148199 259720
rect 116780 259662 148199 259664
rect 116780 259660 116786 259662
rect 148133 259659 148199 259662
rect 156873 259722 156939 259725
rect 181345 259722 181411 259725
rect 189574 259722 189580 259724
rect 156873 259720 181411 259722
rect 156873 259664 156878 259720
rect 156934 259664 181350 259720
rect 181406 259664 181411 259720
rect 156873 259662 181411 259664
rect 156873 259659 156939 259662
rect 181345 259659 181411 259662
rect 181486 259662 189580 259722
rect 121177 259588 121243 259589
rect 121126 259586 121132 259588
rect 121086 259526 121132 259586
rect 121196 259584 121243 259588
rect 121238 259528 121243 259584
rect 121126 259524 121132 259526
rect 121196 259524 121243 259528
rect 123150 259524 123156 259588
rect 123220 259586 123226 259588
rect 123293 259586 123359 259589
rect 123220 259584 123359 259586
rect 123220 259528 123298 259584
rect 123354 259528 123359 259584
rect 123220 259526 123359 259528
rect 123220 259524 123226 259526
rect 121177 259523 121243 259524
rect 123293 259523 123359 259526
rect 123937 259586 124003 259589
rect 124070 259586 124076 259588
rect 123937 259584 124076 259586
rect 123937 259528 123942 259584
rect 123998 259528 124076 259584
rect 123937 259526 124076 259528
rect 123937 259523 124003 259526
rect 124070 259524 124076 259526
rect 124140 259524 124146 259588
rect 155217 259586 155283 259589
rect 181486 259586 181546 259662
rect 189574 259660 189580 259662
rect 189644 259660 189650 259724
rect 155217 259584 181546 259586
rect 155217 259528 155222 259584
rect 155278 259528 181546 259584
rect 155217 259526 181546 259528
rect 185669 259586 185735 259589
rect 186078 259586 186084 259588
rect 185669 259584 186084 259586
rect 185669 259528 185674 259584
rect 185730 259528 186084 259584
rect 185669 259526 186084 259528
rect 155217 259523 155283 259526
rect 185669 259523 185735 259526
rect 186078 259524 186084 259526
rect 186148 259524 186154 259588
rect 122833 259450 122899 259453
rect 122966 259450 122972 259452
rect 122833 259448 122972 259450
rect 122833 259392 122838 259448
rect 122894 259392 122972 259448
rect 122833 259390 122972 259392
rect 122833 259387 122899 259390
rect 122966 259388 122972 259390
rect 123036 259388 123042 259452
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 186078 213828 186084 213892
rect 186148 213890 186154 213892
rect 187417 213890 187483 213893
rect 186148 213888 187483 213890
rect 186148 213832 187422 213888
rect 187478 213832 187483 213888
rect 186148 213830 187483 213832
rect 186148 213828 186154 213830
rect 187417 213827 187483 213830
rect 122557 209674 122623 209677
rect 122782 209674 122788 209676
rect 122557 209672 122788 209674
rect 122557 209616 122562 209672
rect 122618 209616 122788 209672
rect 122557 209614 122788 209616
rect 122557 209611 122623 209614
rect 122782 209612 122788 209614
rect 122852 209612 122858 209676
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 122557 205594 122623 205597
rect 122782 205594 122788 205596
rect 122557 205592 122788 205594
rect 122557 205536 122562 205592
rect 122618 205536 122788 205592
rect 122557 205534 122788 205536
rect 122557 205531 122623 205534
rect 122782 205532 122788 205534
rect 122852 205532 122858 205596
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 104801 201106 104867 201109
rect 122557 201106 122623 201109
rect 104801 201104 122623 201106
rect 104801 201048 104806 201104
rect 104862 201048 122562 201104
rect 122618 201048 122623 201104
rect 104801 201046 122623 201048
rect 104801 201043 104867 201046
rect 122557 201043 122623 201046
rect 123886 200908 123892 200972
rect 123956 200970 123962 200972
rect 123956 200910 131130 200970
rect 123956 200908 123962 200910
rect 131070 200834 131130 200910
rect 153510 200908 153516 200972
rect 153580 200970 153586 200972
rect 170990 200970 170996 200972
rect 153580 200910 170996 200970
rect 153580 200908 153586 200910
rect 170990 200908 170996 200910
rect 171060 200908 171066 200972
rect 158110 200834 158116 200836
rect 131070 200774 158116 200834
rect 158110 200772 158116 200774
rect 158180 200772 158186 200836
rect 124029 200700 124095 200701
rect 124029 200698 124076 200700
rect 123984 200696 124076 200698
rect 123984 200640 124034 200696
rect 123984 200638 124076 200640
rect 124029 200636 124076 200638
rect 124140 200636 124146 200700
rect 156270 200636 156276 200700
rect 156340 200698 156346 200700
rect 173750 200698 173756 200700
rect 156340 200638 173756 200698
rect 156340 200636 156346 200638
rect 173750 200636 173756 200638
rect 173820 200636 173826 200700
rect 124029 200635 124095 200636
rect 122966 200500 122972 200564
rect 123036 200562 123042 200564
rect 124121 200562 124187 200565
rect 123036 200560 124187 200562
rect 123036 200504 124126 200560
rect 124182 200504 124187 200560
rect 123036 200502 124187 200504
rect 123036 200500 123042 200502
rect 124121 200499 124187 200502
rect 132033 200562 132099 200565
rect 142838 200562 142844 200564
rect 132033 200560 142844 200562
rect 132033 200504 132038 200560
rect 132094 200504 142844 200560
rect 132033 200502 142844 200504
rect 132033 200499 132099 200502
rect 142838 200500 142844 200502
rect 142908 200500 142914 200564
rect 180742 200562 180748 200564
rect 151494 200502 180748 200562
rect 107285 200426 107351 200429
rect 126605 200426 126671 200429
rect 107285 200424 126671 200426
rect 107285 200368 107290 200424
rect 107346 200368 126610 200424
rect 126666 200368 126671 200424
rect 107285 200366 126671 200368
rect 107285 200363 107351 200366
rect 126605 200363 126671 200366
rect 131941 200426 132007 200429
rect 138974 200426 138980 200428
rect 131941 200424 138980 200426
rect 131941 200368 131946 200424
rect 132002 200368 138980 200424
rect 131941 200366 138980 200368
rect 131941 200363 132007 200366
rect 138974 200364 138980 200366
rect 139044 200364 139050 200428
rect 128905 200290 128971 200293
rect 128905 200288 148242 200290
rect 128905 200232 128910 200288
rect 128966 200232 148242 200288
rect 128905 200230 148242 200232
rect 128905 200227 128971 200230
rect 107377 200154 107443 200157
rect 130193 200154 130259 200157
rect 107377 200152 130259 200154
rect 107377 200096 107382 200152
rect 107438 200096 130198 200152
rect 130254 200096 130259 200152
rect 107377 200094 130259 200096
rect 107377 200091 107443 200094
rect 130193 200091 130259 200094
rect 131573 200154 131639 200157
rect 131573 200152 145804 200154
rect 131573 200096 131578 200152
rect 131634 200096 145804 200152
rect 131573 200094 145804 200096
rect 131573 200091 131639 200094
rect 131941 200018 132007 200021
rect 131941 200016 136466 200018
rect 131941 199960 131946 200016
rect 132002 199960 136466 200016
rect 131941 199958 136466 199960
rect 131941 199955 132007 199958
rect 132534 199820 132540 199884
rect 132604 199882 132610 199884
rect 132815 199882 132881 199885
rect 132604 199880 132881 199882
rect 132604 199824 132820 199880
rect 132876 199824 132881 199880
rect 132604 199822 132881 199824
rect 132604 199820 132610 199822
rect 132815 199819 132881 199822
rect 133086 199820 133092 199884
rect 133156 199882 133162 199884
rect 133367 199882 133433 199885
rect 133156 199880 133433 199882
rect 133156 199824 133372 199880
rect 133428 199824 133433 199880
rect 133156 199822 133433 199824
rect 133156 199820 133162 199822
rect 133367 199819 133433 199822
rect 134006 199820 134012 199884
rect 134076 199882 134082 199884
rect 134287 199882 134353 199885
rect 134076 199880 134353 199882
rect 134076 199824 134292 199880
rect 134348 199824 134353 199880
rect 134076 199822 134353 199824
rect 134076 199820 134082 199822
rect 134287 199819 134353 199822
rect 134558 199820 134564 199884
rect 134628 199882 134634 199884
rect 134839 199882 134905 199885
rect 134628 199880 134905 199882
rect 134628 199824 134844 199880
rect 134900 199824 134905 199880
rect 134628 199822 134905 199824
rect 134628 199820 134634 199822
rect 134839 199819 134905 199822
rect 135575 199882 135641 199885
rect 136219 199884 136285 199885
rect 135846 199882 135852 199884
rect 135575 199880 135852 199882
rect 135575 199824 135580 199880
rect 135636 199824 135852 199880
rect 135575 199822 135852 199824
rect 135575 199819 135641 199822
rect 135846 199820 135852 199822
rect 135916 199820 135922 199884
rect 136214 199882 136220 199884
rect 136128 199822 136220 199882
rect 136214 199820 136220 199822
rect 136284 199820 136290 199884
rect 136406 199882 136466 199958
rect 136771 199914 136837 199919
rect 136771 199882 136776 199914
rect 136406 199858 136776 199882
rect 136832 199858 136837 199914
rect 137875 199914 137941 199919
rect 137139 199884 137205 199885
rect 137507 199884 137573 199885
rect 137134 199882 137140 199884
rect 136406 199853 136837 199858
rect 136406 199822 136834 199853
rect 137048 199822 137140 199882
rect 137134 199820 137140 199822
rect 137204 199820 137210 199884
rect 137502 199882 137508 199884
rect 137416 199822 137508 199882
rect 137502 199820 137508 199822
rect 137572 199820 137578 199884
rect 137686 199820 137692 199884
rect 137756 199882 137762 199884
rect 137875 199882 137880 199914
rect 137756 199858 137880 199882
rect 137936 199858 137941 199914
rect 142107 199914 142173 199919
rect 137756 199853 137941 199858
rect 138151 199882 138217 199885
rect 138422 199882 138428 199884
rect 138151 199880 138428 199882
rect 137756 199822 137938 199853
rect 138151 199824 138156 199880
rect 138212 199824 138428 199880
rect 138151 199822 138428 199824
rect 137756 199820 137762 199822
rect 136219 199819 136285 199820
rect 137139 199819 137205 199820
rect 137507 199819 137573 199820
rect 138151 199819 138217 199822
rect 138422 199820 138428 199822
rect 138492 199820 138498 199884
rect 141918 199882 141924 199884
rect 140316 199822 141924 199882
rect 121269 199746 121335 199749
rect 140316 199746 140376 199822
rect 141918 199820 141924 199822
rect 141988 199820 141994 199884
rect 142107 199858 142112 199914
rect 142168 199858 142173 199914
rect 142107 199853 142173 199858
rect 142475 199914 142541 199919
rect 142475 199858 142480 199914
rect 142536 199882 142541 199914
rect 143487 199914 143553 199919
rect 142654 199882 142660 199884
rect 142536 199858 142660 199882
rect 142475 199853 142660 199858
rect 121269 199744 140376 199746
rect 121269 199688 121274 199744
rect 121330 199688 140376 199744
rect 121269 199686 140376 199688
rect 121269 199683 121335 199686
rect 140446 199684 140452 199748
rect 140516 199746 140522 199748
rect 142110 199746 142170 199853
rect 142478 199822 142660 199853
rect 142654 199820 142660 199822
rect 142724 199820 142730 199884
rect 142838 199820 142844 199884
rect 142908 199882 142914 199884
rect 143487 199882 143492 199914
rect 142908 199858 143492 199882
rect 143548 199858 143553 199914
rect 144131 199914 144197 199919
rect 144131 199884 144136 199914
rect 144192 199884 144197 199914
rect 144315 199914 144381 199919
rect 142908 199853 143553 199858
rect 142908 199822 143550 199853
rect 142908 199820 142914 199822
rect 144126 199820 144132 199884
rect 144196 199882 144202 199884
rect 144196 199822 144254 199882
rect 144315 199858 144320 199914
rect 144376 199858 144381 199914
rect 144315 199853 144381 199858
rect 144499 199914 144565 199919
rect 144499 199858 144504 199914
rect 144560 199858 144565 199914
rect 145511 199914 145577 199919
rect 144499 199853 144565 199858
rect 144867 199880 144933 199885
rect 144196 199820 144202 199822
rect 144318 199746 144378 199853
rect 140516 199686 142170 199746
rect 142662 199686 144378 199746
rect 144502 199749 144562 199853
rect 144867 199824 144872 199880
rect 144928 199824 144933 199880
rect 145511 199858 145516 199914
rect 145572 199858 145577 199914
rect 145511 199853 145577 199858
rect 145744 199882 145804 200094
rect 147995 199914 148061 199919
rect 145879 199882 145945 199885
rect 147995 199882 148000 199914
rect 145744 199880 145945 199882
rect 144867 199819 144933 199824
rect 144502 199744 144611 199749
rect 144502 199688 144550 199744
rect 144606 199688 144611 199744
rect 144502 199686 144611 199688
rect 140516 199684 140522 199686
rect 128813 199610 128879 199613
rect 142429 199610 142495 199613
rect 128813 199608 142495 199610
rect 128813 199552 128818 199608
rect 128874 199552 142434 199608
rect 142490 199552 142495 199608
rect 128813 199550 142495 199552
rect 128813 199547 128879 199550
rect 142429 199547 142495 199550
rect 126605 199474 126671 199477
rect 135345 199474 135411 199477
rect 126605 199472 135411 199474
rect 126605 199416 126610 199472
rect 126666 199416 135350 199472
rect 135406 199416 135411 199472
rect 126605 199414 135411 199416
rect 126605 199411 126671 199414
rect 135345 199411 135411 199414
rect 136541 199474 136607 199477
rect 137369 199474 137435 199477
rect 136541 199472 137435 199474
rect 136541 199416 136546 199472
rect 136602 199416 137374 199472
rect 137430 199416 137435 199472
rect 136541 199414 137435 199416
rect 136541 199411 136607 199414
rect 137369 199411 137435 199414
rect 138197 199474 138263 199477
rect 138841 199476 138907 199477
rect 138422 199474 138428 199476
rect 138197 199472 138428 199474
rect 138197 199416 138202 199472
rect 138258 199416 138428 199472
rect 138197 199414 138428 199416
rect 138197 199411 138263 199414
rect 138422 199412 138428 199414
rect 138492 199412 138498 199476
rect 138790 199474 138796 199476
rect 138750 199414 138796 199474
rect 138860 199472 138907 199476
rect 138902 199416 138907 199472
rect 138790 199412 138796 199414
rect 138860 199412 138907 199416
rect 138974 199412 138980 199476
rect 139044 199474 139050 199476
rect 142662 199474 142722 199686
rect 144545 199683 144611 199686
rect 144177 199610 144243 199613
rect 144870 199610 144930 199819
rect 145514 199749 145574 199853
rect 145744 199824 145884 199880
rect 145940 199824 145945 199880
rect 145744 199822 145945 199824
rect 145879 199819 145945 199822
rect 146158 199858 148000 199882
rect 148056 199858 148061 199914
rect 146158 199853 148061 199858
rect 146158 199822 148058 199853
rect 145465 199744 145574 199749
rect 145465 199688 145470 199744
rect 145526 199688 145574 199744
rect 145465 199686 145574 199688
rect 145465 199683 145531 199686
rect 144177 199608 144930 199610
rect 144177 199552 144182 199608
rect 144238 199552 144930 199608
rect 144177 199550 144930 199552
rect 144177 199547 144243 199550
rect 139044 199414 142722 199474
rect 145741 199474 145807 199477
rect 146158 199474 146218 199822
rect 146886 199684 146892 199748
rect 146956 199746 146962 199748
rect 147581 199746 147647 199749
rect 146956 199744 147647 199746
rect 146956 199688 147586 199744
rect 147642 199688 147647 199744
rect 146956 199686 147647 199688
rect 146956 199684 146962 199686
rect 147581 199683 147647 199686
rect 148182 199610 148242 200230
rect 148910 199956 148916 200020
rect 148980 200018 148986 200020
rect 148980 199958 150266 200018
rect 148980 199956 148986 199958
rect 148639 199916 148705 199919
rect 148596 199914 148705 199916
rect 148358 199820 148364 199884
rect 148428 199882 148434 199884
rect 148596 199882 148644 199914
rect 148428 199858 148644 199882
rect 148700 199858 148705 199914
rect 149651 199884 149717 199885
rect 150019 199884 150085 199885
rect 149646 199882 149652 199884
rect 148428 199853 148705 199858
rect 148428 199822 148656 199853
rect 149560 199822 149652 199882
rect 148428 199820 148434 199822
rect 149646 199820 149652 199822
rect 149716 199820 149722 199884
rect 150014 199882 150020 199884
rect 149928 199822 150020 199882
rect 150014 199820 150020 199822
rect 150084 199820 150090 199884
rect 150206 199882 150266 199958
rect 151494 199919 151554 200502
rect 180742 200500 180748 200502
rect 180812 200500 180818 200564
rect 178217 200426 178283 200429
rect 152460 200424 178283 200426
rect 152460 200368 178222 200424
rect 178278 200368 178283 200424
rect 152460 200366 178283 200368
rect 150479 199916 150545 199919
rect 150436 199914 150545 199916
rect 150436 199882 150484 199914
rect 150206 199858 150484 199882
rect 150540 199858 150545 199914
rect 151491 199914 151557 199919
rect 150206 199853 150545 199858
rect 151123 199882 151189 199885
rect 151302 199882 151308 199884
rect 151123 199880 151308 199882
rect 150206 199822 150496 199853
rect 151123 199824 151128 199880
rect 151184 199824 151308 199880
rect 151123 199822 151308 199824
rect 149651 199819 149717 199820
rect 150019 199819 150085 199820
rect 151123 199819 151189 199822
rect 151302 199820 151308 199822
rect 151372 199820 151378 199884
rect 151491 199858 151496 199914
rect 151552 199858 151557 199914
rect 151491 199853 151557 199858
rect 152319 199882 152385 199885
rect 152460 199882 152520 200366
rect 178217 200363 178283 200366
rect 168598 200228 168604 200292
rect 168668 200290 168674 200292
rect 201493 200290 201559 200293
rect 168668 200288 201559 200290
rect 168668 200232 201498 200288
rect 201554 200232 201559 200288
rect 168668 200230 201559 200232
rect 168668 200228 168674 200230
rect 201493 200227 201559 200230
rect 154806 200094 161306 200154
rect 154806 199919 154866 200094
rect 161246 200018 161306 200094
rect 161422 200092 161428 200156
rect 161492 200154 161498 200156
rect 161492 200094 169770 200154
rect 161492 200092 161498 200094
rect 165654 200018 165660 200020
rect 161246 199958 165660 200018
rect 165654 199956 165660 199958
rect 165724 199956 165730 200020
rect 154343 199916 154409 199919
rect 154343 199914 154452 199916
rect 152595 199884 152661 199885
rect 152319 199880 152520 199882
rect 152319 199824 152324 199880
rect 152380 199824 152520 199880
rect 152319 199822 152520 199824
rect 152319 199819 152385 199822
rect 152590 199820 152596 199884
rect 152660 199882 152666 199884
rect 152660 199822 152752 199882
rect 152660 199820 152666 199822
rect 153694 199820 153700 199884
rect 153764 199882 153770 199884
rect 153975 199882 154041 199885
rect 153764 199880 154041 199882
rect 153764 199824 153980 199880
rect 154036 199824 154041 199880
rect 154343 199858 154348 199914
rect 154404 199884 154452 199914
rect 154803 199914 154869 199919
rect 154404 199858 154436 199884
rect 154343 199853 154436 199858
rect 153764 199822 154041 199824
rect 154392 199822 154436 199853
rect 153764 199820 153770 199822
rect 152595 199819 152661 199820
rect 153975 199819 154041 199822
rect 154430 199820 154436 199822
rect 154500 199820 154506 199884
rect 154803 199858 154808 199914
rect 154864 199858 154869 199914
rect 154803 199853 154869 199858
rect 155263 199916 155329 199919
rect 155263 199914 155602 199916
rect 155263 199858 155268 199914
rect 155324 199884 155602 199914
rect 156827 199914 156893 199919
rect 155324 199858 155540 199884
rect 155263 199856 155540 199858
rect 155263 199853 155329 199856
rect 155534 199820 155540 199856
rect 155604 199820 155610 199884
rect 155718 199820 155724 199884
rect 155788 199882 155794 199884
rect 155999 199882 156065 199885
rect 156367 199882 156433 199885
rect 156827 199884 156832 199914
rect 156888 199884 156893 199914
rect 158299 199914 158365 199919
rect 155788 199880 156065 199882
rect 155788 199824 156004 199880
rect 156060 199824 156065 199880
rect 155788 199822 156065 199824
rect 155788 199820 155794 199822
rect 155999 199819 156065 199822
rect 156140 199880 156433 199882
rect 156140 199824 156372 199880
rect 156428 199824 156433 199880
rect 156140 199822 156433 199824
rect 150065 199746 150131 199749
rect 155309 199746 155375 199749
rect 155493 199746 155559 199749
rect 155769 199748 155835 199749
rect 155718 199746 155724 199748
rect 150065 199744 155234 199746
rect 150065 199688 150070 199744
rect 150126 199688 155234 199744
rect 150065 199686 155234 199688
rect 150065 199683 150131 199686
rect 150801 199610 150867 199613
rect 148182 199608 150867 199610
rect 148182 199552 150806 199608
rect 150862 199552 150867 199608
rect 148182 199550 150867 199552
rect 150801 199547 150867 199550
rect 152089 199610 152155 199613
rect 153510 199610 153516 199612
rect 152089 199608 153516 199610
rect 152089 199552 152094 199608
rect 152150 199552 153516 199608
rect 152089 199550 153516 199552
rect 152089 199547 152155 199550
rect 153510 199548 153516 199550
rect 153580 199548 153586 199612
rect 153878 199548 153884 199612
rect 153948 199610 153954 199612
rect 154021 199610 154087 199613
rect 153948 199608 154087 199610
rect 153948 199552 154026 199608
rect 154082 199552 154087 199608
rect 153948 199550 154087 199552
rect 155174 199610 155234 199686
rect 155309 199744 155559 199746
rect 155309 199688 155314 199744
rect 155370 199688 155498 199744
rect 155554 199688 155559 199744
rect 155309 199686 155559 199688
rect 155678 199686 155724 199746
rect 155788 199744 155835 199748
rect 155830 199688 155835 199744
rect 155309 199683 155375 199686
rect 155493 199683 155559 199686
rect 155718 199684 155724 199686
rect 155788 199684 155835 199688
rect 156140 199746 156200 199822
rect 156367 199819 156433 199822
rect 156822 199820 156828 199884
rect 156892 199882 156898 199884
rect 157747 199882 157813 199885
rect 158299 199884 158304 199914
rect 158360 199884 158365 199914
rect 165843 199914 165909 199919
rect 157926 199882 157932 199884
rect 156892 199822 156950 199882
rect 157747 199880 157932 199882
rect 157747 199824 157752 199880
rect 157808 199824 157932 199880
rect 157747 199822 157932 199824
rect 156892 199820 156898 199822
rect 157747 199819 157813 199822
rect 157926 199820 157932 199822
rect 157996 199820 158002 199884
rect 158294 199820 158300 199884
rect 158364 199882 158370 199884
rect 158364 199822 158422 199882
rect 158364 199820 158370 199822
rect 158662 199820 158668 199884
rect 158732 199882 158738 199884
rect 159035 199882 159101 199885
rect 159679 199882 159745 199885
rect 158732 199880 159101 199882
rect 158732 199824 159040 199880
rect 159096 199824 159101 199880
rect 158732 199822 159101 199824
rect 158732 199820 158738 199822
rect 159035 199819 159101 199822
rect 159406 199880 159745 199882
rect 159406 199824 159684 199880
rect 159740 199824 159745 199880
rect 159406 199822 159745 199824
rect 156321 199746 156387 199749
rect 156140 199744 156387 199746
rect 156140 199688 156326 199744
rect 156382 199688 156387 199744
rect 156140 199686 156387 199688
rect 155769 199683 155835 199684
rect 156321 199683 156387 199686
rect 158110 199684 158116 199748
rect 158180 199746 158186 199748
rect 158253 199746 158319 199749
rect 158180 199744 158319 199746
rect 158180 199688 158258 199744
rect 158314 199688 158319 199744
rect 158180 199686 158319 199688
rect 158180 199684 158186 199686
rect 158253 199683 158319 199686
rect 159030 199684 159036 199748
rect 159100 199746 159106 199748
rect 159406 199746 159466 199822
rect 159679 199819 159745 199822
rect 160870 199820 160876 199884
rect 160940 199882 160946 199884
rect 161059 199882 161125 199885
rect 163083 199884 163149 199885
rect 163078 199882 163084 199884
rect 160940 199880 161125 199882
rect 160940 199824 161064 199880
rect 161120 199824 161125 199880
rect 160940 199822 161125 199824
rect 162992 199822 163084 199882
rect 160940 199820 160946 199822
rect 161059 199819 161125 199822
rect 163078 199820 163084 199822
rect 163148 199820 163154 199884
rect 163262 199820 163268 199884
rect 163332 199882 163338 199884
rect 163727 199882 163793 199885
rect 163332 199880 163793 199882
rect 163332 199824 163732 199880
rect 163788 199824 163793 199880
rect 163332 199822 163793 199824
rect 163332 199820 163338 199822
rect 163083 199819 163149 199820
rect 163727 199819 163793 199822
rect 164003 199880 164069 199885
rect 164371 199884 164437 199885
rect 164366 199882 164372 199884
rect 164003 199824 164008 199880
rect 164064 199824 164069 199880
rect 164003 199819 164069 199824
rect 164280 199822 164372 199882
rect 164366 199820 164372 199822
rect 164436 199820 164442 199884
rect 164550 199820 164556 199884
rect 164620 199882 164626 199884
rect 164831 199882 164897 199885
rect 164620 199880 164897 199882
rect 164620 199824 164836 199880
rect 164892 199824 164897 199880
rect 164620 199822 164897 199824
rect 164620 199820 164626 199822
rect 164371 199819 164437 199820
rect 164831 199819 164897 199822
rect 165199 199882 165265 199885
rect 165843 199884 165848 199914
rect 165904 199884 165909 199914
rect 166395 199914 166461 199919
rect 166671 199916 166737 199919
rect 169063 199916 169129 199919
rect 165199 199880 165538 199882
rect 165199 199824 165204 199880
rect 165260 199824 165538 199880
rect 165199 199822 165538 199824
rect 165199 199819 165265 199822
rect 164006 199749 164066 199819
rect 159100 199686 159466 199746
rect 159100 199684 159106 199686
rect 159766 199684 159772 199748
rect 159836 199746 159842 199748
rect 160093 199746 160159 199749
rect 160369 199748 160435 199749
rect 160318 199746 160324 199748
rect 159836 199744 160159 199746
rect 159836 199688 160098 199744
rect 160154 199688 160159 199744
rect 159836 199686 160159 199688
rect 160278 199686 160324 199746
rect 160388 199744 160435 199748
rect 160430 199688 160435 199744
rect 159836 199684 159842 199686
rect 160093 199683 160159 199686
rect 160318 199684 160324 199686
rect 160388 199684 160435 199688
rect 162894 199684 162900 199748
rect 162964 199746 162970 199748
rect 163037 199746 163103 199749
rect 162964 199744 163103 199746
rect 162964 199688 163042 199744
rect 163098 199688 163103 199744
rect 162964 199686 163103 199688
rect 162964 199684 162970 199686
rect 160369 199683 160435 199684
rect 163037 199683 163103 199686
rect 163267 199746 163333 199749
rect 163814 199746 163820 199748
rect 163267 199744 163820 199746
rect 163267 199688 163272 199744
rect 163328 199688 163820 199744
rect 163267 199686 163820 199688
rect 163267 199683 163333 199686
rect 163814 199684 163820 199686
rect 163884 199684 163890 199748
rect 163957 199744 164066 199749
rect 163957 199688 163962 199744
rect 164018 199688 164066 199744
rect 163957 199686 164066 199688
rect 165478 199746 165538 199822
rect 165838 199820 165844 199884
rect 165908 199882 165914 199884
rect 165908 199822 165966 199882
rect 166395 199858 166400 199914
rect 166456 199858 166461 199914
rect 166628 199914 166737 199916
rect 166628 199884 166676 199914
rect 166395 199853 166461 199858
rect 165908 199820 165914 199822
rect 166398 199749 166458 199853
rect 166574 199820 166580 199884
rect 166644 199858 166676 199884
rect 166732 199858 166737 199914
rect 169020 199914 169129 199916
rect 166644 199853 166737 199858
rect 166947 199880 167013 199885
rect 166644 199822 166688 199853
rect 166947 199824 166952 199880
rect 167008 199824 167013 199880
rect 166644 199820 166650 199822
rect 166947 199819 167013 199824
rect 168235 199880 168301 199885
rect 168603 199884 168669 199885
rect 168598 199882 168604 199884
rect 168235 199824 168240 199880
rect 168296 199824 168301 199880
rect 168235 199819 168301 199824
rect 168512 199822 168604 199882
rect 168598 199820 168604 199822
rect 168668 199820 168674 199884
rect 168782 199820 168788 199884
rect 168852 199882 168858 199884
rect 169020 199882 169068 199914
rect 168852 199858 169068 199882
rect 169124 199858 169129 199914
rect 168852 199853 169129 199858
rect 169523 199880 169589 199885
rect 168852 199822 169080 199853
rect 169523 199824 169528 199880
rect 169584 199824 169589 199880
rect 168852 199820 168858 199822
rect 168603 199819 168669 199820
rect 169523 199819 169589 199824
rect 165613 199746 165679 199749
rect 165478 199744 165679 199746
rect 165478 199688 165618 199744
rect 165674 199688 165679 199744
rect 165478 199686 165679 199688
rect 163957 199683 164023 199686
rect 165613 199683 165679 199686
rect 166349 199744 166458 199749
rect 166809 199748 166875 199749
rect 166758 199746 166764 199748
rect 166349 199688 166354 199744
rect 166410 199688 166458 199744
rect 166349 199686 166458 199688
rect 166718 199686 166764 199746
rect 166828 199744 166875 199748
rect 166870 199688 166875 199744
rect 166349 199683 166415 199686
rect 166758 199684 166764 199686
rect 166828 199684 166875 199688
rect 166950 199746 167010 199819
rect 167085 199746 167151 199749
rect 166950 199744 167151 199746
rect 166950 199688 167090 199744
rect 167146 199688 167151 199744
rect 166950 199686 167151 199688
rect 166809 199683 166875 199684
rect 167085 199683 167151 199686
rect 167862 199684 167868 199748
rect 167932 199746 167938 199748
rect 168238 199746 168298 199819
rect 167932 199686 168298 199746
rect 167932 199684 167938 199686
rect 169150 199684 169156 199748
rect 169220 199746 169226 199748
rect 169526 199746 169586 199819
rect 169220 199686 169586 199746
rect 169220 199684 169226 199686
rect 169518 199610 169524 199612
rect 155174 199550 169524 199610
rect 153948 199548 153954 199550
rect 154021 199547 154087 199550
rect 169518 199548 169524 199550
rect 169588 199548 169594 199612
rect 169710 199610 169770 200094
rect 169886 200092 169892 200156
rect 169956 200154 169962 200156
rect 178861 200154 178927 200157
rect 201953 200154 202019 200157
rect 169956 200094 176210 200154
rect 169956 200092 169962 200094
rect 170806 200018 170812 200020
rect 170124 199958 170812 200018
rect 169983 199882 170049 199885
rect 170124 199882 170184 199958
rect 170806 199956 170812 199958
rect 170876 199956 170882 200020
rect 176150 200018 176210 200094
rect 178861 200152 202019 200154
rect 178861 200096 178866 200152
rect 178922 200096 201958 200152
rect 202014 200096 202019 200152
rect 178861 200094 202019 200096
rect 178861 200091 178927 200094
rect 201953 200091 202019 200094
rect 178350 200018 178356 200020
rect 176150 199958 178356 200018
rect 178350 199956 178356 199958
rect 178420 199956 178426 200020
rect 171363 199914 171429 199919
rect 170443 199884 170509 199885
rect 170438 199882 170444 199884
rect 169983 199880 170184 199882
rect 169983 199824 169988 199880
rect 170044 199824 170184 199880
rect 169983 199822 170184 199824
rect 170352 199822 170444 199882
rect 169983 199819 170049 199822
rect 170438 199820 170444 199822
rect 170508 199820 170514 199884
rect 170995 199882 171061 199885
rect 171363 199884 171368 199914
rect 171424 199884 171429 199914
rect 174307 199914 174373 199919
rect 170630 199880 171061 199882
rect 170630 199824 171000 199880
rect 171056 199824 171061 199880
rect 170630 199822 171061 199824
rect 170443 199819 170509 199820
rect 170070 199684 170076 199748
rect 170140 199746 170146 199748
rect 170630 199746 170690 199822
rect 170995 199819 171061 199822
rect 171358 199820 171364 199884
rect 171428 199882 171434 199884
rect 171639 199882 171705 199885
rect 171910 199882 171916 199884
rect 171428 199822 171486 199882
rect 171639 199880 171916 199882
rect 171639 199824 171644 199880
rect 171700 199824 171916 199880
rect 171639 199822 171916 199824
rect 171428 199820 171434 199822
rect 171639 199819 171705 199822
rect 171910 199820 171916 199822
rect 171980 199820 171986 199884
rect 172094 199820 172100 199884
rect 172164 199882 172170 199884
rect 172283 199882 172349 199885
rect 172164 199880 172349 199882
rect 172164 199824 172288 199880
rect 172344 199824 172349 199880
rect 172164 199822 172349 199824
rect 172164 199820 172170 199822
rect 172283 199819 172349 199822
rect 172646 199820 172652 199884
rect 172716 199882 172722 199884
rect 173755 199882 173821 199885
rect 172716 199880 173821 199882
rect 172716 199824 173760 199880
rect 173816 199824 173821 199880
rect 174307 199858 174312 199914
rect 174368 199858 174373 199914
rect 174307 199853 174373 199858
rect 172716 199822 173821 199824
rect 172716 199820 172722 199822
rect 173755 199819 173821 199822
rect 170140 199686 170690 199746
rect 170765 199748 170831 199749
rect 171041 199748 171107 199749
rect 172329 199748 172395 199749
rect 170765 199744 170812 199748
rect 170876 199746 170882 199748
rect 170765 199688 170770 199744
rect 170140 199684 170146 199686
rect 170765 199684 170812 199688
rect 170876 199686 170922 199746
rect 170876 199684 170882 199686
rect 170990 199684 170996 199748
rect 171060 199746 171107 199748
rect 172278 199746 172284 199748
rect 171060 199744 171152 199746
rect 171102 199688 171152 199744
rect 171060 199686 171152 199688
rect 172238 199686 172284 199746
rect 172348 199744 172395 199748
rect 172390 199688 172395 199744
rect 171060 199684 171107 199686
rect 172278 199684 172284 199686
rect 172348 199684 172395 199688
rect 174310 199746 174370 199853
rect 174486 199820 174492 199884
rect 174556 199882 174562 199884
rect 175135 199882 175201 199885
rect 174556 199880 175201 199882
rect 174556 199824 175140 199880
rect 175196 199824 175201 199880
rect 174556 199822 175201 199824
rect 174556 199820 174562 199822
rect 175135 199819 175201 199822
rect 175411 199882 175477 199885
rect 175871 199882 175937 199885
rect 176142 199882 176148 199884
rect 175411 199880 175520 199882
rect 175411 199824 175416 199880
rect 175472 199824 175520 199880
rect 175411 199819 175520 199824
rect 175871 199880 176148 199882
rect 175871 199824 175876 199880
rect 175932 199824 176148 199880
rect 175871 199822 176148 199824
rect 175871 199819 175937 199822
rect 176142 199820 176148 199822
rect 176212 199820 176218 199884
rect 176331 199880 176397 199885
rect 176331 199824 176336 199880
rect 176392 199824 176397 199880
rect 176331 199819 176397 199824
rect 176883 199880 176949 199885
rect 176883 199824 176888 199880
rect 176944 199824 176949 199880
rect 176883 199819 176949 199824
rect 177067 199882 177133 199885
rect 190361 199882 190427 199885
rect 177067 199880 190427 199882
rect 177067 199824 177072 199880
rect 177128 199824 190366 199880
rect 190422 199824 190427 199880
rect 177067 199822 190427 199824
rect 177067 199819 177133 199822
rect 190361 199819 190427 199822
rect 175460 199749 175520 199819
rect 176334 199749 176394 199819
rect 174486 199746 174492 199748
rect 174310 199686 174492 199746
rect 174486 199684 174492 199686
rect 174556 199684 174562 199748
rect 175457 199744 175523 199749
rect 175457 199688 175462 199744
rect 175518 199688 175523 199744
rect 170765 199683 170831 199684
rect 171041 199683 171107 199684
rect 172329 199683 172395 199684
rect 175457 199683 175523 199688
rect 175590 199684 175596 199748
rect 175660 199746 175666 199748
rect 175917 199746 175983 199749
rect 175660 199744 175983 199746
rect 175660 199688 175922 199744
rect 175978 199688 175983 199744
rect 175660 199686 175983 199688
rect 175660 199684 175666 199686
rect 175917 199683 175983 199686
rect 176285 199744 176394 199749
rect 176285 199688 176290 199744
rect 176346 199688 176394 199744
rect 176285 199686 176394 199688
rect 176886 199746 176946 199819
rect 200614 199746 200620 199748
rect 176886 199686 200620 199746
rect 176285 199683 176351 199686
rect 200614 199684 200620 199686
rect 200684 199684 200690 199748
rect 180926 199610 180932 199612
rect 169710 199550 180932 199610
rect 180926 199548 180932 199550
rect 180996 199548 181002 199612
rect 154665 199476 154731 199477
rect 154614 199474 154620 199476
rect 145741 199472 146218 199474
rect 145741 199416 145746 199472
rect 145802 199416 146218 199472
rect 145741 199414 146218 199416
rect 154574 199414 154620 199474
rect 154684 199472 154731 199476
rect 154726 199416 154731 199472
rect 139044 199412 139050 199414
rect 138841 199411 138907 199412
rect 145741 199411 145807 199414
rect 154614 199412 154620 199414
rect 154684 199412 154731 199416
rect 154665 199411 154731 199412
rect 155677 199474 155743 199477
rect 156270 199474 156276 199476
rect 155677 199472 156276 199474
rect 155677 199416 155682 199472
rect 155738 199416 156276 199472
rect 155677 199414 156276 199416
rect 155677 199411 155743 199414
rect 156270 199412 156276 199414
rect 156340 199412 156346 199476
rect 156454 199412 156460 199476
rect 156524 199474 156530 199476
rect 157149 199474 157215 199477
rect 156524 199472 157215 199474
rect 156524 199416 157154 199472
rect 157210 199416 157215 199472
rect 156524 199414 157215 199416
rect 156524 199412 156530 199414
rect 157149 199411 157215 199414
rect 158846 199412 158852 199476
rect 158916 199474 158922 199476
rect 159357 199474 159423 199477
rect 158916 199472 159423 199474
rect 158916 199416 159362 199472
rect 159418 199416 159423 199472
rect 158916 199414 159423 199416
rect 158916 199412 158922 199414
rect 159357 199411 159423 199414
rect 161197 199474 161263 199477
rect 162945 199476 163011 199477
rect 161422 199474 161428 199476
rect 161197 199472 161428 199474
rect 161197 199416 161202 199472
rect 161258 199416 161428 199472
rect 161197 199414 161428 199416
rect 161197 199411 161263 199414
rect 161422 199412 161428 199414
rect 161492 199412 161498 199476
rect 162894 199412 162900 199476
rect 162964 199474 163011 199476
rect 163221 199476 163287 199477
rect 163221 199474 163268 199476
rect 162964 199472 163056 199474
rect 163006 199416 163056 199472
rect 162964 199414 163056 199416
rect 163176 199472 163268 199474
rect 163176 199416 163226 199472
rect 163176 199414 163268 199416
rect 162964 199412 163011 199414
rect 162945 199411 163011 199412
rect 163221 199412 163268 199414
rect 163332 199412 163338 199476
rect 169569 199474 169635 199477
rect 169753 199474 169819 199477
rect 169569 199472 169819 199474
rect 169569 199416 169574 199472
rect 169630 199416 169758 199472
rect 169814 199416 169819 199472
rect 169569 199414 169819 199416
rect 163221 199411 163287 199412
rect 169569 199411 169635 199414
rect 169753 199411 169819 199414
rect 169886 199412 169892 199476
rect 169956 199474 169962 199476
rect 170121 199474 170187 199477
rect 170397 199476 170463 199477
rect 170397 199474 170444 199476
rect 169956 199472 170187 199474
rect 169956 199416 170126 199472
rect 170182 199416 170187 199472
rect 169956 199414 170187 199416
rect 170352 199472 170444 199474
rect 170352 199416 170402 199472
rect 170352 199414 170444 199416
rect 169956 199412 169962 199414
rect 170121 199411 170187 199414
rect 170397 199412 170444 199414
rect 170508 199412 170514 199476
rect 170765 199474 170831 199477
rect 170990 199474 170996 199476
rect 170765 199472 170996 199474
rect 170765 199416 170770 199472
rect 170826 199416 170996 199472
rect 170765 199414 170996 199416
rect 170397 199411 170463 199412
rect 170765 199411 170831 199414
rect 170990 199412 170996 199414
rect 171060 199412 171066 199476
rect 171358 199412 171364 199476
rect 171428 199474 171434 199476
rect 172237 199474 172303 199477
rect 171428 199472 172303 199474
rect 171428 199416 172242 199472
rect 172298 199416 172303 199472
rect 171428 199414 172303 199416
rect 171428 199412 171434 199414
rect 172237 199411 172303 199414
rect 172421 199474 172487 199477
rect 172789 199474 172855 199477
rect 173801 199476 173867 199477
rect 173750 199474 173756 199476
rect 172421 199472 172855 199474
rect 172421 199416 172426 199472
rect 172482 199416 172794 199472
rect 172850 199416 172855 199472
rect 172421 199414 172855 199416
rect 173710 199414 173756 199474
rect 173820 199472 173867 199476
rect 173862 199416 173867 199472
rect 172421 199411 172487 199414
rect 172789 199411 172855 199414
rect 173750 199412 173756 199414
rect 173820 199412 173867 199416
rect 173801 199411 173867 199412
rect 133137 199340 133203 199341
rect 133086 199338 133092 199340
rect 133046 199278 133092 199338
rect 133156 199336 133203 199340
rect 133198 199280 133203 199336
rect 133086 199276 133092 199278
rect 133156 199276 133203 199280
rect 139158 199276 139164 199340
rect 139228 199338 139234 199340
rect 139301 199338 139367 199341
rect 140313 199338 140379 199341
rect 139228 199336 139367 199338
rect 139228 199280 139306 199336
rect 139362 199280 139367 199336
rect 139228 199278 139367 199280
rect 139228 199276 139234 199278
rect 133137 199275 133203 199276
rect 139301 199275 139367 199278
rect 139902 199336 140379 199338
rect 139902 199280 140318 199336
rect 140374 199280 140379 199336
rect 139902 199278 140379 199280
rect 108941 199202 109007 199205
rect 136633 199202 136699 199205
rect 108941 199200 136699 199202
rect 108941 199144 108946 199200
rect 109002 199144 136638 199200
rect 136694 199144 136699 199200
rect 108941 199142 136699 199144
rect 108941 199139 109007 199142
rect 136633 199139 136699 199142
rect 136909 199202 136975 199205
rect 139669 199202 139735 199205
rect 136909 199200 139735 199202
rect 136909 199144 136914 199200
rect 136970 199144 139674 199200
rect 139730 199144 139735 199200
rect 136909 199142 139735 199144
rect 136909 199139 136975 199142
rect 139669 199139 139735 199142
rect 129641 199066 129707 199069
rect 133137 199066 133203 199069
rect 129641 199064 133203 199066
rect 129641 199008 129646 199064
rect 129702 199008 133142 199064
rect 133198 199008 133203 199064
rect 129641 199006 133203 199008
rect 129641 199003 129707 199006
rect 133137 199003 133203 199006
rect 137921 199066 137987 199069
rect 139209 199066 139275 199069
rect 137921 199064 139275 199066
rect 137921 199008 137926 199064
rect 137982 199008 139214 199064
rect 139270 199008 139275 199064
rect 137921 199006 139275 199008
rect 137921 199003 137987 199006
rect 139209 199003 139275 199006
rect 130193 198930 130259 198933
rect 136173 198930 136239 198933
rect 130193 198928 136239 198930
rect 130193 198872 130198 198928
rect 130254 198872 136178 198928
rect 136234 198872 136239 198928
rect 130193 198870 136239 198872
rect 130193 198867 130259 198870
rect 136173 198867 136239 198870
rect 136817 198930 136883 198933
rect 137502 198930 137508 198932
rect 136817 198928 137508 198930
rect 136817 198872 136822 198928
rect 136878 198872 137508 198928
rect 136817 198870 137508 198872
rect 136817 198867 136883 198870
rect 137502 198868 137508 198870
rect 137572 198868 137578 198932
rect 139902 198930 139962 199278
rect 140313 199275 140379 199278
rect 140589 199340 140655 199341
rect 140589 199336 140636 199340
rect 140700 199338 140706 199340
rect 140589 199280 140594 199336
rect 140589 199276 140636 199280
rect 140700 199278 140746 199338
rect 140700 199276 140706 199278
rect 141918 199276 141924 199340
rect 141988 199338 141994 199340
rect 153745 199338 153811 199341
rect 156873 199340 156939 199341
rect 141988 199336 153811 199338
rect 141988 199280 153750 199336
rect 153806 199280 153811 199336
rect 141988 199278 153811 199280
rect 141988 199276 141994 199278
rect 140589 199275 140655 199276
rect 153745 199275 153811 199278
rect 156822 199276 156828 199340
rect 156892 199338 156939 199340
rect 157149 199338 157215 199341
rect 182582 199338 182588 199340
rect 156892 199336 156984 199338
rect 156934 199280 156984 199336
rect 156892 199278 156984 199280
rect 157149 199336 182588 199338
rect 157149 199280 157154 199336
rect 157210 199280 182588 199336
rect 157149 199278 182588 199280
rect 156892 199276 156939 199278
rect 156873 199275 156939 199276
rect 157149 199275 157215 199278
rect 182582 199276 182588 199278
rect 182652 199276 182658 199340
rect 140313 199202 140379 199205
rect 140446 199202 140452 199204
rect 140313 199200 140452 199202
rect 140313 199144 140318 199200
rect 140374 199144 140452 199200
rect 140313 199142 140452 199144
rect 140313 199139 140379 199142
rect 140446 199140 140452 199142
rect 140516 199140 140522 199204
rect 152457 199202 152523 199205
rect 183502 199202 183508 199204
rect 152457 199200 183508 199202
rect 152457 199144 152462 199200
rect 152518 199144 183508 199200
rect 152457 199142 183508 199144
rect 152457 199139 152523 199142
rect 183502 199140 183508 199142
rect 183572 199140 183578 199204
rect 140037 199066 140103 199069
rect 140221 199066 140287 199069
rect 140037 199064 140287 199066
rect 140037 199008 140042 199064
rect 140098 199008 140226 199064
rect 140282 199008 140287 199064
rect 140037 199006 140287 199008
rect 140037 199003 140103 199006
rect 140221 199003 140287 199006
rect 146201 199066 146267 199069
rect 178166 199066 178172 199068
rect 146201 199064 178172 199066
rect 146201 199008 146206 199064
rect 146262 199008 178172 199064
rect 146201 199006 178172 199008
rect 146201 199003 146267 199006
rect 178166 199004 178172 199006
rect 178236 199004 178242 199068
rect 140221 198930 140287 198933
rect 183686 198930 183692 198932
rect 139902 198928 140287 198930
rect 139902 198872 140226 198928
rect 140282 198872 140287 198928
rect 139902 198870 140287 198872
rect 140221 198867 140287 198870
rect 150390 198870 183692 198930
rect 131481 198794 131547 198797
rect 138657 198794 138723 198797
rect 131481 198792 138723 198794
rect 131481 198736 131486 198792
rect 131542 198736 138662 198792
rect 138718 198736 138723 198792
rect 131481 198734 138723 198736
rect 131481 198731 131547 198734
rect 138657 198731 138723 198734
rect 148174 198732 148180 198796
rect 148244 198794 148250 198796
rect 148869 198794 148935 198797
rect 148244 198792 148935 198794
rect 148244 198736 148874 198792
rect 148930 198736 148935 198792
rect 148244 198734 148935 198736
rect 148244 198732 148250 198734
rect 148869 198731 148935 198734
rect 149329 198794 149395 198797
rect 150390 198794 150450 198870
rect 183686 198868 183692 198870
rect 183756 198868 183762 198932
rect 155953 198796 156019 198797
rect 149329 198792 150450 198794
rect 149329 198736 149334 198792
rect 149390 198736 150450 198792
rect 149329 198734 150450 198736
rect 149329 198731 149395 198734
rect 155902 198732 155908 198796
rect 155972 198794 156019 198796
rect 156137 198794 156203 198797
rect 184974 198794 184980 198796
rect 155972 198792 156064 198794
rect 156014 198736 156064 198792
rect 155972 198734 156064 198736
rect 156137 198792 184980 198794
rect 156137 198736 156142 198792
rect 156198 198736 184980 198792
rect 156137 198734 184980 198736
rect 155972 198732 156019 198734
rect 155953 198731 156019 198732
rect 156137 198731 156203 198734
rect 184974 198732 184980 198734
rect 185044 198732 185050 198796
rect 167494 198596 167500 198660
rect 167564 198658 167570 198660
rect 167637 198658 167703 198661
rect 167564 198656 167703 198658
rect 167564 198600 167642 198656
rect 167698 198600 167703 198656
rect 167564 198598 167703 198600
rect 167564 198596 167570 198598
rect 167637 198595 167703 198598
rect 171501 198658 171567 198661
rect 171726 198658 171732 198660
rect 171501 198656 171732 198658
rect 171501 198600 171506 198656
rect 171562 198600 171732 198656
rect 171501 198598 171732 198600
rect 171501 198595 171567 198598
rect 171726 198596 171732 198598
rect 171796 198596 171802 198660
rect 171910 198596 171916 198660
rect 171980 198658 171986 198660
rect 189206 198658 189212 198660
rect 171980 198598 189212 198658
rect 171980 198596 171986 198598
rect 189206 198596 189212 198598
rect 189276 198596 189282 198660
rect 195973 198658 196039 198661
rect 196566 198658 196572 198660
rect 195973 198656 196572 198658
rect 195973 198600 195978 198656
rect 196034 198600 196572 198656
rect 195973 198598 196572 198600
rect 195973 198595 196039 198598
rect 196566 198596 196572 198598
rect 196636 198596 196642 198660
rect 133597 198524 133663 198525
rect 133597 198520 133644 198524
rect 133708 198522 133714 198524
rect 133597 198464 133602 198520
rect 133597 198460 133644 198464
rect 133708 198462 133754 198522
rect 133708 198460 133714 198462
rect 153694 198460 153700 198524
rect 153764 198522 153770 198524
rect 158989 198522 159055 198525
rect 153764 198520 159055 198522
rect 153764 198464 158994 198520
rect 159050 198464 159055 198520
rect 153764 198462 159055 198464
rect 153764 198460 153770 198462
rect 133597 198459 133663 198460
rect 158989 198459 159055 198462
rect 169661 198522 169727 198525
rect 186998 198522 187004 198524
rect 169661 198520 187004 198522
rect 169661 198464 169666 198520
rect 169722 198464 187004 198520
rect 169661 198462 187004 198464
rect 169661 198459 169727 198462
rect 186998 198460 187004 198462
rect 187068 198460 187074 198524
rect 126830 198324 126836 198388
rect 126900 198386 126906 198388
rect 139209 198386 139275 198389
rect 126900 198384 139275 198386
rect 126900 198328 139214 198384
rect 139270 198328 139275 198384
rect 126900 198326 139275 198328
rect 126900 198324 126906 198326
rect 139209 198323 139275 198326
rect 156270 198324 156276 198388
rect 156340 198386 156346 198388
rect 156781 198386 156847 198389
rect 156340 198384 156847 198386
rect 156340 198328 156786 198384
rect 156842 198328 156847 198384
rect 156340 198326 156847 198328
rect 156340 198324 156346 198326
rect 156781 198323 156847 198326
rect 159766 198324 159772 198388
rect 159836 198386 159842 198388
rect 162301 198386 162367 198389
rect 159836 198384 162367 198386
rect 159836 198328 162306 198384
rect 162362 198328 162367 198384
rect 159836 198326 162367 198328
rect 159836 198324 159842 198326
rect 162301 198323 162367 198326
rect 170857 198386 170923 198389
rect 190494 198386 190500 198388
rect 170857 198384 190500 198386
rect 170857 198328 170862 198384
rect 170918 198328 190500 198384
rect 170857 198326 190500 198328
rect 170857 198323 170923 198326
rect 190494 198324 190500 198326
rect 190564 198324 190570 198388
rect 145373 198250 145439 198253
rect 142110 198248 145439 198250
rect 142110 198192 145378 198248
rect 145434 198192 145439 198248
rect 142110 198190 145439 198192
rect 125358 198052 125364 198116
rect 125428 198114 125434 198116
rect 142110 198114 142170 198190
rect 145373 198187 145439 198190
rect 163589 198252 163655 198253
rect 163589 198248 163636 198252
rect 163700 198250 163706 198252
rect 181437 198250 181503 198253
rect 194542 198250 194548 198252
rect 163589 198192 163594 198248
rect 163589 198188 163636 198192
rect 163700 198190 163746 198250
rect 167318 198190 176026 198250
rect 163700 198188 163706 198190
rect 163589 198187 163655 198188
rect 125428 198054 138674 198114
rect 125428 198052 125434 198054
rect 126646 197916 126652 197980
rect 126716 197978 126722 197980
rect 126716 197918 138306 197978
rect 126716 197916 126722 197918
rect 138246 197570 138306 197918
rect 138614 197842 138674 198054
rect 141926 198054 142170 198114
rect 157425 198114 157491 198117
rect 167085 198114 167151 198117
rect 157425 198112 167151 198114
rect 157425 198056 157430 198112
rect 157486 198056 167090 198112
rect 167146 198056 167151 198112
rect 157425 198054 167151 198056
rect 141926 197978 141986 198054
rect 157425 198051 157491 198054
rect 167085 198051 167151 198054
rect 140638 197918 141986 197978
rect 146477 197978 146543 197981
rect 167318 197978 167378 198190
rect 169518 198052 169524 198116
rect 169588 198114 169594 198116
rect 169753 198114 169819 198117
rect 169588 198112 169819 198114
rect 169588 198056 169758 198112
rect 169814 198056 169819 198112
rect 169588 198054 169819 198056
rect 169588 198052 169594 198054
rect 169753 198051 169819 198054
rect 171869 198116 171935 198117
rect 171869 198112 171916 198116
rect 171980 198114 171986 198116
rect 171869 198056 171874 198112
rect 171869 198052 171916 198056
rect 171980 198054 172026 198114
rect 171980 198052 171986 198054
rect 174118 198052 174124 198116
rect 174188 198114 174194 198116
rect 174905 198114 174971 198117
rect 174188 198112 174971 198114
rect 174188 198056 174910 198112
rect 174966 198056 174971 198112
rect 174188 198054 174971 198056
rect 175966 198114 176026 198190
rect 181437 198248 194548 198250
rect 181437 198192 181442 198248
rect 181498 198192 194548 198248
rect 181437 198190 194548 198192
rect 181437 198187 181503 198190
rect 194542 198188 194548 198190
rect 194612 198188 194618 198252
rect 176745 198114 176811 198117
rect 175966 198112 176811 198114
rect 175966 198056 176750 198112
rect 176806 198056 176811 198112
rect 175966 198054 176811 198056
rect 174188 198052 174194 198054
rect 171869 198051 171935 198052
rect 174905 198051 174971 198054
rect 176745 198051 176811 198054
rect 146477 197976 167378 197978
rect 146477 197920 146482 197976
rect 146538 197920 167378 197976
rect 146477 197918 167378 197920
rect 140638 197842 140698 197918
rect 146477 197915 146543 197918
rect 179454 197842 179460 197844
rect 138614 197782 140698 197842
rect 176150 197782 179460 197842
rect 139209 197706 139275 197709
rect 145281 197706 145347 197709
rect 139209 197704 145347 197706
rect 139209 197648 139214 197704
rect 139270 197648 145286 197704
rect 145342 197648 145347 197704
rect 139209 197646 145347 197648
rect 139209 197643 139275 197646
rect 145281 197643 145347 197646
rect 145598 197644 145604 197708
rect 145668 197706 145674 197708
rect 147765 197706 147831 197709
rect 145668 197704 147831 197706
rect 145668 197648 147770 197704
rect 147826 197648 147831 197704
rect 145668 197646 147831 197648
rect 145668 197644 145674 197646
rect 147765 197643 147831 197646
rect 167085 197706 167151 197709
rect 176150 197706 176210 197782
rect 179454 197780 179460 197782
rect 179524 197780 179530 197844
rect 167085 197704 176210 197706
rect 167085 197648 167090 197704
rect 167146 197648 176210 197704
rect 167085 197646 176210 197648
rect 167085 197643 167151 197646
rect 146569 197570 146635 197573
rect 138246 197568 146635 197570
rect 138246 197512 146574 197568
rect 146630 197512 146635 197568
rect 138246 197510 146635 197512
rect 146569 197507 146635 197510
rect 176745 197570 176811 197573
rect 179638 197570 179644 197572
rect 176745 197568 179644 197570
rect 176745 197512 176750 197568
rect 176806 197512 179644 197568
rect 176745 197510 179644 197512
rect 176745 197507 176811 197510
rect 179638 197508 179644 197510
rect 179708 197508 179714 197572
rect 132769 197434 132835 197437
rect 133454 197434 133460 197436
rect 132769 197432 133460 197434
rect 132769 197376 132774 197432
rect 132830 197376 133460 197432
rect 132769 197374 133460 197376
rect 132769 197371 132835 197374
rect 133454 197372 133460 197374
rect 133524 197372 133530 197436
rect 134190 197372 134196 197436
rect 134260 197434 134266 197436
rect 135161 197434 135227 197437
rect 134260 197432 135227 197434
rect 134260 197376 135166 197432
rect 135222 197376 135227 197432
rect 134260 197374 135227 197376
rect 134260 197372 134266 197374
rect 135161 197371 135227 197374
rect 140037 197436 140103 197437
rect 156597 197436 156663 197437
rect 140037 197432 140084 197436
rect 140148 197434 140154 197436
rect 140037 197376 140042 197432
rect 140037 197372 140084 197376
rect 140148 197374 140194 197434
rect 156597 197432 156644 197436
rect 156708 197434 156714 197436
rect 156597 197376 156602 197432
rect 140148 197372 140154 197374
rect 156597 197372 156644 197376
rect 156708 197374 156754 197434
rect 156708 197372 156714 197374
rect 140037 197371 140103 197372
rect 156597 197371 156663 197372
rect 129181 197298 129247 197301
rect 153285 197298 153351 197301
rect 129181 197296 153351 197298
rect 129181 197240 129186 197296
rect 129242 197240 153290 197296
rect 153346 197240 153351 197296
rect 129181 197238 153351 197240
rect 129181 197235 129247 197238
rect 153285 197235 153351 197238
rect 153561 197298 153627 197301
rect 154062 197298 154068 197300
rect 153561 197296 154068 197298
rect 153561 197240 153566 197296
rect 153622 197240 154068 197296
rect 153561 197238 154068 197240
rect 153561 197235 153627 197238
rect 154062 197236 154068 197238
rect 154132 197236 154138 197300
rect 166022 197236 166028 197300
rect 166092 197298 166098 197300
rect 166533 197298 166599 197301
rect 166092 197296 166599 197298
rect 166092 197240 166538 197296
rect 166594 197240 166599 197296
rect 166092 197238 166599 197240
rect 166092 197236 166098 197238
rect 166533 197235 166599 197238
rect 130469 197162 130535 197165
rect 154665 197162 154731 197165
rect 130469 197160 154731 197162
rect 130469 197104 130474 197160
rect 130530 197104 154670 197160
rect 154726 197104 154731 197160
rect 130469 197102 154731 197104
rect 130469 197099 130535 197102
rect 154665 197099 154731 197102
rect 165838 197100 165844 197164
rect 165908 197162 165914 197164
rect 183001 197162 183067 197165
rect 165908 197160 183067 197162
rect 165908 197104 183006 197160
rect 183062 197104 183067 197160
rect 165908 197102 183067 197104
rect 165908 197100 165914 197102
rect 183001 197099 183067 197102
rect 108205 197026 108271 197029
rect 137829 197026 137895 197029
rect 108205 197024 137895 197026
rect 108205 196968 108210 197024
rect 108266 196968 137834 197024
rect 137890 196968 137895 197024
rect 108205 196966 137895 196968
rect 108205 196963 108271 196966
rect 137829 196963 137895 196966
rect 161238 196964 161244 197028
rect 161308 197026 161314 197028
rect 169845 197026 169911 197029
rect 161308 197024 169911 197026
rect 161308 196968 169850 197024
rect 169906 196968 169911 197024
rect 161308 196966 169911 196968
rect 161308 196964 161314 196966
rect 169845 196963 169911 196966
rect 176285 197026 176351 197029
rect 197302 197026 197308 197028
rect 176285 197024 197308 197026
rect 176285 196968 176290 197024
rect 176346 196968 197308 197024
rect 176285 196966 197308 196968
rect 176285 196963 176351 196966
rect 197302 196964 197308 196966
rect 197372 196964 197378 197028
rect 104433 196890 104499 196893
rect 134609 196890 134675 196893
rect 104433 196888 134675 196890
rect 104433 196832 104438 196888
rect 104494 196832 134614 196888
rect 134670 196832 134675 196888
rect 104433 196830 134675 196832
rect 104433 196827 104499 196830
rect 134609 196827 134675 196830
rect 163078 196828 163084 196892
rect 163148 196890 163154 196892
rect 171777 196890 171843 196893
rect 163148 196888 171843 196890
rect 163148 196832 171782 196888
rect 171838 196832 171843 196888
rect 163148 196830 171843 196832
rect 163148 196828 163154 196830
rect 171777 196827 171843 196830
rect 108481 196754 108547 196757
rect 138473 196754 138539 196757
rect 108481 196752 138539 196754
rect 108481 196696 108486 196752
rect 108542 196696 138478 196752
rect 138534 196696 138539 196752
rect 108481 196694 138539 196696
rect 108481 196691 108547 196694
rect 138473 196691 138539 196694
rect 169569 196754 169635 196757
rect 203149 196754 203215 196757
rect 169569 196752 203215 196754
rect 169569 196696 169574 196752
rect 169630 196696 203154 196752
rect 203210 196696 203215 196752
rect 169569 196694 203215 196696
rect 169569 196691 169635 196694
rect 203149 196691 203215 196694
rect 107101 196618 107167 196621
rect 138197 196618 138263 196621
rect 107101 196616 138263 196618
rect 107101 196560 107106 196616
rect 107162 196560 138202 196616
rect 138258 196560 138263 196616
rect 107101 196558 138263 196560
rect 107101 196555 107167 196558
rect 138197 196555 138263 196558
rect 164969 196618 165035 196621
rect 198917 196618 198983 196621
rect 164969 196616 198983 196618
rect 164969 196560 164974 196616
rect 165030 196560 198922 196616
rect 198978 196560 198983 196616
rect 164969 196558 198983 196560
rect 164969 196555 165035 196558
rect 198917 196555 198983 196558
rect 174629 196484 174695 196485
rect 174629 196480 174676 196484
rect 174740 196482 174746 196484
rect 174629 196424 174634 196480
rect 174629 196420 174676 196424
rect 174740 196422 174786 196482
rect 174740 196420 174746 196422
rect 174629 196419 174695 196420
rect 135846 196284 135852 196348
rect 135916 196346 135922 196348
rect 136173 196346 136239 196349
rect 135916 196344 136239 196346
rect 135916 196288 136178 196344
rect 136234 196288 136239 196344
rect 135916 196286 136239 196288
rect 135916 196284 135922 196286
rect 136173 196283 136239 196286
rect 135846 196148 135852 196212
rect 135916 196210 135922 196212
rect 135989 196210 136055 196213
rect 135916 196208 136055 196210
rect 135916 196152 135994 196208
rect 136050 196152 136055 196208
rect 135916 196150 136055 196152
rect 135916 196148 135922 196150
rect 135989 196147 136055 196150
rect 122557 196074 122623 196077
rect 136265 196076 136331 196077
rect 139209 196076 139275 196077
rect 122782 196074 122788 196076
rect 122557 196072 122788 196074
rect 122557 196016 122562 196072
rect 122618 196016 122788 196072
rect 122557 196014 122788 196016
rect 122557 196011 122623 196014
rect 122782 196012 122788 196014
rect 122852 196012 122858 196076
rect 136214 196012 136220 196076
rect 136284 196074 136331 196076
rect 136284 196072 136376 196074
rect 136326 196016 136376 196072
rect 136284 196014 136376 196016
rect 136284 196012 136331 196014
rect 139158 196012 139164 196076
rect 139228 196074 139275 196076
rect 149053 196074 149119 196077
rect 158662 196074 158668 196076
rect 139228 196072 139320 196074
rect 139270 196016 139320 196072
rect 139228 196014 139320 196016
rect 149053 196072 158668 196074
rect 149053 196016 149058 196072
rect 149114 196016 158668 196072
rect 149053 196014 158668 196016
rect 139228 196012 139275 196014
rect 136265 196011 136331 196012
rect 139209 196011 139275 196012
rect 149053 196011 149119 196014
rect 158662 196012 158668 196014
rect 158732 196012 158738 196076
rect 117681 195938 117747 195941
rect 138013 195938 138079 195941
rect 151537 195940 151603 195941
rect 151486 195938 151492 195940
rect 117681 195936 138079 195938
rect 117681 195880 117686 195936
rect 117742 195880 138018 195936
rect 138074 195880 138079 195936
rect 117681 195878 138079 195880
rect 151446 195878 151492 195938
rect 151556 195936 151603 195940
rect 151598 195880 151603 195936
rect 117681 195875 117747 195878
rect 138013 195875 138079 195878
rect 151486 195876 151492 195878
rect 151556 195876 151603 195880
rect 151537 195875 151603 195876
rect 155861 195938 155927 195941
rect 160277 195940 160343 195941
rect 156086 195938 156092 195940
rect 155861 195936 156092 195938
rect 155861 195880 155866 195936
rect 155922 195880 156092 195936
rect 155861 195878 156092 195880
rect 155861 195875 155927 195878
rect 156086 195876 156092 195878
rect 156156 195876 156162 195940
rect 160277 195938 160324 195940
rect 160232 195936 160324 195938
rect 160232 195880 160282 195936
rect 160232 195878 160324 195880
rect 160277 195876 160324 195878
rect 160388 195876 160394 195940
rect 162710 195876 162716 195940
rect 162780 195938 162786 195940
rect 163037 195938 163103 195941
rect 162780 195936 163103 195938
rect 162780 195880 163042 195936
rect 163098 195880 163103 195936
rect 162780 195878 163103 195880
rect 162780 195876 162786 195878
rect 160277 195875 160343 195876
rect 163037 195875 163103 195878
rect 131982 195740 131988 195804
rect 132052 195802 132058 195804
rect 149237 195802 149303 195805
rect 132052 195800 149303 195802
rect 132052 195744 149242 195800
rect 149298 195744 149303 195800
rect 132052 195742 149303 195744
rect 132052 195740 132058 195742
rect 149237 195739 149303 195742
rect 128118 195604 128124 195668
rect 128188 195666 128194 195668
rect 146937 195666 147003 195669
rect 128188 195664 147003 195666
rect 128188 195608 146942 195664
rect 146998 195608 147003 195664
rect 128188 195606 147003 195608
rect 128188 195604 128194 195606
rect 146937 195603 147003 195606
rect 175273 195666 175339 195669
rect 187182 195666 187188 195668
rect 175273 195664 187188 195666
rect 175273 195608 175278 195664
rect 175334 195608 187188 195664
rect 175273 195606 187188 195608
rect 175273 195603 175339 195606
rect 187182 195604 187188 195606
rect 187252 195604 187258 195668
rect 127934 195468 127940 195532
rect 128004 195530 128010 195532
rect 148041 195530 148107 195533
rect 149697 195532 149763 195533
rect 128004 195528 148107 195530
rect 128004 195472 148046 195528
rect 148102 195472 148107 195528
rect 128004 195470 148107 195472
rect 128004 195468 128010 195470
rect 148041 195467 148107 195470
rect 149646 195468 149652 195532
rect 149716 195530 149763 195532
rect 149973 195532 150039 195533
rect 149973 195530 150020 195532
rect 149716 195528 149808 195530
rect 149758 195472 149808 195528
rect 149716 195470 149808 195472
rect 149928 195528 150020 195530
rect 149928 195472 149978 195528
rect 149928 195470 150020 195472
rect 149716 195468 149763 195470
rect 149697 195467 149763 195468
rect 149973 195468 150020 195470
rect 150084 195468 150090 195532
rect 153878 195468 153884 195532
rect 153948 195530 153954 195532
rect 154389 195530 154455 195533
rect 153948 195528 154455 195530
rect 153948 195472 154394 195528
rect 154450 195472 154455 195528
rect 153948 195470 154455 195472
rect 153948 195468 153954 195470
rect 149973 195467 150039 195468
rect 154389 195467 154455 195470
rect 167361 195530 167427 195533
rect 168046 195530 168052 195532
rect 167361 195528 168052 195530
rect 167361 195472 167366 195528
rect 167422 195472 168052 195528
rect 167361 195470 168052 195472
rect 167361 195467 167427 195470
rect 168046 195468 168052 195470
rect 168116 195468 168122 195532
rect 168373 195530 168439 195533
rect 169150 195530 169156 195532
rect 168373 195528 169156 195530
rect 168373 195472 168378 195528
rect 168434 195472 169156 195528
rect 168373 195470 169156 195472
rect 168373 195467 168439 195470
rect 169150 195468 169156 195470
rect 169220 195468 169226 195532
rect 170673 195530 170739 195533
rect 172094 195530 172100 195532
rect 170673 195528 172100 195530
rect 170673 195472 170678 195528
rect 170734 195472 172100 195528
rect 170673 195470 172100 195472
rect 170673 195467 170739 195470
rect 172094 195468 172100 195470
rect 172164 195468 172170 195532
rect 174997 195530 175063 195533
rect 191782 195530 191788 195532
rect 174997 195528 191788 195530
rect 174997 195472 175002 195528
rect 175058 195472 191788 195528
rect 174997 195470 191788 195472
rect 174997 195467 175063 195470
rect 191782 195468 191788 195470
rect 191852 195468 191858 195532
rect 112437 195394 112503 195397
rect 142337 195394 142403 195397
rect 112437 195392 142403 195394
rect 112437 195336 112442 195392
rect 112498 195336 142342 195392
rect 142398 195336 142403 195392
rect 112437 195334 142403 195336
rect 112437 195331 112503 195334
rect 142337 195331 142403 195334
rect 145230 195332 145236 195396
rect 145300 195394 145306 195396
rect 162945 195394 163011 195397
rect 145300 195392 163011 195394
rect 145300 195336 162950 195392
rect 163006 195336 163011 195392
rect 145300 195334 163011 195336
rect 145300 195332 145306 195334
rect 162945 195331 163011 195334
rect 167678 195332 167684 195396
rect 167748 195394 167754 195396
rect 167913 195394 167979 195397
rect 167748 195392 167979 195394
rect 167748 195336 167918 195392
rect 167974 195336 167979 195392
rect 167748 195334 167979 195336
rect 167748 195332 167754 195334
rect 167913 195331 167979 195334
rect 168741 195394 168807 195397
rect 202965 195394 203031 195397
rect 168741 195392 203031 195394
rect 168741 195336 168746 195392
rect 168802 195336 202970 195392
rect 203026 195336 203031 195392
rect 168741 195334 203031 195336
rect 168741 195331 168807 195334
rect 202965 195331 203031 195334
rect 121310 195196 121316 195260
rect 121380 195258 121386 195260
rect 132033 195258 132099 195261
rect 121380 195256 132099 195258
rect 121380 195200 132038 195256
rect 132094 195200 132099 195256
rect 121380 195198 132099 195200
rect 121380 195196 121386 195198
rect 132033 195195 132099 195198
rect 132166 195196 132172 195260
rect 132236 195258 132242 195260
rect 148910 195258 148916 195260
rect 132236 195198 148916 195258
rect 132236 195196 132242 195198
rect 148910 195196 148916 195198
rect 148980 195196 148986 195260
rect 150709 195258 150775 195261
rect 151118 195258 151124 195260
rect 150709 195256 151124 195258
rect 150709 195200 150714 195256
rect 150770 195200 151124 195256
rect 150709 195198 151124 195200
rect 150709 195195 150775 195198
rect 151118 195196 151124 195198
rect 151188 195196 151194 195260
rect 153510 195196 153516 195260
rect 153580 195258 153586 195260
rect 153653 195258 153719 195261
rect 153580 195256 153719 195258
rect 153580 195200 153658 195256
rect 153714 195200 153719 195256
rect 153580 195198 153719 195200
rect 153580 195196 153586 195198
rect 153653 195195 153719 195198
rect 154297 195258 154363 195261
rect 154430 195258 154436 195260
rect 154297 195256 154436 195258
rect 154297 195200 154302 195256
rect 154358 195200 154436 195256
rect 154297 195198 154436 195200
rect 154297 195195 154363 195198
rect 154430 195196 154436 195198
rect 154500 195196 154506 195260
rect 162894 195196 162900 195260
rect 162964 195258 162970 195260
rect 164049 195258 164115 195261
rect 162964 195256 164115 195258
rect 162964 195200 164054 195256
rect 164110 195200 164115 195256
rect 162964 195198 164115 195200
rect 162964 195196 162970 195198
rect 164049 195195 164115 195198
rect 164693 195260 164759 195261
rect 164693 195256 164740 195260
rect 164804 195258 164810 195260
rect 164693 195200 164698 195256
rect 164693 195196 164740 195200
rect 164804 195198 164850 195258
rect 164804 195196 164810 195198
rect 166574 195196 166580 195260
rect 166644 195258 166650 195260
rect 200481 195258 200547 195261
rect 166644 195256 200547 195258
rect 166644 195200 200486 195256
rect 200542 195200 200547 195256
rect 166644 195198 200547 195200
rect 166644 195196 166650 195198
rect 164693 195195 164759 195196
rect 200481 195195 200547 195198
rect 130878 195060 130884 195124
rect 130948 195122 130954 195124
rect 143901 195122 143967 195125
rect 130948 195120 143967 195122
rect 130948 195064 143906 195120
rect 143962 195064 143967 195120
rect 130948 195062 143967 195064
rect 130948 195060 130954 195062
rect 143901 195059 143967 195062
rect 149646 195060 149652 195124
rect 149716 195122 149722 195124
rect 150341 195122 150407 195125
rect 149716 195120 150407 195122
rect 149716 195064 150346 195120
rect 150402 195064 150407 195120
rect 149716 195062 150407 195064
rect 149716 195060 149722 195062
rect 150341 195059 150407 195062
rect 152590 195060 152596 195124
rect 152660 195122 152666 195124
rect 161841 195122 161907 195125
rect 152660 195120 161907 195122
rect 152660 195064 161846 195120
rect 161902 195064 161907 195120
rect 152660 195062 161907 195064
rect 152660 195060 152666 195062
rect 161841 195059 161907 195062
rect 164366 195060 164372 195124
rect 164436 195122 164442 195124
rect 178309 195122 178375 195125
rect 164436 195120 178375 195122
rect 164436 195064 178314 195120
rect 178370 195064 178375 195120
rect 164436 195062 178375 195064
rect 164436 195060 164442 195062
rect 178309 195059 178375 195062
rect 136214 194924 136220 194988
rect 136284 194986 136290 194988
rect 136449 194986 136515 194989
rect 137185 194988 137251 194989
rect 136284 194984 136515 194986
rect 136284 194928 136454 194984
rect 136510 194928 136515 194984
rect 136284 194926 136515 194928
rect 136284 194924 136290 194926
rect 136449 194923 136515 194926
rect 137134 194924 137140 194988
rect 137204 194986 137251 194988
rect 137204 194984 137296 194986
rect 137246 194928 137296 194984
rect 137204 194926 137296 194928
rect 137204 194924 137251 194926
rect 138054 194924 138060 194988
rect 138124 194986 138130 194988
rect 138381 194986 138447 194989
rect 138124 194984 138447 194986
rect 138124 194928 138386 194984
rect 138442 194928 138447 194984
rect 138124 194926 138447 194928
rect 138124 194924 138130 194926
rect 137185 194923 137251 194924
rect 138381 194923 138447 194926
rect 139117 194988 139183 194989
rect 139117 194984 139164 194988
rect 139228 194986 139234 194988
rect 139117 194928 139122 194984
rect 139117 194924 139164 194928
rect 139228 194926 139274 194986
rect 139228 194924 139234 194926
rect 148726 194924 148732 194988
rect 148796 194986 148802 194988
rect 160645 194986 160711 194989
rect 164509 194988 164575 194989
rect 164509 194986 164556 194988
rect 148796 194984 160711 194986
rect 148796 194928 160650 194984
rect 160706 194928 160711 194984
rect 148796 194926 160711 194928
rect 164464 194984 164556 194986
rect 164464 194928 164514 194984
rect 164464 194926 164556 194928
rect 148796 194924 148802 194926
rect 139117 194923 139183 194924
rect 160645 194923 160711 194926
rect 164509 194924 164556 194926
rect 164620 194924 164626 194988
rect 165654 194924 165660 194988
rect 165724 194986 165730 194988
rect 189257 194986 189323 194989
rect 165724 194984 189323 194986
rect 165724 194928 189262 194984
rect 189318 194928 189323 194984
rect 165724 194926 189323 194928
rect 165724 194924 165730 194926
rect 164509 194923 164575 194924
rect 189257 194923 189323 194926
rect 138422 194788 138428 194852
rect 138492 194850 138498 194852
rect 138565 194850 138631 194853
rect 138492 194848 138631 194850
rect 138492 194792 138570 194848
rect 138626 194792 138631 194848
rect 138492 194790 138631 194792
rect 138492 194788 138498 194790
rect 138565 194787 138631 194790
rect 175406 194788 175412 194852
rect 175476 194850 175482 194852
rect 175641 194850 175707 194853
rect 175476 194848 175707 194850
rect 175476 194792 175646 194848
rect 175702 194792 175707 194848
rect 175476 194790 175707 194792
rect 175476 194788 175482 194790
rect 175641 194787 175707 194790
rect 186405 194850 186471 194853
rect 187366 194850 187372 194852
rect 186405 194848 187372 194850
rect 186405 194792 186410 194848
rect 186466 194792 187372 194848
rect 186405 194790 187372 194792
rect 186405 194787 186471 194790
rect 187366 194788 187372 194790
rect 187436 194788 187442 194852
rect 104617 194170 104683 194173
rect 133045 194170 133111 194173
rect 152273 194172 152339 194173
rect 152222 194170 152228 194172
rect 104617 194168 133111 194170
rect 104617 194112 104622 194168
rect 104678 194112 133050 194168
rect 133106 194112 133111 194168
rect 104617 194110 133111 194112
rect 152182 194110 152228 194170
rect 152292 194168 152339 194172
rect 152334 194112 152339 194168
rect 104617 194107 104683 194110
rect 133045 194107 133111 194110
rect 152222 194108 152228 194110
rect 152292 194108 152339 194112
rect 152273 194107 152339 194108
rect 124990 193972 124996 194036
rect 125060 194034 125066 194036
rect 145465 194034 145531 194037
rect 125060 194032 145531 194034
rect 125060 193976 145470 194032
rect 145526 193976 145531 194032
rect 125060 193974 145531 193976
rect 125060 193972 125066 193974
rect 145465 193971 145531 193974
rect 157977 194034 158043 194037
rect 158478 194034 158484 194036
rect 157977 194032 158484 194034
rect 157977 193976 157982 194032
rect 158038 193976 158484 194032
rect 157977 193974 158484 193976
rect 157977 193971 158043 193974
rect 158478 193972 158484 193974
rect 158548 193972 158554 194036
rect 100661 193898 100727 193901
rect 133270 193898 133276 193900
rect 100661 193896 133276 193898
rect 100661 193840 100666 193896
rect 100722 193840 133276 193896
rect 100661 193838 133276 193840
rect 100661 193835 100727 193838
rect 133270 193836 133276 193838
rect 133340 193836 133346 193900
rect 115197 192810 115263 192813
rect 142245 192810 142311 192813
rect 115197 192808 142311 192810
rect 115197 192752 115202 192808
rect 115258 192752 142250 192808
rect 142306 192752 142311 192808
rect 115197 192750 142311 192752
rect 115197 192747 115263 192750
rect 142245 192747 142311 192750
rect 106181 192674 106247 192677
rect 137277 192674 137343 192677
rect 106181 192672 137343 192674
rect 106181 192616 106186 192672
rect 106242 192616 137282 192672
rect 137338 192616 137343 192672
rect 106181 192614 137343 192616
rect 106181 192611 106247 192614
rect 137277 192611 137343 192614
rect 190361 192674 190427 192677
rect 204437 192674 204503 192677
rect 190361 192672 204503 192674
rect 190361 192616 190366 192672
rect 190422 192616 204442 192672
rect 204498 192616 204503 192672
rect 190361 192614 204503 192616
rect 190361 192611 190427 192614
rect 204437 192611 204503 192614
rect 103237 192538 103303 192541
rect 136725 192538 136791 192541
rect 103237 192536 136791 192538
rect 103237 192480 103242 192536
rect 103298 192480 136730 192536
rect 136786 192480 136791 192536
rect 103237 192478 136791 192480
rect 103237 192475 103303 192478
rect 136725 192475 136791 192478
rect 175457 192538 175523 192541
rect 205633 192538 205699 192541
rect 175457 192536 205699 192538
rect 175457 192480 175462 192536
rect 175518 192480 205638 192536
rect 205694 192480 205699 192536
rect 175457 192478 205699 192480
rect 175457 192475 175523 192478
rect 205633 192475 205699 192478
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 151854 191524 151860 191588
rect 151924 191586 151930 191588
rect 152089 191586 152155 191589
rect 151924 191584 152155 191586
rect 151924 191528 152094 191584
rect 152150 191528 152155 191584
rect 151924 191526 152155 191528
rect 151924 191524 151930 191526
rect 152089 191523 152155 191526
rect 148910 191388 148916 191452
rect 148980 191450 148986 191452
rect 160461 191450 160527 191453
rect 148980 191448 160527 191450
rect 148980 191392 160466 191448
rect 160522 191392 160527 191448
rect 148980 191390 160527 191392
rect 148980 191388 148986 191390
rect 160461 191387 160527 191390
rect 149462 191252 149468 191316
rect 149532 191314 149538 191316
rect 160185 191314 160251 191317
rect 149532 191312 160251 191314
rect 149532 191256 160190 191312
rect 160246 191256 160251 191312
rect 149532 191254 160251 191256
rect 149532 191252 149538 191254
rect 160185 191251 160251 191254
rect 173157 191314 173223 191317
rect 173382 191314 173388 191316
rect 173157 191312 173388 191314
rect 173157 191256 173162 191312
rect 173218 191256 173388 191312
rect 173157 191254 173388 191256
rect 173157 191251 173223 191254
rect 173382 191252 173388 191254
rect 173452 191252 173458 191316
rect 140998 191116 141004 191180
rect 141068 191178 141074 191180
rect 142061 191178 142127 191181
rect 141068 191176 142127 191178
rect 141068 191120 142066 191176
rect 142122 191120 142127 191176
rect 141068 191118 142127 191120
rect 141068 191116 141074 191118
rect 142061 191115 142127 191118
rect 145414 191116 145420 191180
rect 145484 191178 145490 191180
rect 146109 191178 146175 191181
rect 145484 191176 146175 191178
rect 145484 191120 146114 191176
rect 146170 191120 146175 191176
rect 145484 191118 146175 191120
rect 145484 191116 145490 191118
rect 146109 191115 146175 191118
rect 147070 191116 147076 191180
rect 147140 191178 147146 191180
rect 147213 191178 147279 191181
rect 147140 191176 147279 191178
rect 147140 191120 147218 191176
rect 147274 191120 147279 191176
rect 147140 191118 147279 191120
rect 147140 191116 147146 191118
rect 147213 191115 147279 191118
rect 150341 191178 150407 191181
rect 156086 191178 156092 191180
rect 150341 191176 156092 191178
rect 150341 191120 150346 191176
rect 150402 191120 156092 191176
rect 150341 191118 156092 191120
rect 150341 191115 150407 191118
rect 156086 191116 156092 191118
rect 156156 191116 156162 191180
rect 158110 191116 158116 191180
rect 158180 191178 158186 191180
rect 158529 191178 158595 191181
rect 158180 191176 158595 191178
rect 158180 191120 158534 191176
rect 158590 191120 158595 191176
rect 158180 191118 158595 191120
rect 158180 191116 158186 191118
rect 158529 191115 158595 191118
rect 160737 191178 160803 191181
rect 161054 191178 161060 191180
rect 160737 191176 161060 191178
rect 160737 191120 160742 191176
rect 160798 191120 161060 191176
rect 160737 191118 161060 191120
rect 160737 191115 160803 191118
rect 161054 191116 161060 191118
rect 161124 191116 161130 191180
rect 162158 191116 162164 191180
rect 162228 191178 162234 191180
rect 162669 191178 162735 191181
rect 162228 191176 162735 191178
rect 162228 191120 162674 191176
rect 162730 191120 162735 191176
rect 162228 191118 162735 191120
rect 162228 191116 162234 191118
rect 162669 191115 162735 191118
rect 165838 191116 165844 191180
rect 165908 191178 165914 191180
rect 166901 191178 166967 191181
rect 165908 191176 166967 191178
rect 165908 191120 166906 191176
rect 166962 191120 166967 191176
rect 165908 191118 166967 191120
rect 165908 191116 165914 191118
rect 166901 191115 166967 191118
rect 169293 191180 169359 191181
rect 169293 191176 169340 191180
rect 169404 191178 169410 191180
rect 169293 191120 169298 191176
rect 169293 191116 169340 191120
rect 169404 191118 169450 191178
rect 169404 191116 169410 191118
rect 171542 191116 171548 191180
rect 171612 191178 171618 191180
rect 172053 191178 172119 191181
rect 171612 191176 172119 191178
rect 171612 191120 172058 191176
rect 172114 191120 172119 191176
rect 171612 191118 172119 191120
rect 171612 191116 171618 191118
rect 169293 191115 169359 191116
rect 172053 191115 172119 191118
rect 172973 191180 173039 191181
rect 172973 191176 173020 191180
rect 173084 191178 173090 191180
rect 172973 191120 172978 191176
rect 172973 191116 173020 191120
rect 173084 191118 173130 191178
rect 173084 191116 173090 191118
rect 175774 191116 175780 191180
rect 175844 191178 175850 191180
rect 176469 191178 176535 191181
rect 175844 191176 176535 191178
rect 175844 191120 176474 191176
rect 176530 191120 176535 191176
rect 175844 191118 176535 191120
rect 175844 191116 175850 191118
rect 172973 191115 173039 191116
rect 176469 191115 176535 191118
rect 142153 191042 142219 191045
rect 142470 191042 142476 191044
rect 142153 191040 142476 191042
rect 142153 190984 142158 191040
rect 142214 190984 142476 191040
rect 142153 190982 142476 190984
rect 142153 190979 142219 190982
rect 142470 190980 142476 190982
rect 142540 190980 142546 191044
rect 150014 190980 150020 191044
rect 150084 191042 150090 191044
rect 159081 191042 159147 191045
rect 150084 191040 159147 191042
rect 150084 190984 159086 191040
rect 159142 190984 159147 191040
rect 150084 190982 159147 190984
rect 150084 190980 150090 190982
rect 159081 190979 159147 190982
rect 160870 190980 160876 191044
rect 160940 191042 160946 191044
rect 161381 191042 161447 191045
rect 160940 191040 161447 191042
rect 160940 190984 161386 191040
rect 161442 190984 161447 191040
rect 160940 190982 161447 190984
rect 160940 190980 160946 190982
rect 161381 190979 161447 190982
rect 172830 190980 172836 191044
rect 172900 191042 172906 191044
rect 173709 191042 173775 191045
rect 172900 191040 173775 191042
rect 172900 190984 173714 191040
rect 173770 190984 173775 191040
rect 172900 190982 173775 190984
rect 172900 190980 172906 190982
rect 173709 190979 173775 190982
rect 122557 190498 122623 190501
rect 122782 190498 122788 190500
rect 122557 190496 122788 190498
rect 122557 190440 122562 190496
rect 122618 190440 122788 190496
rect 122557 190438 122788 190440
rect 122557 190435 122623 190438
rect 122782 190436 122788 190438
rect 122852 190436 122858 190500
rect 122557 190362 122623 190365
rect 122782 190362 122788 190364
rect 122557 190360 122788 190362
rect 122557 190304 122562 190360
rect 122618 190304 122788 190360
rect 122557 190302 122788 190304
rect 122557 190299 122623 190302
rect 122782 190300 122788 190302
rect 122852 190300 122858 190364
rect 140814 190300 140820 190364
rect 140884 190362 140890 190364
rect 141693 190362 141759 190365
rect 140884 190360 141759 190362
rect 140884 190304 141698 190360
rect 141754 190304 141759 190360
rect 140884 190302 141759 190304
rect 140884 190300 140890 190302
rect 141693 190299 141759 190302
rect 165981 190090 166047 190093
rect 166206 190090 166212 190092
rect 165981 190088 166212 190090
rect 165981 190032 165986 190088
rect 166042 190032 166212 190088
rect 165981 190030 166212 190032
rect 165981 190027 166047 190030
rect 166206 190028 166212 190030
rect 166276 190028 166282 190092
rect 154941 189954 155007 189957
rect 155718 189954 155724 189956
rect 154941 189952 155724 189954
rect 154941 189896 154946 189952
rect 155002 189896 155724 189952
rect 154941 189894 155724 189896
rect 154941 189891 155007 189894
rect 155718 189892 155724 189894
rect 155788 189892 155794 189956
rect 157006 189212 157012 189276
rect 157076 189274 157082 189276
rect 158897 189274 158963 189277
rect 157076 189272 158963 189274
rect 157076 189216 158902 189272
rect 158958 189216 158963 189272
rect 157076 189214 158963 189216
rect 157076 189212 157082 189214
rect 158897 189211 158963 189214
rect 170397 189274 170463 189277
rect 170806 189274 170812 189276
rect 170397 189272 170812 189274
rect 170397 189216 170402 189272
rect 170458 189216 170812 189272
rect 170397 189214 170812 189216
rect 170397 189211 170463 189214
rect 170806 189212 170812 189214
rect 170876 189212 170882 189276
rect 133965 189138 134031 189141
rect 134374 189138 134380 189140
rect 133965 189136 134380 189138
rect 133965 189080 133970 189136
rect 134026 189080 134380 189136
rect 133965 189078 134380 189080
rect 133965 189075 134031 189078
rect 134374 189076 134380 189078
rect 134444 189076 134450 189140
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect 152549 188868 152615 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 138422 188804 138428 188868
rect 138492 188866 138498 188868
rect 143574 188866 143580 188868
rect 138492 188806 143580 188866
rect 138492 188804 138498 188806
rect 143574 188804 143580 188806
rect 143644 188804 143650 188868
rect 152549 188864 152596 188868
rect 152660 188866 152666 188868
rect 152549 188808 152554 188864
rect 152549 188804 152596 188808
rect 152660 188806 152706 188866
rect 152660 188804 152666 188806
rect 152549 188803 152615 188804
rect 138790 188532 138796 188596
rect 138860 188594 138866 188596
rect 138933 188594 138999 188597
rect 138860 188592 138999 188594
rect 138860 188536 138938 188592
rect 138994 188536 138999 188592
rect 138860 188534 138999 188536
rect 138860 188532 138866 188534
rect 138933 188531 138999 188534
rect 139761 188594 139827 188597
rect 140446 188594 140452 188596
rect 139761 188592 140452 188594
rect 139761 188536 139766 188592
rect 139822 188536 140452 188592
rect 139761 188534 140452 188536
rect 139761 188531 139827 188534
rect 140446 188532 140452 188534
rect 140516 188532 140522 188596
rect 164969 188594 165035 188597
rect 165102 188594 165108 188596
rect 164969 188592 165108 188594
rect 164969 188536 164974 188592
rect 165030 188536 165108 188592
rect 164969 188534 165108 188536
rect 164969 188531 165035 188534
rect 165102 188532 165108 188534
rect 165172 188532 165178 188596
rect 131614 188396 131620 188460
rect 131684 188458 131690 188460
rect 132309 188458 132375 188461
rect 131684 188456 132375 188458
rect 131684 188400 132314 188456
rect 132370 188400 132375 188456
rect 131684 188398 132375 188400
rect 131684 188396 131690 188398
rect 132309 188395 132375 188398
rect 135621 188458 135687 188461
rect 136030 188458 136036 188460
rect 135621 188456 136036 188458
rect 135621 188400 135626 188456
rect 135682 188400 136036 188456
rect 135621 188398 136036 188400
rect 135621 188395 135687 188398
rect 136030 188396 136036 188398
rect 136100 188396 136106 188460
rect 136582 188396 136588 188460
rect 136652 188458 136658 188460
rect 137001 188458 137067 188461
rect 136652 188456 137067 188458
rect 136652 188400 137006 188456
rect 137062 188400 137067 188456
rect 136652 188398 137067 188400
rect 136652 188396 136658 188398
rect 137001 188395 137067 188398
rect 137502 188396 137508 188460
rect 137572 188458 137578 188460
rect 137645 188458 137711 188461
rect 137572 188456 137711 188458
rect 137572 188400 137650 188456
rect 137706 188400 137711 188456
rect 137572 188398 137711 188400
rect 137572 188396 137578 188398
rect 137645 188395 137711 188398
rect 138422 188396 138428 188460
rect 138492 188458 138498 188460
rect 138841 188458 138907 188461
rect 138492 188456 138907 188458
rect 138492 188400 138846 188456
rect 138902 188400 138907 188456
rect 138492 188398 138907 188400
rect 138492 188396 138498 188398
rect 138841 188395 138907 188398
rect 140262 188396 140268 188460
rect 140332 188458 140338 188460
rect 140405 188458 140471 188461
rect 140332 188456 140471 188458
rect 140332 188400 140410 188456
rect 140466 188400 140471 188456
rect 140332 188398 140471 188400
rect 140332 188396 140338 188398
rect 140405 188395 140471 188398
rect 149830 188396 149836 188460
rect 149900 188458 149906 188460
rect 149973 188458 150039 188461
rect 149900 188456 150039 188458
rect 149900 188400 149978 188456
rect 150034 188400 150039 188456
rect 149900 188398 150039 188400
rect 149900 188396 149906 188398
rect 149973 188395 150039 188398
rect 176193 188458 176259 188461
rect 176510 188458 176516 188460
rect 176193 188456 176516 188458
rect 176193 188400 176198 188456
rect 176254 188400 176516 188456
rect 176193 188398 176516 188400
rect 176193 188395 176259 188398
rect 176510 188396 176516 188398
rect 176580 188396 176586 188460
rect 176878 188396 176884 188460
rect 176948 188458 176954 188460
rect 177481 188458 177547 188461
rect 176948 188456 177547 188458
rect 176948 188400 177486 188456
rect 177542 188400 177547 188456
rect 176948 188398 177547 188400
rect 176948 188396 176954 188398
rect 177481 188395 177547 188398
rect 130510 188260 130516 188324
rect 130580 188322 130586 188324
rect 144453 188322 144519 188325
rect 130580 188320 144519 188322
rect 130580 188264 144458 188320
rect 144514 188264 144519 188320
rect 130580 188262 144519 188264
rect 130580 188260 130586 188262
rect 144453 188259 144519 188262
rect 176694 188260 176700 188324
rect 176764 188322 176770 188324
rect 177297 188322 177363 188325
rect 176764 188320 177363 188322
rect 176764 188264 177302 188320
rect 177358 188264 177363 188320
rect 176764 188262 177363 188264
rect 176764 188260 176770 188262
rect 177297 188259 177363 188262
rect 130694 188124 130700 188188
rect 130764 188186 130770 188188
rect 144126 188186 144132 188188
rect 130764 188126 144132 188186
rect 130764 188124 130770 188126
rect 144126 188124 144132 188126
rect 144196 188124 144202 188188
rect 137277 188050 137343 188053
rect 138606 188050 138612 188052
rect 137277 188048 138612 188050
rect 137277 187992 137282 188048
rect 137338 187992 138612 188048
rect 137277 187990 138612 187992
rect 137277 187987 137343 187990
rect 138606 187988 138612 187990
rect 138676 187988 138682 188052
rect 176653 188050 176719 188053
rect 198774 188050 198780 188052
rect 176653 188048 198780 188050
rect 176653 187992 176658 188048
rect 176714 187992 198780 188048
rect 176653 187990 198780 187992
rect 176653 187987 176719 187990
rect 198774 187988 198780 187990
rect 198844 187988 198850 188052
rect 175457 187778 175523 187781
rect 176142 187778 176148 187780
rect 175457 187776 176148 187778
rect 175457 187720 175462 187776
rect 175518 187720 176148 187776
rect 175457 187718 176148 187720
rect 175457 187715 175523 187718
rect 176142 187716 176148 187718
rect 176212 187716 176218 187780
rect 137185 187642 137251 187645
rect 142286 187642 142292 187644
rect 137185 187640 142292 187642
rect 137185 187584 137190 187640
rect 137246 187584 142292 187640
rect 137185 187582 142292 187584
rect 137185 187579 137251 187582
rect 142286 187580 142292 187582
rect 142356 187580 142362 187644
rect 161974 187444 161980 187508
rect 162044 187506 162050 187508
rect 162485 187506 162551 187509
rect 162044 187504 162551 187506
rect 162044 187448 162490 187504
rect 162546 187448 162551 187504
rect 162044 187446 162551 187448
rect 162044 187444 162050 187446
rect 162485 187443 162551 187446
rect 152733 187372 152799 187373
rect 152733 187368 152780 187372
rect 152844 187370 152850 187372
rect 152733 187312 152738 187368
rect 152733 187308 152780 187312
rect 152844 187310 152890 187370
rect 152844 187308 152850 187310
rect 163262 187308 163268 187372
rect 163332 187370 163338 187372
rect 163865 187370 163931 187373
rect 163332 187368 163931 187370
rect 163332 187312 163870 187368
rect 163926 187312 163931 187368
rect 163332 187310 163931 187312
rect 163332 187308 163338 187310
rect 152733 187307 152799 187308
rect 163865 187307 163931 187310
rect 135437 187098 135503 187101
rect 136398 187098 136404 187100
rect 135437 187096 136404 187098
rect 135437 187040 135442 187096
rect 135498 187040 136404 187096
rect 135437 187038 136404 187040
rect 135437 187035 135503 187038
rect 136398 187036 136404 187038
rect 136468 187036 136474 187100
rect 161933 187098 161999 187101
rect 178534 187098 178540 187100
rect 161933 187096 178540 187098
rect 161933 187040 161938 187096
rect 161994 187040 178540 187096
rect 161933 187038 178540 187040
rect 161933 187035 161999 187038
rect 178534 187036 178540 187038
rect 178604 187036 178610 187100
rect 137461 186282 137527 186285
rect 137686 186282 137692 186284
rect 137461 186280 137692 186282
rect 137461 186224 137466 186280
rect 137522 186224 137692 186280
rect 137461 186222 137692 186224
rect 137461 186219 137527 186222
rect 137686 186220 137692 186222
rect 137756 186220 137762 186284
rect 165286 185812 165292 185876
rect 165356 185874 165362 185876
rect 165429 185874 165495 185877
rect 165356 185872 165495 185874
rect 165356 185816 165434 185872
rect 165490 185816 165495 185872
rect 165356 185814 165495 185816
rect 165356 185812 165362 185814
rect 165429 185811 165495 185814
rect 168741 185874 168807 185877
rect 168966 185874 168972 185876
rect 168741 185872 168972 185874
rect 168741 185816 168746 185872
rect 168802 185816 168972 185872
rect 168741 185814 168972 185816
rect 168741 185811 168807 185814
rect 168966 185812 168972 185814
rect 169036 185812 169042 185876
rect 147438 184044 147444 184108
rect 147508 184106 147514 184108
rect 159357 184106 159423 184109
rect 147508 184104 159423 184106
rect 147508 184048 159362 184104
rect 159418 184048 159423 184104
rect 147508 184046 159423 184048
rect 147508 184044 147514 184046
rect 159357 184043 159423 184046
rect 125174 183772 125180 183836
rect 125244 183834 125250 183836
rect 144637 183834 144703 183837
rect 125244 183832 144703 183834
rect 125244 183776 144642 183832
rect 144698 183776 144703 183832
rect 125244 183774 144703 183776
rect 125244 183772 125250 183774
rect 144637 183771 144703 183774
rect 164918 182548 164924 182612
rect 164988 182610 164994 182612
rect 165245 182610 165311 182613
rect 164988 182608 165311 182610
rect 164988 182552 165250 182608
rect 165306 182552 165311 182608
rect 164988 182550 165311 182552
rect 164988 182548 164994 182550
rect 165245 182547 165311 182550
rect 142102 180916 142108 180980
rect 142172 180916 142178 180980
rect 142110 180845 142170 180916
rect 122557 180842 122623 180845
rect 122966 180842 122972 180844
rect 122557 180840 122972 180842
rect 122557 180784 122562 180840
rect 122618 180784 122972 180840
rect 122557 180782 122972 180784
rect 122557 180779 122623 180782
rect 122966 180780 122972 180782
rect 123036 180780 123042 180844
rect 142061 180842 142170 180845
rect 142016 180840 142170 180842
rect 142016 180784 142066 180840
rect 142122 180784 142170 180840
rect 142016 180782 142170 180784
rect 142061 180779 142127 180782
rect 142061 180708 142127 180709
rect 142061 180706 142108 180708
rect 142016 180704 142108 180706
rect 142172 180706 142178 180708
rect 142016 180648 142066 180704
rect 142016 180646 142108 180648
rect 142061 180644 142108 180646
rect 142172 180646 142254 180706
rect 142172 180644 142178 180646
rect 142061 180643 142127 180644
rect 195513 179346 195579 179349
rect 196014 179346 196020 179348
rect 195513 179344 196020 179346
rect 195513 179288 195518 179344
rect 195574 179288 196020 179344
rect 195513 179286 196020 179288
rect 195513 179283 195579 179286
rect 196014 179284 196020 179286
rect 196084 179284 196090 179348
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 142102 171260 142108 171324
rect 142172 171260 142178 171324
rect 142110 171189 142170 171260
rect 142061 171186 142170 171189
rect 142016 171184 142170 171186
rect 142016 171128 142066 171184
rect 142122 171128 142170 171184
rect 142016 171126 142170 171128
rect 142061 171123 142127 171126
rect 142061 171050 142127 171053
rect 142016 171048 142170 171050
rect 142016 170992 142066 171048
rect 142122 170992 142170 171048
rect 142016 170990 142170 170992
rect 142061 170987 142170 170990
rect 142110 170916 142170 170987
rect 142102 170852 142108 170916
rect 142172 170852 142178 170916
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 142061 161532 142127 161533
rect 142061 161530 142108 161532
rect 142016 161528 142108 161530
rect 142172 161530 142178 161532
rect 142016 161472 142066 161528
rect 142016 161470 142108 161472
rect 142061 161468 142108 161470
rect 142172 161470 142254 161530
rect 142172 161468 142178 161470
rect 142061 161467 142127 161468
rect 142061 161396 142127 161397
rect 142061 161394 142108 161396
rect 142016 161392 142108 161394
rect 142172 161394 142178 161396
rect 142016 161336 142066 161392
rect 142016 161334 142108 161336
rect 142061 161332 142108 161334
rect 142172 161334 142254 161394
rect 142172 161332 142178 161334
rect 142061 161331 142127 161332
rect 162342 154396 162348 154460
rect 162412 154458 162418 154460
rect 168465 154458 168531 154461
rect 162412 154456 168531 154458
rect 162412 154400 168470 154456
rect 168526 154400 168531 154456
rect 162412 154398 168531 154400
rect 162412 154396 162418 154398
rect 168465 154395 168531 154398
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 580349 152627 580415 152630
rect 165889 152554 165955 152557
rect 186078 152554 186084 152556
rect 165889 152552 186084 152554
rect 165889 152496 165894 152552
rect 165950 152496 186084 152552
rect 165889 152494 186084 152496
rect 165889 152491 165955 152494
rect 186078 152492 186084 152494
rect 186148 152492 186154 152556
rect 583520 152540 584960 152630
rect 168281 152418 168347 152421
rect 202137 152418 202203 152421
rect 168281 152416 202203 152418
rect 168281 152360 168286 152416
rect 168342 152360 202142 152416
rect 202198 152360 202203 152416
rect 168281 152358 202203 152360
rect 168281 152355 168347 152358
rect 202137 152355 202203 152358
rect 142102 151948 142108 152012
rect 142172 151948 142178 152012
rect 142110 151877 142170 151948
rect 142061 151874 142170 151877
rect 142016 151872 142170 151874
rect 142016 151816 142066 151872
rect 142122 151816 142170 151872
rect 142016 151814 142170 151816
rect 142061 151811 142127 151814
rect 142061 151738 142127 151741
rect 142016 151736 142170 151738
rect 142016 151680 142066 151736
rect 142122 151680 142170 151736
rect 142016 151678 142170 151680
rect 142061 151675 142170 151678
rect 142110 151604 142170 151675
rect 142102 151540 142108 151604
rect 142172 151540 142178 151604
rect 117681 151194 117747 151197
rect 142654 151194 142660 151196
rect 117681 151192 142660 151194
rect 117681 151136 117686 151192
rect 117742 151136 142660 151192
rect 117681 151134 142660 151136
rect 117681 151131 117747 151134
rect 142654 151132 142660 151134
rect 142724 151132 142730 151196
rect 116301 151058 116367 151061
rect 142470 151058 142476 151060
rect 116301 151056 142476 151058
rect 116301 151000 116306 151056
rect 116362 151000 142476 151056
rect 116301 150998 142476 151000
rect 116301 150995 116367 150998
rect 142470 150996 142476 150998
rect 142540 150996 142546 151060
rect 157609 150378 157675 150381
rect 182766 150378 182772 150380
rect 157609 150376 182772 150378
rect 157609 150320 157614 150376
rect 157670 150320 182772 150376
rect 157609 150318 182772 150320
rect 157609 150315 157675 150318
rect 182766 150316 182772 150318
rect 182836 150316 182842 150380
rect 201401 150378 201467 150381
rect 201718 150378 201724 150380
rect 201401 150376 201724 150378
rect 201401 150320 201406 150376
rect 201462 150320 201724 150376
rect 201401 150318 201724 150320
rect 201401 150315 201467 150318
rect 201718 150316 201724 150318
rect 201788 150316 201794 150380
rect 202781 150378 202847 150381
rect 203006 150378 203012 150380
rect 202781 150376 203012 150378
rect 202781 150320 202786 150376
rect 202842 150320 203012 150376
rect 202781 150318 203012 150320
rect 202781 150315 202847 150318
rect 203006 150316 203012 150318
rect 203076 150316 203082 150380
rect 157425 150242 157491 150245
rect 183870 150242 183876 150244
rect 157425 150240 183876 150242
rect 157425 150184 157430 150240
rect 157486 150184 183876 150240
rect 157425 150182 183876 150184
rect 157425 150179 157491 150182
rect 183870 150180 183876 150182
rect 183940 150180 183946 150244
rect 174261 150106 174327 150109
rect 201534 150106 201540 150108
rect 174261 150104 201540 150106
rect 174261 150048 174266 150104
rect 174322 150048 201540 150104
rect 174261 150046 201540 150048
rect 174261 150043 174327 150046
rect 201534 150044 201540 150046
rect 201604 150044 201610 150108
rect 157241 149970 157307 149973
rect 185158 149970 185164 149972
rect 157241 149968 185164 149970
rect -960 149834 480 149924
rect 157241 149912 157246 149968
rect 157302 149912 185164 149968
rect 157241 149910 185164 149912
rect 157241 149907 157307 149910
rect 185158 149908 185164 149910
rect 185228 149908 185234 149972
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 154941 149834 155007 149837
rect 184054 149834 184060 149836
rect 154941 149832 184060 149834
rect 154941 149776 154946 149832
rect 155002 149776 184060 149832
rect 154941 149774 184060 149776
rect 154941 149771 155007 149774
rect 184054 149772 184060 149774
rect 184124 149772 184130 149836
rect 150341 149698 150407 149701
rect 185342 149698 185348 149700
rect 150341 149696 185348 149698
rect 150341 149640 150346 149696
rect 150402 149640 185348 149696
rect 150341 149638 185348 149640
rect 150341 149635 150407 149638
rect 185342 149636 185348 149638
rect 185412 149636 185418 149700
rect 157793 149562 157859 149565
rect 181110 149562 181116 149564
rect 157793 149560 181116 149562
rect 157793 149504 157798 149560
rect 157854 149504 181116 149560
rect 157793 149502 181116 149504
rect 157793 149499 157859 149502
rect 181110 149500 181116 149502
rect 181180 149500 181186 149564
rect 122833 149020 122899 149021
rect 122782 148956 122788 149020
rect 122852 149018 122899 149020
rect 122852 149016 122944 149018
rect 122894 148960 122944 149016
rect 122852 148958 122944 148960
rect 122852 148956 122899 148958
rect 122833 148955 122899 148956
rect 125225 148610 125291 148613
rect 145741 148610 145807 148613
rect 125225 148608 145807 148610
rect 125225 148552 125230 148608
rect 125286 148552 145746 148608
rect 145802 148552 145807 148608
rect 125225 148550 145807 148552
rect 125225 148547 125291 148550
rect 145741 148547 145807 148550
rect 122966 148412 122972 148476
rect 123036 148474 123042 148476
rect 153377 148474 153443 148477
rect 123036 148472 153443 148474
rect 123036 148416 153382 148472
rect 153438 148416 153443 148472
rect 123036 148414 153443 148416
rect 123036 148412 123042 148414
rect 153377 148411 153443 148414
rect 100477 148338 100543 148341
rect 133045 148338 133111 148341
rect 100477 148336 133111 148338
rect 100477 148280 100482 148336
rect 100538 148280 133050 148336
rect 133106 148280 133111 148336
rect 100477 148278 133111 148280
rect 100477 148275 100543 148278
rect 133045 148275 133111 148278
rect 197854 147732 197860 147796
rect 197924 147794 197930 147796
rect 198181 147794 198247 147797
rect 197924 147792 198247 147794
rect 197924 147736 198186 147792
rect 198242 147736 198247 147792
rect 197924 147734 198247 147736
rect 197924 147732 197930 147734
rect 198181 147731 198247 147734
rect 156045 147386 156111 147389
rect 182950 147386 182956 147388
rect 156045 147384 182956 147386
rect 156045 147328 156050 147384
rect 156106 147328 182956 147384
rect 156045 147326 182956 147328
rect 156045 147323 156111 147326
rect 182950 147324 182956 147326
rect 183020 147324 183026 147388
rect 154757 147250 154823 147253
rect 181294 147250 181300 147252
rect 154757 147248 181300 147250
rect 154757 147192 154762 147248
rect 154818 147192 181300 147248
rect 154757 147190 181300 147192
rect 154757 147187 154823 147190
rect 181294 147188 181300 147190
rect 181364 147188 181370 147252
rect 172605 147114 172671 147117
rect 202822 147114 202828 147116
rect 172605 147112 202828 147114
rect 172605 147056 172610 147112
rect 172666 147056 202828 147112
rect 172605 147054 202828 147056
rect 172605 147051 172671 147054
rect 202822 147052 202828 147054
rect 202892 147052 202898 147116
rect 113449 146978 113515 146981
rect 143574 146978 143580 146980
rect 113449 146976 143580 146978
rect 113449 146920 113454 146976
rect 113510 146920 143580 146976
rect 113449 146918 143580 146920
rect 113449 146915 113515 146918
rect 143574 146916 143580 146918
rect 143644 146916 143650 146980
rect 147581 146978 147647 146981
rect 179822 146978 179828 146980
rect 147581 146976 179828 146978
rect 147581 146920 147586 146976
rect 147642 146920 179828 146976
rect 147581 146918 179828 146920
rect 147581 146915 147647 146918
rect 179822 146916 179828 146918
rect 179892 146916 179898 146980
rect 126973 146434 127039 146437
rect 580257 146434 580323 146437
rect 126973 146432 580323 146434
rect 126973 146376 126978 146432
rect 127034 146376 580262 146432
rect 580318 146376 580323 146432
rect 126973 146374 580323 146376
rect 126973 146371 127039 146374
rect 580257 146371 580323 146374
rect 116894 146236 116900 146300
rect 116964 146298 116970 146300
rect 130285 146298 130351 146301
rect 116964 146296 130351 146298
rect 116964 146240 130290 146296
rect 130346 146240 130351 146296
rect 116964 146238 130351 146240
rect 116964 146236 116970 146238
rect 130285 146235 130351 146238
rect 174077 146298 174143 146301
rect 188521 146298 188587 146301
rect 174077 146296 188587 146298
rect 174077 146240 174082 146296
rect 174138 146240 188526 146296
rect 188582 146240 188587 146296
rect 174077 146238 188587 146240
rect 174077 146235 174143 146238
rect 188521 146235 188587 146238
rect 193857 146298 193923 146301
rect 193990 146298 193996 146300
rect 193857 146296 193996 146298
rect 193857 146240 193862 146296
rect 193918 146240 193996 146296
rect 193857 146238 193996 146240
rect 193857 146235 193923 146238
rect 193990 146236 193996 146238
rect 194060 146236 194066 146300
rect 198733 146298 198799 146301
rect 199326 146298 199332 146300
rect 198733 146296 199332 146298
rect 198733 146240 198738 146296
rect 198794 146240 199332 146296
rect 198733 146238 199332 146240
rect 198733 146235 198799 146238
rect 199326 146236 199332 146238
rect 199396 146236 199402 146300
rect 112846 146100 112852 146164
rect 112916 146162 112922 146164
rect 129825 146162 129891 146165
rect 112916 146160 129891 146162
rect 112916 146104 129830 146160
rect 129886 146104 129891 146160
rect 112916 146102 129891 146104
rect 112916 146100 112922 146102
rect 129825 146099 129891 146102
rect 173893 146162 173959 146165
rect 193121 146162 193187 146165
rect 173893 146160 193187 146162
rect 173893 146104 173898 146160
rect 173954 146104 193126 146160
rect 193182 146104 193187 146160
rect 173893 146102 193187 146104
rect 173893 146099 173959 146102
rect 193121 146099 193187 146102
rect 193806 146100 193812 146164
rect 193876 146162 193882 146164
rect 194041 146162 194107 146165
rect 193876 146160 194107 146162
rect 193876 146104 194046 146160
rect 194102 146104 194107 146160
rect 193876 146102 194107 146104
rect 193876 146100 193882 146102
rect 194041 146099 194107 146102
rect 111558 145964 111564 146028
rect 111628 146026 111634 146028
rect 129917 146026 129983 146029
rect 111628 146024 129983 146026
rect 111628 145968 129922 146024
rect 129978 145968 129983 146024
rect 111628 145966 129983 145968
rect 111628 145964 111634 145966
rect 129917 145963 129983 145966
rect 164417 146026 164483 146029
rect 195053 146026 195119 146029
rect 164417 146024 195119 146026
rect 164417 145968 164422 146024
rect 164478 145968 195058 146024
rect 195114 145968 195119 146024
rect 164417 145966 195119 145968
rect 164417 145963 164483 145966
rect 195053 145963 195119 145966
rect 111374 145828 111380 145892
rect 111444 145890 111450 145892
rect 131113 145890 131179 145893
rect 111444 145888 131179 145890
rect 111444 145832 131118 145888
rect 131174 145832 131179 145888
rect 111444 145830 131179 145832
rect 111444 145828 111450 145830
rect 131113 145827 131179 145830
rect 162301 145890 162367 145893
rect 194726 145890 194732 145892
rect 162301 145888 194732 145890
rect 162301 145832 162306 145888
rect 162362 145832 194732 145888
rect 162301 145830 194732 145832
rect 162301 145827 162367 145830
rect 194726 145828 194732 145830
rect 194796 145828 194802 145892
rect 116710 145692 116716 145756
rect 116780 145754 116786 145756
rect 116853 145754 116919 145757
rect 116780 145752 116919 145754
rect 116780 145696 116858 145752
rect 116914 145696 116919 145752
rect 116780 145694 116919 145696
rect 116780 145692 116786 145694
rect 116853 145691 116919 145694
rect 118366 145692 118372 145756
rect 118436 145754 118442 145756
rect 146293 145754 146359 145757
rect 118436 145752 146359 145754
rect 118436 145696 146298 145752
rect 146354 145696 146359 145752
rect 118436 145694 146359 145696
rect 118436 145692 118442 145694
rect 146293 145691 146359 145694
rect 160645 145754 160711 145757
rect 193254 145754 193260 145756
rect 160645 145752 193260 145754
rect 160645 145696 160650 145752
rect 160706 145696 193260 145752
rect 160645 145694 193260 145696
rect 160645 145691 160711 145694
rect 193254 145692 193260 145694
rect 193324 145692 193330 145756
rect 118182 145556 118188 145620
rect 118252 145618 118258 145620
rect 147673 145618 147739 145621
rect 118252 145616 147739 145618
rect 118252 145560 147678 145616
rect 147734 145560 147739 145616
rect 118252 145558 147739 145560
rect 118252 145556 118258 145558
rect 147673 145555 147739 145558
rect 153285 145618 153351 145621
rect 187141 145618 187207 145621
rect 153285 145616 187207 145618
rect 153285 145560 153290 145616
rect 153346 145560 187146 145616
rect 187202 145560 187207 145616
rect 153285 145558 187207 145560
rect 153285 145555 153351 145558
rect 187141 145555 187207 145558
rect 193121 145618 193187 145621
rect 199561 145618 199627 145621
rect 193121 145616 199627 145618
rect 193121 145560 193126 145616
rect 193182 145560 199566 145616
rect 199622 145560 199627 145616
rect 193121 145558 199627 145560
rect 193121 145555 193187 145558
rect 199561 145555 199627 145558
rect 119654 144740 119660 144804
rect 119724 144802 119730 144804
rect 119981 144802 120047 144805
rect 119724 144800 120047 144802
rect 119724 144744 119986 144800
rect 120042 144744 120047 144800
rect 119724 144742 120047 144744
rect 119724 144740 119730 144742
rect 119981 144739 120047 144742
rect 168005 144802 168071 144805
rect 196198 144802 196204 144804
rect 168005 144800 196204 144802
rect 168005 144744 168010 144800
rect 168066 144744 196204 144800
rect 168005 144742 196204 144744
rect 168005 144739 168071 144742
rect 196198 144740 196204 144742
rect 196268 144740 196274 144804
rect 113950 144604 113956 144668
rect 114020 144666 114026 144668
rect 140865 144666 140931 144669
rect 114020 144664 140931 144666
rect 114020 144608 140870 144664
rect 140926 144608 140931 144664
rect 114020 144606 140931 144608
rect 114020 144604 114026 144606
rect 140865 144603 140931 144606
rect 166349 144666 166415 144669
rect 197486 144666 197492 144668
rect 166349 144664 197492 144666
rect 166349 144608 166354 144664
rect 166410 144608 197492 144664
rect 166349 144606 197492 144608
rect 166349 144603 166415 144606
rect 197486 144604 197492 144606
rect 197556 144604 197562 144668
rect 114134 144468 114140 144532
rect 114204 144530 114210 144532
rect 142521 144530 142587 144533
rect 114204 144528 142587 144530
rect 114204 144472 142526 144528
rect 142582 144472 142587 144528
rect 114204 144470 142587 144472
rect 114204 144468 114210 144470
rect 142521 144467 142587 144470
rect 162209 144530 162275 144533
rect 193438 144530 193444 144532
rect 162209 144528 193444 144530
rect 162209 144472 162214 144528
rect 162270 144472 193444 144528
rect 162209 144470 193444 144472
rect 162209 144467 162275 144470
rect 193438 144468 193444 144470
rect 193508 144468 193514 144532
rect 115422 144332 115428 144396
rect 115492 144394 115498 144396
rect 144177 144394 144243 144397
rect 115492 144392 144243 144394
rect 115492 144336 144182 144392
rect 144238 144336 144243 144392
rect 115492 144334 144243 144336
rect 115492 144332 115498 144334
rect 144177 144331 144243 144334
rect 154481 144394 154547 144397
rect 187918 144394 187924 144396
rect 154481 144392 187924 144394
rect 154481 144336 154486 144392
rect 154542 144336 187924 144392
rect 154481 144334 187924 144336
rect 154481 144331 154547 144334
rect 187918 144332 187924 144334
rect 187988 144332 187994 144396
rect 115790 144196 115796 144260
rect 115860 144258 115866 144260
rect 145833 144258 145899 144261
rect 115860 144256 145899 144258
rect 115860 144200 145838 144256
rect 145894 144200 145899 144256
rect 115860 144198 145899 144200
rect 115860 144196 115866 144198
rect 145833 144195 145899 144198
rect 159449 144258 159515 144261
rect 193622 144258 193628 144260
rect 159449 144256 193628 144258
rect 159449 144200 159454 144256
rect 159510 144200 193628 144256
rect 159449 144198 193628 144200
rect 159449 144195 159515 144198
rect 193622 144196 193628 144198
rect 193692 144196 193698 144260
rect 119838 144060 119844 144124
rect 119908 144122 119914 144124
rect 151077 144122 151143 144125
rect 119908 144120 151143 144122
rect 119908 144064 151082 144120
rect 151138 144064 151143 144120
rect 119908 144062 151143 144064
rect 119908 144060 119914 144062
rect 151077 144059 151143 144062
rect 158069 144122 158135 144125
rect 192334 144122 192340 144124
rect 158069 144120 192340 144122
rect 158069 144064 158074 144120
rect 158130 144064 192340 144120
rect 158069 144062 192340 144064
rect 158069 144059 158135 144062
rect 192334 144060 192340 144062
rect 192404 144060 192410 144124
rect 113766 143924 113772 143988
rect 113836 143986 113842 143988
rect 138657 143986 138723 143989
rect 113836 143984 138723 143986
rect 113836 143928 138662 143984
rect 138718 143928 138723 143984
rect 113836 143926 138723 143928
rect 113836 143924 113842 143926
rect 138657 143923 138723 143926
rect 165521 143986 165587 143989
rect 192150 143986 192156 143988
rect 165521 143984 192156 143986
rect 165521 143928 165526 143984
rect 165582 143928 192156 143984
rect 165521 143926 192156 143928
rect 165521 143923 165587 143926
rect 192150 143924 192156 143926
rect 192220 143924 192226 143988
rect 113030 143788 113036 143852
rect 113100 143850 113106 143852
rect 139393 143850 139459 143853
rect 113100 143848 139459 143850
rect 113100 143792 139398 143848
rect 139454 143792 139459 143848
rect 113100 143790 139459 143792
rect 113100 143788 113106 143790
rect 139393 143787 139459 143790
rect 120717 143442 120783 143445
rect 126789 143442 126855 143445
rect 120717 143440 126855 143442
rect 120717 143384 120722 143440
rect 120778 143384 126794 143440
rect 126850 143384 126855 143440
rect 120717 143382 126855 143384
rect 120717 143379 120783 143382
rect 126789 143379 126855 143382
rect 165245 143442 165311 143445
rect 187969 143442 188035 143445
rect 165245 143440 188035 143442
rect 165245 143384 165250 143440
rect 165306 143384 187974 143440
rect 188030 143384 188035 143440
rect 165245 143382 188035 143384
rect 165245 143379 165311 143382
rect 187969 143379 188035 143382
rect 121729 143306 121795 143309
rect 143073 143306 143139 143309
rect 121729 143304 143139 143306
rect 121729 143248 121734 143304
rect 121790 143248 143078 143304
rect 143134 143248 143139 143304
rect 121729 143246 143139 143248
rect 121729 143243 121795 143246
rect 143073 143243 143139 143246
rect 163589 143306 163655 143309
rect 188102 143306 188108 143308
rect 163589 143304 188108 143306
rect 163589 143248 163594 143304
rect 163650 143248 188108 143304
rect 163589 143246 188108 143248
rect 163589 143243 163655 143246
rect 188102 143244 188108 143246
rect 188172 143244 188178 143308
rect 122414 143108 122420 143172
rect 122484 143170 122490 143172
rect 146385 143170 146451 143173
rect 122484 143168 146451 143170
rect 122484 143112 146390 143168
rect 146446 143112 146451 143168
rect 122484 143110 146451 143112
rect 122484 143108 122490 143110
rect 146385 143107 146451 143110
rect 161933 143170 161999 143173
rect 188286 143170 188292 143172
rect 161933 143168 188292 143170
rect 161933 143112 161938 143168
rect 161994 143112 188292 143168
rect 161933 143110 188292 143112
rect 161933 143107 161999 143110
rect 188286 143108 188292 143110
rect 188356 143108 188362 143172
rect 120942 142972 120948 143036
rect 121012 143034 121018 143036
rect 145005 143034 145071 143037
rect 121012 143032 145071 143034
rect 121012 142976 145010 143032
rect 145066 142976 145071 143032
rect 121012 142974 145071 142976
rect 121012 142972 121018 142974
rect 145005 142971 145071 142974
rect 160001 143034 160067 143037
rect 188061 143034 188127 143037
rect 160001 143032 188127 143034
rect 160001 142976 160006 143032
rect 160062 142976 188066 143032
rect 188122 142976 188127 143032
rect 160001 142974 188127 142976
rect 160001 142971 160067 142974
rect 188061 142971 188127 142974
rect 121126 142836 121132 142900
rect 121196 142898 121202 142900
rect 148041 142898 148107 142901
rect 121196 142896 148107 142898
rect 121196 142840 148046 142896
rect 148102 142840 148107 142896
rect 121196 142838 148107 142840
rect 121196 142836 121202 142838
rect 148041 142835 148107 142838
rect 155125 142898 155191 142901
rect 187734 142898 187740 142900
rect 155125 142896 187740 142898
rect 155125 142840 155130 142896
rect 155186 142840 187740 142896
rect 155125 142838 187740 142840
rect 155125 142835 155191 142838
rect 187734 142836 187740 142838
rect 187804 142836 187810 142900
rect 122230 142700 122236 142764
rect 122300 142762 122306 142764
rect 149697 142762 149763 142765
rect 122300 142760 149763 142762
rect 122300 142704 149702 142760
rect 149758 142704 149763 142760
rect 122300 142702 149763 142704
rect 122300 142700 122306 142702
rect 149697 142699 149763 142702
rect 156965 142762 157031 142765
rect 189022 142762 189028 142764
rect 156965 142760 189028 142762
rect 156965 142704 156970 142760
rect 157026 142704 189028 142760
rect 156965 142702 189028 142704
rect 156965 142699 157031 142702
rect 189022 142700 189028 142702
rect 189092 142700 189098 142764
rect 142061 142356 142127 142357
rect 142061 142354 142108 142356
rect 142016 142352 142108 142354
rect 142172 142354 142178 142356
rect 142016 142296 142066 142352
rect 142016 142294 142108 142296
rect 142061 142292 142108 142294
rect 142172 142294 142254 142354
rect 142172 142292 142178 142294
rect 142061 142291 142127 142292
rect 126789 142218 126855 142221
rect 191598 142218 191604 142220
rect 126789 142216 191604 142218
rect 126789 142160 126794 142216
rect 126850 142160 191604 142216
rect 126789 142158 191604 142160
rect 126789 142155 126855 142158
rect 191598 142156 191604 142158
rect 191668 142156 191674 142220
rect 157333 142082 157399 142085
rect 189574 142082 189580 142084
rect 157333 142080 189580 142082
rect 157333 142024 157338 142080
rect 157394 142024 189580 142080
rect 157333 142022 189580 142024
rect 157333 142019 157399 142022
rect 189574 142020 189580 142022
rect 189644 142020 189650 142084
rect 115606 141612 115612 141676
rect 115676 141674 115682 141676
rect 125593 141674 125659 141677
rect 143625 141674 143691 141677
rect 115676 141672 125659 141674
rect 115676 141616 125598 141672
rect 125654 141616 125659 141672
rect 115676 141614 125659 141616
rect 115676 141612 115682 141614
rect 125593 141611 125659 141614
rect 132450 141672 143691 141674
rect 132450 141616 143630 141672
rect 143686 141616 143691 141672
rect 132450 141614 143691 141616
rect 118550 141476 118556 141540
rect 118620 141538 118626 141540
rect 132450 141538 132510 141614
rect 143625 141611 143691 141614
rect 176653 141674 176719 141677
rect 177614 141674 177620 141676
rect 176653 141672 177620 141674
rect 176653 141616 176658 141672
rect 176714 141616 177620 141672
rect 176653 141614 177620 141616
rect 176653 141611 176719 141614
rect 177614 141612 177620 141614
rect 177684 141612 177690 141676
rect 118620 141478 132510 141538
rect 141417 141538 141483 141541
rect 141734 141538 141740 141540
rect 141417 141536 141740 141538
rect 141417 141480 141422 141536
rect 141478 141480 141740 141536
rect 141417 141478 141740 141480
rect 118620 141476 118626 141478
rect 141417 141475 141483 141478
rect 141734 141476 141740 141478
rect 141804 141476 141810 141540
rect 164141 141538 164207 141541
rect 191966 141538 191972 141540
rect 164141 141536 191972 141538
rect 164141 141480 164146 141536
rect 164202 141480 191972 141536
rect 164141 141478 191972 141480
rect 164141 141475 164207 141478
rect 191966 141476 191972 141478
rect 192036 141476 192042 141540
rect 117078 141340 117084 141404
rect 117148 141402 117154 141404
rect 150433 141402 150499 141405
rect 117148 141400 150499 141402
rect 117148 141344 150438 141400
rect 150494 141344 150499 141400
rect 117148 141342 150499 141344
rect 117148 141340 117154 141342
rect 150433 141339 150499 141342
rect 157149 141402 157215 141405
rect 189390 141402 189396 141404
rect 157149 141400 189396 141402
rect 157149 141344 157154 141400
rect 157210 141344 189396 141400
rect 157149 141342 189396 141344
rect 157149 141339 157215 141342
rect 189390 141340 189396 141342
rect 189460 141340 189466 141404
rect 141366 141204 141372 141268
rect 141436 141266 141442 141268
rect 141601 141266 141667 141269
rect 141436 141264 141667 141266
rect 141436 141208 141606 141264
rect 141662 141208 141667 141264
rect 141436 141206 141667 141208
rect 141436 141204 141442 141206
rect 141601 141203 141667 141206
rect 176745 141266 176811 141269
rect 177430 141266 177436 141268
rect 176745 141264 177436 141266
rect 176745 141208 176750 141264
rect 176806 141208 177436 141264
rect 176745 141206 177436 141208
rect 176745 141203 176811 141206
rect 177430 141204 177436 141206
rect 177500 141204 177506 141268
rect 127341 141130 127407 141133
rect 188286 141130 188292 141132
rect 127341 141128 188292 141130
rect 127341 141072 127346 141128
rect 127402 141072 188292 141128
rect 127341 141070 188292 141072
rect 127341 141067 127407 141070
rect 188286 141068 188292 141070
rect 188356 141068 188362 141132
rect 124029 140994 124095 140997
rect 189758 140994 189764 140996
rect 124029 140992 189764 140994
rect 124029 140936 124034 140992
rect 124090 140936 189764 140992
rect 124029 140934 189764 140936
rect 124029 140931 124095 140934
rect 189758 140932 189764 140934
rect 189828 140932 189834 140996
rect 125409 140858 125475 140861
rect 192334 140858 192340 140860
rect 125409 140856 192340 140858
rect 125409 140800 125414 140856
rect 125470 140800 192340 140856
rect 125409 140798 192340 140800
rect 125409 140795 125475 140798
rect 192334 140796 192340 140798
rect 192404 140796 192410 140860
rect 120574 140524 120580 140588
rect 120644 140586 120650 140588
rect 182265 140586 182331 140589
rect 120644 140584 182331 140586
rect 120644 140528 182270 140584
rect 182326 140528 182331 140584
rect 120644 140526 182331 140528
rect 120644 140524 120650 140526
rect 182265 140523 182331 140526
rect 169753 140450 169819 140453
rect 190678 140450 190684 140452
rect 169753 140448 190684 140450
rect 169753 140392 169758 140448
rect 169814 140392 190684 140448
rect 169753 140390 190684 140392
rect 169753 140387 169819 140390
rect 190678 140388 190684 140390
rect 190748 140388 190754 140452
rect 122373 140314 122439 140317
rect 125225 140314 125291 140317
rect 122373 140312 125291 140314
rect 122373 140256 122378 140312
rect 122434 140256 125230 140312
rect 125286 140256 125291 140312
rect 122373 140254 125291 140256
rect 122373 140251 122439 140254
rect 125225 140251 125291 140254
rect 126278 140252 126284 140316
rect 126348 140314 126354 140316
rect 126697 140314 126763 140317
rect 126348 140312 126763 140314
rect 126348 140256 126702 140312
rect 126758 140256 126763 140312
rect 126348 140254 126763 140256
rect 126348 140252 126354 140254
rect 126697 140251 126763 140254
rect 169937 140314 170003 140317
rect 191281 140314 191347 140317
rect 169937 140312 191347 140314
rect 169937 140256 169942 140312
rect 169998 140256 191286 140312
rect 191342 140256 191347 140312
rect 169937 140254 191347 140256
rect 169937 140251 170003 140254
rect 191281 140251 191347 140254
rect 128905 140178 128971 140181
rect 122790 140176 128971 140178
rect 122790 140120 128910 140176
rect 128966 140120 128971 140176
rect 122790 140118 128971 140120
rect 122598 139980 122604 140044
rect 122668 140042 122674 140044
rect 122790 140042 122850 140118
rect 128905 140115 128971 140118
rect 157057 140178 157123 140181
rect 178718 140178 178724 140180
rect 157057 140176 178724 140178
rect 157057 140120 157062 140176
rect 157118 140120 178724 140176
rect 157057 140118 178724 140120
rect 157057 140115 157123 140118
rect 178718 140116 178724 140118
rect 178788 140116 178794 140180
rect 179045 140178 179111 140181
rect 185853 140180 185919 140181
rect 185853 140178 185900 140180
rect 179045 140176 180810 140178
rect 179045 140120 179050 140176
rect 179106 140120 180810 140176
rect 179045 140118 180810 140120
rect 185808 140176 185900 140178
rect 185808 140120 185858 140176
rect 185808 140118 185900 140120
rect 179045 140115 179111 140118
rect 122668 139982 122850 140042
rect 122668 139980 122674 139982
rect 123518 139980 123524 140044
rect 123588 140042 123594 140044
rect 129181 140042 129247 140045
rect 123588 140040 129247 140042
rect 123588 139984 129186 140040
rect 129242 139984 129247 140040
rect 123588 139982 129247 139984
rect 123588 139980 123594 139982
rect 129181 139979 129247 139982
rect 158529 140042 158595 140045
rect 180006 140042 180012 140044
rect 158529 140040 180012 140042
rect 158529 139984 158534 140040
rect 158590 139984 180012 140040
rect 158529 139982 180012 139984
rect 158529 139979 158595 139982
rect 180006 139980 180012 139982
rect 180076 139980 180082 140044
rect 119838 139844 119844 139908
rect 119908 139906 119914 139908
rect 125041 139906 125107 139909
rect 119908 139904 125107 139906
rect 119908 139848 125046 139904
rect 125102 139848 125107 139904
rect 119908 139846 125107 139848
rect 180750 139906 180810 140118
rect 185853 140116 185900 140118
rect 185964 140116 185970 140180
rect 186221 140178 186287 140181
rect 189022 140178 189028 140180
rect 186221 140176 189028 140178
rect 186221 140120 186226 140176
rect 186282 140120 189028 140176
rect 186221 140118 189028 140120
rect 185853 140115 185919 140116
rect 186221 140115 186287 140118
rect 189022 140116 189028 140118
rect 189092 140116 189098 140180
rect 181621 140044 181687 140045
rect 181621 140042 181668 140044
rect 181576 140040 181668 140042
rect 181576 139984 181626 140040
rect 181576 139982 181668 139984
rect 181621 139980 181668 139982
rect 181732 139980 181738 140044
rect 183461 140042 183527 140045
rect 188654 140042 188660 140044
rect 183461 140040 188660 140042
rect 183461 139984 183466 140040
rect 183522 139984 188660 140040
rect 183461 139982 188660 139984
rect 181621 139979 181687 139980
rect 183461 139979 183527 139982
rect 188654 139980 188660 139982
rect 188724 139980 188730 140044
rect 191966 139906 191972 139908
rect 180750 139846 191972 139906
rect 119908 139844 119914 139846
rect 125041 139843 125107 139846
rect 191966 139844 191972 139846
rect 192036 139844 192042 139908
rect 180149 139770 180215 139773
rect 186221 139770 186287 139773
rect 180149 139768 186287 139770
rect 180149 139712 180154 139768
rect 180210 139712 186226 139768
rect 186282 139712 186287 139768
rect 180149 139710 186287 139712
rect 180149 139707 180215 139710
rect 186221 139707 186287 139710
rect 187734 139708 187740 139772
rect 187804 139770 187810 139772
rect 188705 139770 188771 139773
rect 187804 139768 188771 139770
rect 187804 139712 188710 139768
rect 188766 139712 188771 139768
rect 187804 139710 188771 139712
rect 187804 139708 187810 139710
rect 188705 139707 188771 139710
rect 122046 139572 122052 139636
rect 122116 139634 122122 139636
rect 184013 139634 184079 139637
rect 122116 139632 184079 139634
rect 122116 139576 184018 139632
rect 184074 139576 184079 139632
rect 122116 139574 184079 139576
rect 122116 139572 122122 139574
rect 184013 139571 184079 139574
rect 184657 139634 184723 139637
rect 327717 139634 327783 139637
rect 184657 139632 327783 139634
rect 184657 139576 184662 139632
rect 184718 139576 327722 139632
rect 327778 139576 327783 139632
rect 184657 139574 327783 139576
rect 184657 139571 184723 139574
rect 327717 139571 327783 139574
rect 120758 139436 120764 139500
rect 120828 139498 120834 139500
rect 183829 139498 183895 139501
rect 184381 139498 184447 139501
rect 120828 139496 184447 139498
rect 120828 139440 183834 139496
rect 183890 139440 184386 139496
rect 184442 139440 184447 139496
rect 120828 139438 184447 139440
rect 120828 139436 120834 139438
rect 183829 139435 183895 139438
rect 184381 139435 184447 139438
rect 184565 139498 184631 139501
rect 576117 139498 576183 139501
rect 184565 139496 576183 139498
rect 184565 139440 184570 139496
rect 184626 139440 576122 139496
rect 576178 139440 576183 139496
rect 184565 139438 576183 139440
rect 184565 139435 184631 139438
rect 576117 139435 576183 139438
rect 122414 139300 122420 139364
rect 122484 139362 122490 139364
rect 124489 139362 124555 139365
rect 122484 139360 124555 139362
rect 122484 139304 124494 139360
rect 124550 139304 124555 139360
rect 122484 139302 124555 139304
rect 122484 139300 122490 139302
rect 124489 139299 124555 139302
rect 124806 139300 124812 139364
rect 124876 139362 124882 139364
rect 125501 139362 125567 139365
rect 125961 139362 126027 139365
rect 124876 139360 125567 139362
rect 124876 139304 125506 139360
rect 125562 139304 125567 139360
rect 124876 139302 125567 139304
rect 124876 139300 124882 139302
rect 125501 139299 125567 139302
rect 125734 139360 126027 139362
rect 125734 139304 125966 139360
rect 126022 139304 126027 139360
rect 125734 139302 126027 139304
rect 122189 139090 122255 139093
rect 125734 139090 125794 139302
rect 125961 139299 126027 139302
rect 126145 139362 126211 139365
rect 126462 139362 126468 139364
rect 126145 139360 126468 139362
rect 126145 139304 126150 139360
rect 126206 139304 126468 139360
rect 126145 139302 126468 139304
rect 126145 139299 126211 139302
rect 126462 139300 126468 139302
rect 126532 139300 126538 139364
rect 127617 139362 127683 139365
rect 130009 139362 130075 139365
rect 126838 139360 127683 139362
rect 126838 139304 127622 139360
rect 127678 139304 127683 139360
rect 126838 139302 127683 139304
rect 122189 139088 125794 139090
rect 122189 139032 122194 139088
rect 122250 139032 125794 139088
rect 122189 139030 125794 139032
rect 122189 139027 122255 139030
rect 119797 138954 119863 138957
rect 126838 138954 126898 139302
rect 127617 139299 127683 139302
rect 127758 139360 130075 139362
rect 127758 139304 130014 139360
rect 130070 139304 130075 139360
rect 127758 139302 130075 139304
rect 119797 138952 126898 138954
rect 119797 138896 119802 138952
rect 119858 138896 126898 138952
rect 119797 138894 126898 138896
rect 119797 138891 119863 138894
rect 120809 138818 120875 138821
rect 127758 138818 127818 139302
rect 130009 139299 130075 139302
rect 130326 139300 130332 139364
rect 130396 139362 130402 139364
rect 131021 139362 131087 139365
rect 130396 139360 131087 139362
rect 130396 139304 131026 139360
rect 131082 139304 131087 139360
rect 130396 139302 131087 139304
rect 130396 139300 130402 139302
rect 131021 139299 131087 139302
rect 131798 139300 131804 139364
rect 131868 139362 131874 139364
rect 132217 139362 132283 139365
rect 149605 139362 149671 139365
rect 150985 139364 151051 139365
rect 150934 139362 150940 139364
rect 131868 139360 132283 139362
rect 131868 139304 132222 139360
rect 132278 139304 132283 139360
rect 131868 139302 132283 139304
rect 131868 139300 131874 139302
rect 132217 139299 132283 139302
rect 142110 139360 149671 139362
rect 142110 139304 149610 139360
rect 149666 139304 149671 139360
rect 142110 139302 149671 139304
rect 150894 139302 150940 139362
rect 151004 139360 151051 139364
rect 151046 139304 151051 139360
rect 120809 138816 127818 138818
rect 120809 138760 120814 138816
rect 120870 138760 127818 138816
rect 120809 138758 127818 138760
rect 120809 138755 120875 138758
rect 119654 138620 119660 138684
rect 119724 138682 119730 138684
rect 142110 138682 142170 139302
rect 149605 139299 149671 139302
rect 150934 139300 150940 139302
rect 151004 139300 151051 139304
rect 154798 139300 154804 139364
rect 154868 139362 154874 139364
rect 155217 139362 155283 139365
rect 154868 139360 155283 139362
rect 154868 139304 155222 139360
rect 155278 139304 155283 139360
rect 154868 139302 155283 139304
rect 154868 139300 154874 139302
rect 150985 139299 151051 139300
rect 155217 139299 155283 139302
rect 155350 139300 155356 139364
rect 155420 139362 155426 139364
rect 155769 139362 155835 139365
rect 155420 139360 155835 139362
rect 155420 139304 155774 139360
rect 155830 139304 155835 139360
rect 155420 139302 155835 139304
rect 155420 139300 155426 139302
rect 155769 139299 155835 139302
rect 159214 139300 159220 139364
rect 159284 139362 159290 139364
rect 159541 139362 159607 139365
rect 159284 139360 159607 139362
rect 159284 139304 159546 139360
rect 159602 139304 159607 139360
rect 159284 139302 159607 139304
rect 159284 139300 159290 139302
rect 159541 139299 159607 139302
rect 159817 139362 159883 139365
rect 159950 139362 159956 139364
rect 159817 139360 159956 139362
rect 159817 139304 159822 139360
rect 159878 139304 159956 139360
rect 159817 139302 159956 139304
rect 159817 139299 159883 139302
rect 159950 139300 159956 139302
rect 160020 139300 160026 139364
rect 165337 139362 165403 139365
rect 178861 139362 178927 139365
rect 180149 139362 180215 139365
rect 188245 139362 188311 139365
rect 191097 139362 191163 139365
rect 165337 139360 171150 139362
rect 165337 139304 165342 139360
rect 165398 139304 171150 139360
rect 165337 139302 171150 139304
rect 165337 139299 165403 139302
rect 119724 138622 142170 138682
rect 171090 138682 171150 139302
rect 178861 139360 179890 139362
rect 178861 139304 178866 139360
rect 178922 139304 179890 139360
rect 178861 139302 179890 139304
rect 178861 139299 178927 139302
rect 179830 139090 179890 139302
rect 180149 139360 188311 139362
rect 180149 139304 180154 139360
rect 180210 139304 188250 139360
rect 188306 139304 188311 139360
rect 180149 139302 188311 139304
rect 180149 139299 180215 139302
rect 188245 139299 188311 139302
rect 190410 139360 191163 139362
rect 190410 139304 191102 139360
rect 191158 139304 191163 139360
rect 190410 139302 191163 139304
rect 186865 139226 186931 139229
rect 190410 139226 190470 139302
rect 191097 139299 191163 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 186865 139224 190470 139226
rect 186865 139168 186870 139224
rect 186926 139168 190470 139224
rect 583520 139212 584960 139302
rect 186865 139166 190470 139168
rect 186865 139163 186931 139166
rect 186865 139090 186931 139093
rect 179830 139088 186931 139090
rect 179830 139032 186870 139088
rect 186926 139032 186931 139088
rect 179830 139030 186931 139032
rect 186865 139027 186931 139030
rect 187417 139090 187483 139093
rect 196801 139090 196867 139093
rect 187417 139088 196867 139090
rect 187417 139032 187422 139088
rect 187478 139032 196806 139088
rect 196862 139032 196867 139088
rect 187417 139030 196867 139032
rect 187417 139027 187483 139030
rect 196801 139027 196867 139030
rect 185894 138892 185900 138956
rect 185964 138954 185970 138956
rect 198181 138954 198247 138957
rect 185964 138952 198247 138954
rect 185964 138896 198186 138952
rect 198242 138896 198247 138952
rect 185964 138894 198247 138896
rect 185964 138892 185970 138894
rect 198181 138891 198247 138894
rect 181662 138756 181668 138820
rect 181732 138818 181738 138820
rect 200113 138818 200179 138821
rect 181732 138816 200179 138818
rect 181732 138760 200118 138816
rect 200174 138760 200179 138816
rect 181732 138758 200179 138760
rect 181732 138756 181738 138758
rect 200113 138755 200179 138758
rect 191189 138682 191255 138685
rect 171090 138680 191255 138682
rect 171090 138624 191194 138680
rect 191250 138624 191255 138680
rect 171090 138622 191255 138624
rect 119724 138620 119730 138622
rect 191189 138619 191255 138622
rect 118877 138138 118943 138141
rect 119470 138138 119476 138140
rect 118877 138136 119476 138138
rect 118877 138080 118882 138136
rect 118938 138080 119476 138136
rect 118877 138078 119476 138080
rect 118877 138075 118943 138078
rect 119470 138076 119476 138078
rect 119540 138076 119546 138140
rect 200798 138076 200804 138140
rect 200868 138138 200874 138140
rect 200941 138138 201007 138141
rect 200868 138136 201007 138138
rect 200868 138080 200946 138136
rect 201002 138080 201007 138136
rect 200868 138078 201007 138080
rect 200868 138076 200874 138078
rect 200941 138075 201007 138078
rect 186078 137940 186084 138004
rect 186148 138002 186154 138004
rect 192661 138002 192727 138005
rect 186148 138000 192727 138002
rect 186148 137944 192666 138000
rect 192722 137944 192727 138000
rect 186148 137942 192727 137944
rect 186148 137940 186154 137942
rect 192661 137939 192727 137942
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 122373 132562 122439 132565
rect 122782 132562 122788 132564
rect 122373 132560 122788 132562
rect 122373 132504 122378 132560
rect 122434 132504 122788 132560
rect 122373 132502 122788 132504
rect 122373 132499 122439 132502
rect 122782 132500 122788 132502
rect 122852 132500 122858 132564
rect 122373 132426 122439 132429
rect 122782 132426 122788 132428
rect 122373 132424 122788 132426
rect 122373 132368 122378 132424
rect 122434 132368 122788 132424
rect 122373 132366 122788 132368
rect 122373 132363 122439 132366
rect 122782 132364 122788 132366
rect 122852 132364 122858 132428
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 188654 125564 188660 125628
rect 188724 125626 188730 125628
rect 583526 125626 583586 125838
rect 188724 125566 583586 125626
rect 188724 125564 188730 125566
rect -960 123572 480 123812
rect 122373 122906 122439 122909
rect 122782 122906 122788 122908
rect 122373 122904 122788 122906
rect 122373 122848 122378 122904
rect 122434 122848 122788 122904
rect 122373 122846 122788 122848
rect 122373 122843 122439 122846
rect 122782 122844 122788 122846
rect 122852 122844 122858 122908
rect 122373 122770 122439 122773
rect 122782 122770 122788 122772
rect 122373 122768 122788 122770
rect 122373 122712 122378 122768
rect 122434 122712 122788 122768
rect 122373 122710 122788 122712
rect 122373 122707 122439 122710
rect 122782 122708 122788 122710
rect 122852 122708 122858 122772
rect 122373 113250 122439 113253
rect 122782 113250 122788 113252
rect 122373 113248 122788 113250
rect 122373 113192 122378 113248
rect 122434 113192 122788 113248
rect 122373 113190 122788 113192
rect 122373 113187 122439 113190
rect 122782 113188 122788 113190
rect 122852 113188 122858 113252
rect 122373 113114 122439 113117
rect 122782 113114 122788 113116
rect 122373 113112 122788 113114
rect 122373 113056 122378 113112
rect 122434 113056 122788 113112
rect 122373 113054 122788 113056
rect 122373 113051 122439 113054
rect 122782 113052 122788 113054
rect 122852 113052 122858 113116
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 188286 111828 188292 111892
rect 188356 111890 188362 111892
rect 583526 111890 583586 112646
rect 188356 111830 583586 111890
rect 188356 111828 188362 111830
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 122373 103594 122439 103597
rect 122782 103594 122788 103596
rect 122373 103592 122788 103594
rect 122373 103536 122378 103592
rect 122434 103536 122788 103592
rect 122373 103534 122788 103536
rect 122373 103531 122439 103534
rect 122782 103532 122788 103534
rect 122852 103532 122858 103596
rect 122373 103458 122439 103461
rect 122782 103458 122788 103460
rect 122373 103456 122788 103458
rect 122373 103400 122378 103456
rect 122434 103400 122788 103456
rect 122373 103398 122788 103400
rect 122373 103395 122439 103398
rect 122782 103396 122788 103398
rect 122852 103396 122858 103460
rect 580257 99514 580323 99517
rect 583520 99514 584960 99604
rect 580257 99512 584960 99514
rect 580257 99456 580262 99512
rect 580318 99456 584960 99512
rect 580257 99454 584960 99456
rect 580257 99451 580323 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 120574 96658 120580 96660
rect 6870 96598 120580 96658
rect 120574 96596 120580 96598
rect 120644 96596 120650 96660
rect 122373 93938 122439 93941
rect 122782 93938 122788 93940
rect 122373 93936 122788 93938
rect 122373 93880 122378 93936
rect 122434 93880 122788 93936
rect 122373 93878 122788 93880
rect 122373 93875 122439 93878
rect 122782 93876 122788 93878
rect 122852 93876 122858 93940
rect 122373 93802 122439 93805
rect 122782 93802 122788 93804
rect 122373 93800 122788 93802
rect 122373 93744 122378 93800
rect 122434 93744 122788 93800
rect 122373 93742 122788 93744
rect 122373 93739 122439 93742
rect 122782 93740 122788 93742
rect 122852 93740 122858 93804
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 122373 84282 122439 84285
rect 122782 84282 122788 84284
rect 122373 84280 122788 84282
rect 122373 84224 122378 84280
rect 122434 84224 122788 84280
rect 122373 84222 122788 84224
rect 122373 84219 122439 84222
rect 122782 84220 122788 84222
rect 122852 84220 122858 84284
rect 122373 84146 122439 84149
rect 122782 84146 122788 84148
rect 122373 84144 122788 84146
rect 122373 84088 122378 84144
rect 122434 84088 122788 84144
rect 122373 84086 122788 84088
rect 122373 84083 122439 84086
rect 122782 84084 122788 84086
rect 122852 84084 122858 84148
rect 137134 81636 137140 81700
rect 137204 81698 137210 81700
rect 142286 81698 142292 81700
rect 137204 81638 142292 81698
rect 137204 81636 137210 81638
rect 142286 81636 142292 81638
rect 142356 81636 142362 81700
rect 77293 81562 77359 81565
rect 138238 81562 138244 81564
rect 77293 81560 138244 81562
rect 77293 81504 77298 81560
rect 77354 81504 138244 81560
rect 77293 81502 138244 81504
rect 77293 81499 77359 81502
rect 138238 81500 138244 81502
rect 138308 81500 138314 81564
rect 130510 81228 130516 81292
rect 130580 81290 130586 81292
rect 144678 81290 144684 81292
rect 130580 81230 144684 81290
rect 130580 81228 130586 81230
rect 144678 81228 144684 81230
rect 144748 81228 144754 81292
rect 174118 81228 174124 81292
rect 174188 81290 174194 81292
rect 174854 81290 174860 81292
rect 174188 81230 174860 81290
rect 174188 81228 174194 81230
rect 174854 81228 174860 81230
rect 174924 81228 174930 81292
rect 126830 81092 126836 81156
rect 126900 81154 126906 81156
rect 145046 81154 145052 81156
rect 126900 81094 145052 81154
rect 126900 81092 126906 81094
rect 145046 81092 145052 81094
rect 145116 81092 145122 81156
rect 150014 81092 150020 81156
rect 150084 81154 150090 81156
rect 158662 81154 158668 81156
rect 150084 81094 158668 81154
rect 150084 81092 150090 81094
rect 158662 81092 158668 81094
rect 158732 81092 158738 81156
rect 171358 81092 171364 81156
rect 171428 81154 171434 81156
rect 191281 81154 191347 81157
rect 171428 81152 191347 81154
rect 171428 81096 191286 81152
rect 191342 81096 191347 81152
rect 171428 81094 191347 81096
rect 171428 81092 171434 81094
rect 191281 81091 191347 81094
rect 125174 80956 125180 81020
rect 125244 81018 125250 81020
rect 144494 81018 144500 81020
rect 125244 80958 144500 81018
rect 125244 80956 125250 80958
rect 144494 80956 144500 80958
rect 144564 80956 144570 81020
rect 159398 80956 159404 81020
rect 159468 81018 159474 81020
rect 180006 81018 180012 81020
rect 159468 80958 180012 81018
rect 159468 80956 159474 80958
rect 180006 80956 180012 80958
rect 180076 80956 180082 81020
rect 126646 80820 126652 80884
rect 126716 80882 126722 80884
rect 146334 80882 146340 80884
rect 126716 80822 146340 80882
rect 126716 80820 126722 80822
rect 146334 80820 146340 80822
rect 146404 80820 146410 80884
rect 162526 80820 162532 80884
rect 162596 80882 162602 80884
rect 168414 80882 168420 80884
rect 162596 80822 168420 80882
rect 162596 80820 162602 80822
rect 168414 80820 168420 80822
rect 168484 80820 168490 80884
rect 170622 80820 170628 80884
rect 170692 80882 170698 80884
rect 193949 80882 194015 80885
rect 170692 80880 194015 80882
rect 170692 80824 193954 80880
rect 194010 80824 194015 80880
rect 170692 80822 194015 80824
rect 170692 80820 170698 80822
rect 193949 80819 194015 80822
rect 145966 80746 145972 80748
rect 128310 80686 145972 80746
rect 126278 80412 126284 80476
rect 126348 80474 126354 80476
rect 128310 80474 128370 80686
rect 145966 80684 145972 80686
rect 146036 80684 146042 80748
rect 167678 80684 167684 80748
rect 167748 80746 167754 80748
rect 177246 80746 177252 80748
rect 167748 80686 177252 80746
rect 167748 80684 167754 80686
rect 177246 80684 177252 80686
rect 177316 80684 177322 80748
rect 177430 80684 177436 80748
rect 177500 80746 177506 80748
rect 177757 80746 177823 80749
rect 177500 80744 177823 80746
rect 177500 80688 177762 80744
rect 177818 80688 177823 80744
rect 177500 80686 177823 80688
rect 177500 80684 177506 80686
rect 177757 80683 177823 80686
rect 177941 80746 178007 80749
rect 178401 80746 178467 80749
rect 182541 80748 182607 80749
rect 178534 80746 178540 80748
rect 177941 80744 178050 80746
rect 177941 80688 177946 80744
rect 178002 80688 178050 80744
rect 177941 80683 178050 80688
rect 178401 80744 178540 80746
rect 178401 80688 178406 80744
rect 178462 80688 178540 80744
rect 178401 80686 178540 80688
rect 178401 80683 178467 80686
rect 178534 80684 178540 80686
rect 178604 80684 178610 80748
rect 182541 80744 182588 80748
rect 182652 80746 182658 80748
rect 206461 80746 206527 80749
rect 182541 80688 182546 80744
rect 182541 80684 182588 80688
rect 182652 80686 182698 80746
rect 186270 80744 206527 80746
rect 186270 80688 206466 80744
rect 206522 80688 206527 80744
rect 186270 80686 206527 80688
rect 182652 80684 182658 80686
rect 182541 80683 182607 80684
rect 130694 80548 130700 80612
rect 130764 80610 130770 80612
rect 143574 80610 143580 80612
rect 130764 80550 143580 80610
rect 130764 80548 130770 80550
rect 143574 80548 143580 80550
rect 143644 80548 143650 80612
rect 175222 80548 175228 80612
rect 175292 80610 175298 80612
rect 177990 80610 178050 80683
rect 175292 80550 178050 80610
rect 178125 80610 178191 80613
rect 186270 80610 186330 80686
rect 206461 80683 206527 80686
rect 178125 80608 186330 80610
rect 178125 80552 178130 80608
rect 178186 80552 186330 80608
rect 178125 80550 186330 80552
rect 175292 80548 175298 80550
rect 178125 80547 178191 80550
rect 131849 80476 131915 80477
rect 131798 80474 131804 80476
rect 126348 80414 128370 80474
rect 131758 80414 131804 80474
rect 131868 80472 131915 80476
rect 131910 80416 131915 80472
rect 126348 80412 126354 80414
rect 131798 80412 131804 80414
rect 131868 80412 131915 80416
rect 131849 80411 131915 80412
rect 132125 80474 132191 80477
rect 135662 80474 135668 80476
rect 132125 80472 135668 80474
rect 132125 80416 132130 80472
rect 132186 80416 135668 80472
rect 132125 80414 135668 80416
rect 132125 80411 132191 80414
rect 135662 80412 135668 80414
rect 135732 80412 135738 80476
rect 148542 80474 148548 80476
rect 135854 80414 148548 80474
rect 123518 80276 123524 80340
rect 123588 80338 123594 80340
rect 124121 80338 124187 80341
rect 123588 80336 124187 80338
rect 123588 80280 124126 80336
rect 124182 80280 124187 80336
rect 123588 80278 124187 80280
rect 123588 80276 123594 80278
rect 124121 80275 124187 80278
rect 120533 80202 120599 80205
rect 135854 80202 135914 80414
rect 148542 80412 148548 80414
rect 148612 80412 148618 80476
rect 162710 80474 162716 80476
rect 161982 80414 162716 80474
rect 149462 80276 149468 80340
rect 149532 80338 149538 80340
rect 160502 80338 160508 80340
rect 149532 80278 160508 80338
rect 149532 80276 149538 80278
rect 160502 80276 160508 80278
rect 160572 80276 160578 80340
rect 120533 80200 135914 80202
rect 120533 80144 120538 80200
rect 120594 80144 135914 80200
rect 120533 80142 135914 80144
rect 135992 80142 137386 80202
rect 120533 80139 120599 80142
rect 134374 80066 134380 80068
rect 133922 80006 134380 80066
rect 132815 79964 132881 79967
rect 133183 79964 133249 79967
rect 133551 79964 133617 79967
rect 132815 79962 132924 79964
rect 131757 79930 131823 79933
rect 132815 79930 132820 79962
rect 131757 79928 132820 79930
rect 131757 79872 131762 79928
rect 131818 79906 132820 79928
rect 132876 79932 132924 79962
rect 133183 79962 133292 79964
rect 132876 79906 132908 79932
rect 131818 79872 132908 79906
rect 131757 79870 132908 79872
rect 131757 79867 131823 79870
rect 132902 79868 132908 79870
rect 132972 79868 132978 79932
rect 133183 79906 133188 79962
rect 133244 79932 133292 79962
rect 133551 79962 133660 79964
rect 133244 79906 133276 79932
rect 133183 79901 133276 79906
rect 133232 79870 133276 79901
rect 133270 79868 133276 79870
rect 133340 79868 133346 79932
rect 133551 79906 133556 79962
rect 133612 79932 133660 79962
rect 133922 79933 133982 80006
rect 134374 80004 134380 80006
rect 134444 80004 134450 80068
rect 135110 80004 135116 80068
rect 135180 80066 135186 80068
rect 135180 80004 135224 80066
rect 135662 80004 135668 80068
rect 135732 80066 135738 80068
rect 135992 80066 136052 80142
rect 135732 80006 136052 80066
rect 137326 80066 137386 80142
rect 139894 80140 139900 80204
rect 139964 80202 139970 80204
rect 139964 80142 147644 80202
rect 139964 80140 139970 80142
rect 137326 80006 138030 80066
rect 135732 80004 135738 80006
rect 135164 79933 135224 80004
rect 137139 79964 137205 79967
rect 137139 79962 137262 79964
rect 133612 79906 133644 79932
rect 133551 79901 133644 79906
rect 133600 79870 133644 79901
rect 133638 79868 133644 79870
rect 133708 79868 133714 79932
rect 133919 79928 133985 79933
rect 133919 79872 133924 79928
rect 133980 79872 133985 79928
rect 133919 79867 133985 79872
rect 134287 79930 134353 79933
rect 134558 79930 134564 79932
rect 134287 79928 134564 79930
rect 134287 79872 134292 79928
rect 134348 79872 134564 79928
rect 134287 79870 134564 79872
rect 134287 79867 134353 79870
rect 134558 79868 134564 79870
rect 134628 79868 134634 79932
rect 135164 79928 135273 79933
rect 135164 79872 135212 79928
rect 135268 79872 135273 79928
rect 135164 79870 135273 79872
rect 135207 79867 135273 79870
rect 136214 79868 136220 79932
rect 136284 79930 136290 79932
rect 136495 79930 136561 79933
rect 136771 79932 136837 79933
rect 137139 79932 137144 79962
rect 137200 79932 137262 79962
rect 137970 79933 138030 80006
rect 140078 80004 140084 80068
rect 140148 80004 140154 80068
rect 140814 80004 140820 80068
rect 140884 80066 140890 80068
rect 140884 80006 141112 80066
rect 140884 80004 140890 80006
rect 138427 79962 138493 79967
rect 136766 79930 136772 79932
rect 136284 79928 136561 79930
rect 136284 79872 136500 79928
rect 136556 79872 136561 79928
rect 136284 79870 136561 79872
rect 136680 79870 136772 79930
rect 136284 79868 136290 79870
rect 136495 79867 136561 79870
rect 136766 79868 136772 79870
rect 136836 79868 136842 79932
rect 137134 79868 137140 79932
rect 137204 79904 137262 79932
rect 137323 79930 137389 79933
rect 137686 79930 137692 79932
rect 137323 79928 137692 79930
rect 137204 79868 137210 79904
rect 137323 79872 137328 79928
rect 137384 79872 137692 79928
rect 137323 79870 137692 79872
rect 136771 79867 136837 79868
rect 137323 79867 137389 79870
rect 137686 79868 137692 79870
rect 137756 79868 137762 79932
rect 137967 79928 138033 79933
rect 137967 79872 137972 79928
rect 138028 79872 138033 79928
rect 137967 79867 138033 79872
rect 138238 79868 138244 79932
rect 138308 79930 138314 79932
rect 138427 79930 138432 79962
rect 138308 79906 138432 79930
rect 138488 79906 138493 79962
rect 138308 79901 138493 79906
rect 138703 79964 138769 79967
rect 138703 79962 138812 79964
rect 138703 79906 138708 79962
rect 138764 79932 138812 79962
rect 140086 79933 140146 80004
rect 140359 79964 140425 79967
rect 140316 79962 140425 79964
rect 138764 79906 138796 79932
rect 138703 79901 138796 79906
rect 138308 79870 138490 79901
rect 138752 79870 138796 79901
rect 138308 79868 138314 79870
rect 138790 79868 138796 79870
rect 138860 79868 138866 79932
rect 138974 79868 138980 79932
rect 139044 79930 139050 79932
rect 139255 79930 139321 79933
rect 139044 79928 139321 79930
rect 139044 79872 139260 79928
rect 139316 79872 139321 79928
rect 139044 79870 139321 79872
rect 139044 79868 139050 79870
rect 139212 79867 139321 79870
rect 140083 79930 140149 79933
rect 140316 79932 140364 79962
rect 140083 79928 140192 79930
rect 140083 79872 140088 79928
rect 140144 79872 140192 79928
rect 140083 79867 140192 79872
rect 140262 79868 140268 79932
rect 140332 79906 140364 79932
rect 140420 79906 140425 79962
rect 140332 79901 140425 79906
rect 140543 79964 140609 79967
rect 140543 79962 140652 79964
rect 140543 79906 140548 79962
rect 140604 79930 140652 79962
rect 140604 79906 140882 79930
rect 140543 79901 140882 79906
rect 140332 79870 140376 79901
rect 140592 79870 140882 79901
rect 140332 79868 140338 79870
rect 116393 79794 116459 79797
rect 116393 79792 138030 79794
rect 116393 79736 116398 79792
rect 116454 79736 138030 79792
rect 116393 79734 138030 79736
rect 116393 79731 116459 79734
rect 131246 79596 131252 79660
rect 131316 79658 131322 79660
rect 131614 79658 131620 79660
rect 131316 79598 131620 79658
rect 131316 79596 131322 79598
rect 131614 79596 131620 79598
rect 131684 79658 131690 79660
rect 132217 79658 132283 79661
rect 131684 79656 132283 79658
rect 131684 79600 132222 79656
rect 132278 79600 132283 79656
rect 131684 79598 132283 79600
rect 131684 79596 131690 79598
rect 132217 79595 132283 79598
rect 133321 79658 133387 79661
rect 134241 79660 134307 79661
rect 133454 79658 133460 79660
rect 133321 79656 133460 79658
rect 133321 79600 133326 79656
rect 133382 79600 133460 79656
rect 133321 79598 133460 79600
rect 133321 79595 133387 79598
rect 133454 79596 133460 79598
rect 133524 79596 133530 79660
rect 134190 79658 134196 79660
rect 134114 79598 134196 79658
rect 134260 79658 134307 79660
rect 135161 79658 135227 79661
rect 134260 79656 135227 79658
rect 134302 79600 135166 79656
rect 135222 79600 135227 79656
rect 134190 79596 134196 79598
rect 134260 79598 135227 79600
rect 134260 79596 134307 79598
rect 134241 79595 134307 79596
rect 135161 79595 135227 79598
rect 135713 79658 135779 79661
rect 135897 79658 135963 79661
rect 136030 79658 136036 79660
rect 135713 79656 136036 79658
rect 135713 79600 135718 79656
rect 135774 79600 135902 79656
rect 135958 79600 136036 79656
rect 135713 79598 136036 79600
rect 135713 79595 135779 79598
rect 135897 79595 135963 79598
rect 136030 79596 136036 79598
rect 136100 79596 136106 79660
rect 136582 79596 136588 79660
rect 136652 79658 136658 79660
rect 136725 79658 136791 79661
rect 137001 79658 137067 79661
rect 136652 79656 137067 79658
rect 136652 79600 136730 79656
rect 136786 79600 137006 79656
rect 137062 79600 137067 79656
rect 136652 79598 137067 79600
rect 136652 79596 136658 79598
rect 136725 79595 136791 79598
rect 137001 79595 137067 79598
rect 137134 79596 137140 79660
rect 137204 79658 137210 79660
rect 137369 79658 137435 79661
rect 137204 79656 137435 79658
rect 137204 79600 137374 79656
rect 137430 79600 137435 79656
rect 137204 79598 137435 79600
rect 137204 79596 137210 79598
rect 137369 79595 137435 79598
rect 124806 79460 124812 79524
rect 124876 79522 124882 79524
rect 130837 79522 130903 79525
rect 132217 79522 132283 79525
rect 124876 79520 132283 79522
rect 124876 79464 130842 79520
rect 130898 79464 132222 79520
rect 132278 79464 132283 79520
rect 124876 79462 132283 79464
rect 124876 79460 124882 79462
rect 130837 79459 130903 79462
rect 132217 79459 132283 79462
rect 133597 79522 133663 79525
rect 135529 79524 135595 79525
rect 134742 79522 134748 79524
rect 133597 79520 134748 79522
rect 133597 79464 133602 79520
rect 133658 79464 134748 79520
rect 133597 79462 134748 79464
rect 133597 79459 133663 79462
rect 134742 79460 134748 79462
rect 134812 79460 134818 79524
rect 135478 79522 135484 79524
rect 135438 79462 135484 79522
rect 135548 79520 135595 79524
rect 135590 79464 135595 79520
rect 135478 79460 135484 79462
rect 135548 79460 135595 79464
rect 135529 79459 135595 79460
rect 135713 79522 135779 79525
rect 135846 79522 135852 79524
rect 135713 79520 135852 79522
rect 135713 79464 135718 79520
rect 135774 79464 135852 79520
rect 135713 79462 135852 79464
rect 135713 79459 135779 79462
rect 135846 79460 135852 79462
rect 135916 79460 135922 79524
rect 137001 79522 137067 79525
rect 137318 79522 137324 79524
rect 137001 79520 137324 79522
rect 137001 79464 137006 79520
rect 137062 79464 137324 79520
rect 137001 79462 137324 79464
rect 137001 79459 137067 79462
rect 137318 79460 137324 79462
rect 137388 79460 137394 79524
rect 137502 79460 137508 79524
rect 137572 79522 137578 79524
rect 137645 79522 137711 79525
rect 137572 79520 137711 79522
rect 137572 79464 137650 79520
rect 137706 79464 137711 79520
rect 137572 79462 137711 79464
rect 137970 79522 138030 79734
rect 138238 79732 138244 79796
rect 138308 79794 138314 79796
rect 138519 79794 138585 79797
rect 138308 79792 138585 79794
rect 138308 79736 138524 79792
rect 138580 79736 138585 79792
rect 138308 79734 138585 79736
rect 138308 79732 138314 79734
rect 138519 79731 138585 79734
rect 139212 79661 139272 79867
rect 140132 79797 140192 79867
rect 139531 79796 139597 79797
rect 139526 79794 139532 79796
rect 139440 79734 139532 79794
rect 139526 79732 139532 79734
rect 139596 79732 139602 79796
rect 140129 79792 140195 79797
rect 140589 79796 140655 79797
rect 140589 79794 140636 79796
rect 140129 79736 140134 79792
rect 140190 79736 140195 79792
rect 139531 79731 139597 79732
rect 140129 79731 140195 79736
rect 140544 79792 140636 79794
rect 140544 79736 140594 79792
rect 140544 79734 140636 79736
rect 140589 79732 140636 79734
rect 140700 79732 140706 79796
rect 140589 79731 140655 79732
rect 138473 79658 138539 79661
rect 138606 79658 138612 79660
rect 138473 79656 138612 79658
rect 138473 79600 138478 79656
rect 138534 79600 138612 79656
rect 138473 79598 138612 79600
rect 138473 79595 138539 79598
rect 138606 79596 138612 79598
rect 138676 79596 138682 79660
rect 139209 79656 139275 79661
rect 139209 79600 139214 79656
rect 139270 79600 139275 79656
rect 139209 79595 139275 79600
rect 139342 79596 139348 79660
rect 139412 79658 139418 79660
rect 140221 79658 140287 79661
rect 139412 79656 140287 79658
rect 139412 79600 140226 79656
rect 140282 79600 140287 79656
rect 139412 79598 140287 79600
rect 139412 79596 139418 79598
rect 140221 79595 140287 79598
rect 140497 79658 140563 79661
rect 140822 79658 140882 79870
rect 140497 79656 140882 79658
rect 140497 79600 140502 79656
rect 140558 79600 140882 79656
rect 140497 79598 140882 79600
rect 141052 79658 141112 80006
rect 144494 80004 144500 80068
rect 144564 80066 144570 80068
rect 144564 80006 144746 80066
rect 144564 80004 144570 80006
rect 142659 79962 142725 79967
rect 141182 79868 141188 79932
rect 141252 79930 141258 79932
rect 142015 79930 142081 79933
rect 141252 79928 142081 79930
rect 141252 79872 142020 79928
rect 142076 79872 142081 79928
rect 142659 79906 142664 79962
rect 142720 79930 142725 79962
rect 143027 79962 143093 79967
rect 142838 79930 142844 79932
rect 142720 79906 142844 79930
rect 142659 79901 142844 79906
rect 141252 79870 142081 79872
rect 142662 79870 142844 79901
rect 141252 79868 141258 79870
rect 142015 79867 142081 79870
rect 142838 79868 142844 79870
rect 142908 79868 142914 79932
rect 143027 79906 143032 79962
rect 143088 79930 143093 79962
rect 144686 79933 144746 80006
rect 146702 80004 146708 80068
rect 146772 80066 146778 80068
rect 147584 80066 147644 80142
rect 148358 80140 148364 80204
rect 148428 80202 148434 80204
rect 149094 80202 149100 80204
rect 148428 80142 149100 80202
rect 148428 80140 148434 80142
rect 149094 80140 149100 80142
rect 149164 80140 149170 80204
rect 149278 80140 149284 80204
rect 149348 80202 149354 80204
rect 151118 80202 151124 80204
rect 149348 80142 150450 80202
rect 149348 80140 149354 80142
rect 146772 80006 146954 80066
rect 147584 80006 149162 80066
rect 146772 80004 146778 80006
rect 146155 79962 146221 79967
rect 143763 79932 143829 79933
rect 144499 79932 144565 79933
rect 143206 79930 143212 79932
rect 143088 79906 143212 79930
rect 143027 79901 143212 79906
rect 143030 79870 143212 79901
rect 143206 79868 143212 79870
rect 143276 79868 143282 79932
rect 143758 79930 143764 79932
rect 143672 79870 143764 79930
rect 143758 79868 143764 79870
rect 143828 79868 143834 79932
rect 144494 79930 144500 79932
rect 144408 79870 144500 79930
rect 144494 79868 144500 79870
rect 144564 79868 144570 79932
rect 144683 79928 144749 79933
rect 144683 79872 144688 79928
rect 144744 79872 144749 79928
rect 143763 79867 143829 79868
rect 144499 79867 144565 79868
rect 144683 79867 144749 79872
rect 145143 79930 145209 79933
rect 145143 79928 145252 79930
rect 145143 79872 145148 79928
rect 145204 79872 145252 79928
rect 145143 79867 145252 79872
rect 145414 79868 145420 79932
rect 145484 79930 145490 79932
rect 146155 79930 146160 79962
rect 145484 79906 146160 79930
rect 146216 79906 146221 79962
rect 146894 79933 146954 80006
rect 147351 79964 147417 79967
rect 147351 79962 147460 79964
rect 145484 79901 146221 79906
rect 145484 79870 146218 79901
rect 145484 79868 145490 79870
rect 146334 79868 146340 79932
rect 146404 79930 146410 79932
rect 146404 79899 146632 79930
rect 146891 79928 146957 79933
rect 146404 79894 146681 79899
rect 146404 79870 146620 79894
rect 146404 79868 146410 79870
rect 141739 79792 141805 79797
rect 141739 79736 141744 79792
rect 141800 79736 141805 79792
rect 141739 79731 141805 79736
rect 142843 79794 142909 79797
rect 143022 79794 143028 79796
rect 142843 79792 143028 79794
rect 142843 79736 142848 79792
rect 142904 79736 143028 79792
rect 142843 79734 143028 79736
rect 142843 79731 142909 79734
rect 143022 79732 143028 79734
rect 143092 79732 143098 79796
rect 143625 79794 143691 79797
rect 144407 79794 144473 79797
rect 144678 79794 144684 79796
rect 143625 79792 144684 79794
rect 143625 79736 143630 79792
rect 143686 79736 144412 79792
rect 144468 79736 144684 79792
rect 143625 79734 144684 79736
rect 143625 79731 143691 79734
rect 144407 79731 144473 79734
rect 144678 79732 144684 79734
rect 144748 79732 144754 79796
rect 141742 79658 141802 79731
rect 141052 79598 141802 79658
rect 142705 79658 142771 79661
rect 143165 79658 143231 79661
rect 142705 79656 143231 79658
rect 142705 79600 142710 79656
rect 142766 79600 143170 79656
rect 143226 79600 143231 79656
rect 142705 79598 143231 79600
rect 140497 79595 140563 79598
rect 142705 79595 142771 79598
rect 143165 79595 143231 79598
rect 143574 79596 143580 79660
rect 143644 79658 143650 79660
rect 143809 79658 143875 79661
rect 143644 79656 143875 79658
rect 143644 79600 143814 79656
rect 143870 79600 143875 79656
rect 143644 79598 143875 79600
rect 145192 79658 145252 79867
rect 146572 79838 146620 79870
rect 146676 79838 146681 79894
rect 146891 79872 146896 79928
rect 146952 79872 146957 79928
rect 147351 79906 147356 79962
rect 147412 79932 147460 79962
rect 147627 79932 147693 79933
rect 147995 79932 148061 79933
rect 147412 79906 147444 79932
rect 147351 79901 147444 79906
rect 146891 79867 146957 79872
rect 147400 79870 147444 79901
rect 147438 79868 147444 79870
rect 147508 79868 147514 79932
rect 147622 79868 147628 79932
rect 147692 79930 147698 79932
rect 147990 79930 147996 79932
rect 147692 79870 147784 79930
rect 147904 79870 147996 79930
rect 147692 79868 147698 79870
rect 147990 79868 147996 79870
rect 148060 79868 148066 79932
rect 148179 79894 148245 79899
rect 147627 79867 147693 79868
rect 147995 79867 148061 79868
rect 146572 79836 146681 79838
rect 146615 79833 146681 79836
rect 148179 79838 148184 79894
rect 148240 79838 148245 79894
rect 148358 79868 148364 79932
rect 148428 79930 148434 79932
rect 148639 79930 148705 79933
rect 148428 79928 148705 79930
rect 148428 79872 148644 79928
rect 148700 79872 148705 79928
rect 148428 79870 148705 79872
rect 148428 79868 148434 79870
rect 148639 79867 148705 79870
rect 148179 79833 148245 79838
rect 145327 79794 145393 79797
rect 146201 79794 146267 79797
rect 145327 79792 146267 79794
rect 145327 79736 145332 79792
rect 145388 79736 146206 79792
rect 146262 79736 146267 79792
rect 145327 79734 146267 79736
rect 145327 79731 145393 79734
rect 146201 79731 146267 79734
rect 146886 79732 146892 79796
rect 146956 79794 146962 79796
rect 147397 79794 147463 79797
rect 146956 79792 147463 79794
rect 146956 79736 147402 79792
rect 147458 79736 147463 79792
rect 146956 79734 147463 79736
rect 146956 79732 146962 79734
rect 147397 79731 147463 79734
rect 148182 79661 148242 79833
rect 148869 79792 148935 79797
rect 148869 79736 148874 79792
rect 148930 79736 148935 79792
rect 148869 79731 148935 79736
rect 145373 79658 145439 79661
rect 145192 79656 145439 79658
rect 145192 79600 145378 79656
rect 145434 79600 145439 79656
rect 145192 79598 145439 79600
rect 143644 79596 143650 79598
rect 143809 79595 143875 79598
rect 145373 79595 145439 79598
rect 145598 79596 145604 79660
rect 145668 79658 145674 79660
rect 147857 79658 147923 79661
rect 145668 79656 147923 79658
rect 145668 79600 147862 79656
rect 147918 79600 147923 79656
rect 145668 79598 147923 79600
rect 145668 79596 145674 79598
rect 147857 79595 147923 79598
rect 148133 79656 148242 79661
rect 148133 79600 148138 79656
rect 148194 79600 148242 79656
rect 148133 79598 148242 79600
rect 148133 79595 148199 79598
rect 148358 79596 148364 79660
rect 148428 79658 148434 79660
rect 148872 79658 148932 79731
rect 148428 79598 148932 79658
rect 149102 79658 149162 80006
rect 150198 80004 150204 80068
rect 150268 80004 150274 80068
rect 149375 79964 149441 79967
rect 149375 79962 149484 79964
rect 149375 79906 149380 79962
rect 149436 79906 149484 79962
rect 150019 79962 150085 79967
rect 149375 79901 149484 79906
rect 149424 79797 149484 79901
rect 149830 79868 149836 79932
rect 149900 79930 149906 79932
rect 150019 79930 150024 79962
rect 149900 79906 150024 79930
rect 150080 79906 150085 79962
rect 150206 79933 150266 80004
rect 150390 79967 150450 80142
rect 150942 80142 151124 80202
rect 150942 80066 151002 80142
rect 151118 80140 151124 80142
rect 151188 80140 151194 80204
rect 156454 80140 156460 80204
rect 156524 80202 156530 80204
rect 156524 80142 157074 80202
rect 156524 80140 156530 80142
rect 150896 80006 151002 80066
rect 150896 79967 150956 80006
rect 151118 80004 151124 80068
rect 151188 80066 151194 80068
rect 151670 80066 151676 80068
rect 151188 80006 151324 80066
rect 151188 80004 151194 80006
rect 150387 79962 150453 79967
rect 149900 79901 150085 79906
rect 150203 79928 150269 79933
rect 149900 79870 150082 79901
rect 150203 79872 150208 79928
rect 150264 79872 150269 79928
rect 150387 79906 150392 79962
rect 150448 79906 150453 79962
rect 150847 79962 150956 79967
rect 150387 79901 150453 79906
rect 150571 79928 150637 79933
rect 149900 79868 149906 79870
rect 150203 79867 150269 79872
rect 150571 79872 150576 79928
rect 150632 79872 150637 79928
rect 150847 79906 150852 79962
rect 150908 79906 150956 79962
rect 151264 79967 151324 80006
rect 151494 80006 151676 80066
rect 151264 79962 151373 79967
rect 150847 79901 150956 79906
rect 150571 79867 150637 79872
rect 150574 79797 150634 79867
rect 150896 79797 150956 79901
rect 151123 79928 151189 79933
rect 151123 79872 151128 79928
rect 151184 79872 151189 79928
rect 151264 79906 151312 79962
rect 151368 79906 151373 79962
rect 151264 79904 151373 79906
rect 151307 79901 151373 79904
rect 151494 79930 151554 80006
rect 151670 80004 151676 80006
rect 151740 80004 151746 80068
rect 155350 80004 155356 80068
rect 155420 80066 155426 80068
rect 155420 80006 155878 80066
rect 155420 80004 155426 80006
rect 152595 79962 152661 79967
rect 154711 79964 154777 79967
rect 151767 79930 151833 79933
rect 151494 79928 151833 79930
rect 151123 79867 151189 79872
rect 151494 79872 151772 79928
rect 151828 79872 151833 79928
rect 151494 79870 151833 79872
rect 151767 79867 151833 79870
rect 152406 79868 152412 79932
rect 152476 79930 152482 79932
rect 152595 79930 152600 79962
rect 152476 79906 152600 79930
rect 152656 79906 152661 79962
rect 154530 79962 154777 79964
rect 152476 79901 152661 79906
rect 152476 79870 152658 79901
rect 152476 79868 152482 79870
rect 152774 79868 152780 79932
rect 152844 79930 152850 79932
rect 153607 79930 153673 79933
rect 154246 79930 154252 79932
rect 152844 79870 152938 79930
rect 153607 79928 154252 79930
rect 153607 79872 153612 79928
rect 153668 79872 154252 79928
rect 153607 79870 154252 79872
rect 152844 79868 152850 79870
rect 149421 79792 149487 79797
rect 149421 79736 149426 79792
rect 149482 79736 149487 79792
rect 149421 79731 149487 79736
rect 150574 79792 150683 79797
rect 150574 79736 150622 79792
rect 150678 79736 150683 79792
rect 150574 79734 150683 79736
rect 150617 79731 150683 79734
rect 150893 79792 150959 79797
rect 150893 79736 150898 79792
rect 150954 79736 150959 79792
rect 150893 79731 150959 79736
rect 151126 79794 151186 79867
rect 152779 79838 152784 79868
rect 152840 79838 152845 79868
rect 153607 79867 153673 79870
rect 154246 79868 154252 79870
rect 154316 79868 154322 79932
rect 154530 79906 154716 79962
rect 154772 79906 154777 79962
rect 154530 79904 154777 79906
rect 152779 79833 152845 79838
rect 151261 79796 151327 79797
rect 151261 79794 151308 79796
rect 151126 79792 151308 79794
rect 151372 79794 151378 79796
rect 151126 79736 151266 79792
rect 151126 79734 151308 79736
rect 151261 79732 151308 79734
rect 151372 79734 151454 79794
rect 151675 79792 151741 79797
rect 151675 79736 151680 79792
rect 151736 79736 151741 79792
rect 151372 79732 151378 79734
rect 151261 79731 151327 79732
rect 151675 79731 151741 79736
rect 151854 79732 151860 79796
rect 151924 79794 151930 79796
rect 152227 79794 152293 79797
rect 151924 79792 152293 79794
rect 151924 79736 152232 79792
rect 152288 79736 152293 79792
rect 151924 79734 152293 79736
rect 151924 79732 151930 79734
rect 152227 79731 152293 79734
rect 151678 79661 151738 79731
rect 149789 79658 149855 79661
rect 150065 79658 150131 79661
rect 149102 79656 150131 79658
rect 149102 79600 149794 79656
rect 149850 79600 150070 79656
rect 150126 79600 150131 79656
rect 149102 79598 150131 79600
rect 148428 79596 148434 79598
rect 149789 79595 149855 79598
rect 150065 79595 150131 79598
rect 150934 79596 150940 79660
rect 151004 79658 151010 79660
rect 151678 79658 151787 79661
rect 152457 79658 152523 79661
rect 152590 79658 152596 79660
rect 151004 79656 151868 79658
rect 151004 79600 151726 79656
rect 151782 79600 151868 79656
rect 151004 79598 151868 79600
rect 152457 79656 152596 79658
rect 152457 79600 152462 79656
rect 152518 79600 152596 79656
rect 152457 79598 152596 79600
rect 151004 79596 151010 79598
rect 151721 79595 151787 79598
rect 152457 79595 152523 79598
rect 152590 79596 152596 79598
rect 152660 79596 152666 79660
rect 152782 79658 152842 79833
rect 153878 79732 153884 79796
rect 153948 79794 153954 79796
rect 154297 79794 154363 79797
rect 153948 79792 154363 79794
rect 153948 79736 154302 79792
rect 154358 79736 154363 79792
rect 153948 79734 154363 79736
rect 154530 79794 154590 79904
rect 154711 79901 154777 79904
rect 155079 79964 155145 79967
rect 155079 79962 155188 79964
rect 155079 79906 155084 79962
rect 155140 79930 155188 79962
rect 155818 79933 155878 80006
rect 156091 79962 156157 79967
rect 155350 79930 155356 79932
rect 155140 79906 155356 79930
rect 155079 79901 155356 79906
rect 155128 79870 155356 79901
rect 155350 79868 155356 79870
rect 155420 79868 155426 79932
rect 155631 79930 155697 79933
rect 155815 79930 155881 79933
rect 155631 79928 155740 79930
rect 155631 79872 155636 79928
rect 155692 79872 155740 79928
rect 155631 79867 155740 79872
rect 155815 79928 155924 79930
rect 155815 79872 155820 79928
rect 155876 79872 155924 79928
rect 156091 79906 156096 79962
rect 156152 79906 156157 79962
rect 156459 79962 156525 79967
rect 156459 79932 156464 79962
rect 156520 79932 156525 79962
rect 156091 79901 156157 79906
rect 155815 79867 155924 79872
rect 154895 79828 154961 79831
rect 154895 79826 155004 79828
rect 154530 79734 154682 79794
rect 154895 79770 154900 79826
rect 154956 79794 155004 79826
rect 155125 79794 155191 79797
rect 154956 79792 155191 79794
rect 154956 79770 155130 79792
rect 154895 79765 155130 79770
rect 154944 79736 155130 79765
rect 155186 79736 155191 79792
rect 154944 79734 155191 79736
rect 153948 79732 153954 79734
rect 154297 79731 154363 79734
rect 152917 79658 152983 79661
rect 152782 79656 152983 79658
rect 152782 79600 152922 79656
rect 152978 79600 152983 79656
rect 152782 79598 152983 79600
rect 152917 79595 152983 79598
rect 153837 79658 153903 79661
rect 154481 79658 154547 79661
rect 153837 79656 154547 79658
rect 153837 79600 153842 79656
rect 153898 79600 154486 79656
rect 154542 79600 154547 79656
rect 153837 79598 154547 79600
rect 153837 79595 153903 79598
rect 154481 79595 154547 79598
rect 154622 79525 154682 79734
rect 155125 79731 155191 79734
rect 155263 79794 155329 79797
rect 155680 79796 155740 79867
rect 155534 79794 155540 79796
rect 155263 79792 155540 79794
rect 155263 79736 155268 79792
rect 155324 79736 155540 79792
rect 155263 79734 155540 79736
rect 155263 79731 155329 79734
rect 155534 79732 155540 79734
rect 155604 79732 155610 79796
rect 155680 79734 155724 79796
rect 155718 79732 155724 79734
rect 155788 79732 155794 79796
rect 155864 79661 155924 79867
rect 154849 79660 154915 79661
rect 154798 79658 154804 79660
rect 154758 79598 154804 79658
rect 154868 79658 154915 79660
rect 155585 79658 155651 79661
rect 154868 79656 155651 79658
rect 154910 79600 155590 79656
rect 155646 79600 155651 79656
rect 154798 79596 154804 79598
rect 154868 79598 155651 79600
rect 154868 79596 154915 79598
rect 154849 79595 154915 79596
rect 155585 79595 155651 79598
rect 155861 79656 155927 79661
rect 155861 79600 155866 79656
rect 155922 79600 155927 79656
rect 155861 79595 155927 79600
rect 137970 79462 149530 79522
rect 137572 79460 137578 79462
rect 137645 79459 137711 79462
rect 130326 79324 130332 79388
rect 130396 79386 130402 79388
rect 139894 79386 139900 79388
rect 130396 79326 139900 79386
rect 130396 79324 130402 79326
rect 139894 79324 139900 79326
rect 139964 79324 139970 79388
rect 140037 79386 140103 79389
rect 140446 79386 140452 79388
rect 140037 79384 140452 79386
rect 140037 79328 140042 79384
rect 140098 79328 140452 79384
rect 140037 79326 140452 79328
rect 140037 79323 140103 79326
rect 140446 79324 140452 79326
rect 140516 79324 140522 79388
rect 140865 79386 140931 79389
rect 141325 79388 141391 79389
rect 140998 79386 141004 79388
rect 140865 79384 141004 79386
rect 140865 79328 140870 79384
rect 140926 79328 141004 79384
rect 140865 79326 141004 79328
rect 140865 79323 140931 79326
rect 140998 79324 141004 79326
rect 141068 79324 141074 79388
rect 141325 79386 141372 79388
rect 141280 79384 141372 79386
rect 141280 79328 141330 79384
rect 141280 79326 141372 79328
rect 141325 79324 141372 79326
rect 141436 79324 141442 79388
rect 141601 79386 141667 79389
rect 141734 79386 141740 79388
rect 141601 79384 141740 79386
rect 141601 79328 141606 79384
rect 141662 79328 141740 79384
rect 141601 79326 141740 79328
rect 141325 79323 141391 79324
rect 141601 79323 141667 79326
rect 141734 79324 141740 79326
rect 141804 79324 141810 79388
rect 143574 79324 143580 79388
rect 143644 79386 143650 79388
rect 144821 79386 144887 79389
rect 143644 79384 144887 79386
rect 143644 79328 144826 79384
rect 144882 79328 144887 79384
rect 143644 79326 144887 79328
rect 143644 79324 143650 79326
rect 144821 79323 144887 79326
rect 145046 79324 145052 79388
rect 145116 79386 145122 79388
rect 145281 79386 145347 79389
rect 145116 79384 145347 79386
rect 145116 79328 145286 79384
rect 145342 79328 145347 79384
rect 145116 79326 145347 79328
rect 145116 79324 145122 79326
rect 145281 79323 145347 79326
rect 145966 79324 145972 79388
rect 146036 79386 146042 79388
rect 146753 79386 146819 79389
rect 146036 79384 146819 79386
rect 146036 79328 146758 79384
rect 146814 79328 146819 79384
rect 146036 79326 146819 79328
rect 146036 79324 146042 79326
rect 146753 79323 146819 79326
rect 147070 79324 147076 79388
rect 147140 79386 147146 79388
rect 147489 79386 147555 79389
rect 148041 79388 148107 79389
rect 147140 79384 147555 79386
rect 147140 79328 147494 79384
rect 147550 79328 147555 79384
rect 147140 79326 147555 79328
rect 147140 79324 147146 79326
rect 147489 79323 147555 79326
rect 147990 79324 147996 79388
rect 148060 79386 148107 79388
rect 148060 79384 148152 79386
rect 148102 79328 148152 79384
rect 148060 79326 148152 79328
rect 148060 79324 148107 79326
rect 148542 79324 148548 79388
rect 148612 79386 148618 79388
rect 148685 79386 148751 79389
rect 149470 79386 149530 79462
rect 149646 79460 149652 79524
rect 149716 79522 149722 79524
rect 150249 79522 150315 79525
rect 150433 79522 150499 79525
rect 149716 79520 150499 79522
rect 149716 79464 150254 79520
rect 150310 79464 150438 79520
rect 150494 79464 150499 79520
rect 149716 79462 150499 79464
rect 149716 79460 149722 79462
rect 150249 79459 150315 79462
rect 150433 79459 150499 79462
rect 151353 79522 151419 79525
rect 151486 79522 151492 79524
rect 151353 79520 151492 79522
rect 151353 79464 151358 79520
rect 151414 79464 151492 79520
rect 151353 79462 151492 79464
rect 151353 79459 151419 79462
rect 151486 79460 151492 79462
rect 151556 79460 151562 79524
rect 152222 79460 152228 79524
rect 152292 79522 152298 79524
rect 153101 79522 153167 79525
rect 152292 79520 153167 79522
rect 152292 79464 153106 79520
rect 153162 79464 153167 79520
rect 152292 79462 153167 79464
rect 152292 79460 152298 79462
rect 153101 79459 153167 79462
rect 153469 79524 153535 79525
rect 153469 79520 153516 79524
rect 153580 79522 153586 79524
rect 153469 79464 153474 79520
rect 153469 79460 153516 79464
rect 153580 79462 153626 79522
rect 153580 79460 153586 79462
rect 153694 79460 153700 79524
rect 153764 79522 153770 79524
rect 153929 79522 153995 79525
rect 153764 79520 153995 79522
rect 153764 79464 153934 79520
rect 153990 79464 153995 79520
rect 153764 79462 153995 79464
rect 153764 79460 153770 79462
rect 153469 79459 153535 79460
rect 153929 79459 153995 79462
rect 154573 79520 154682 79525
rect 154573 79464 154578 79520
rect 154634 79464 154682 79520
rect 154573 79462 154682 79464
rect 156094 79522 156154 79901
rect 156454 79868 156460 79932
rect 156524 79930 156530 79932
rect 157014 79930 157074 80142
rect 157190 80004 157196 80068
rect 157260 80066 157266 80068
rect 157260 80006 158776 80066
rect 157260 80004 157266 80006
rect 157195 79930 157261 79933
rect 156524 79870 156582 79930
rect 157014 79928 157261 79930
rect 157014 79872 157200 79928
rect 157256 79872 157261 79928
rect 157014 79870 157261 79872
rect 156524 79868 156530 79870
rect 157195 79867 157261 79870
rect 157696 79868 157702 79932
rect 157766 79930 157772 79932
rect 157839 79930 157905 79933
rect 157766 79928 157905 79930
rect 157766 79872 157844 79928
rect 157900 79872 157905 79928
rect 157766 79870 157905 79872
rect 157766 79868 157772 79870
rect 157839 79867 157905 79870
rect 158110 79868 158116 79932
rect 158180 79930 158186 79932
rect 158575 79930 158641 79933
rect 158180 79928 158641 79930
rect 158180 79872 158580 79928
rect 158636 79872 158641 79928
rect 158180 79870 158641 79872
rect 158180 79868 158186 79870
rect 158575 79867 158641 79870
rect 157011 79796 157077 79797
rect 157006 79794 157012 79796
rect 156920 79734 157012 79794
rect 157006 79732 157012 79734
rect 157076 79732 157082 79796
rect 157011 79731 157077 79732
rect 156270 79596 156276 79660
rect 156340 79658 156346 79660
rect 156597 79658 156663 79661
rect 156340 79656 156663 79658
rect 156340 79600 156602 79656
rect 156658 79600 156663 79656
rect 156340 79598 156663 79600
rect 156340 79596 156346 79598
rect 156597 79595 156663 79598
rect 156505 79522 156571 79525
rect 156094 79520 156571 79522
rect 156094 79464 156510 79520
rect 156566 79464 156571 79520
rect 156094 79462 156571 79464
rect 157198 79522 157258 79867
rect 158299 79796 158365 79797
rect 158294 79794 158300 79796
rect 158164 79734 158300 79794
rect 158164 79661 158224 79734
rect 158294 79732 158300 79734
rect 158364 79732 158370 79796
rect 158716 79794 158776 80006
rect 159214 80004 159220 80068
rect 159284 80066 159290 80068
rect 161054 80066 161060 80068
rect 159284 80006 159834 80066
rect 159284 80004 159290 80006
rect 159774 79933 159834 80006
rect 160832 80006 161060 80066
rect 160832 79967 160892 80006
rect 161054 80004 161060 80006
rect 161124 80004 161130 80068
rect 160783 79962 160892 79967
rect 158846 79868 158852 79932
rect 158916 79930 158922 79932
rect 158916 79870 159466 79930
rect 158916 79868 158922 79870
rect 159406 79797 159466 79870
rect 159771 79928 159837 79933
rect 159771 79872 159776 79928
rect 159832 79872 159837 79928
rect 159771 79867 159837 79872
rect 160507 79928 160573 79933
rect 160507 79872 160512 79928
rect 160568 79872 160573 79928
rect 160783 79906 160788 79962
rect 160844 79906 160892 79962
rect 160783 79904 160892 79906
rect 161243 79962 161309 79967
rect 161243 79906 161248 79962
rect 161304 79906 161309 79962
rect 160783 79901 160849 79904
rect 161243 79901 161309 79906
rect 161611 79930 161677 79933
rect 161611 79928 161812 79930
rect 160507 79867 160573 79872
rect 160510 79797 160570 79867
rect 158624 79734 159282 79794
rect 158299 79731 158365 79732
rect 158624 79661 158684 79734
rect 157517 79658 157583 79661
rect 157517 79656 157626 79658
rect 157517 79600 157522 79656
rect 157578 79600 157626 79656
rect 157517 79595 157626 79600
rect 158161 79656 158227 79661
rect 158437 79660 158503 79661
rect 158437 79658 158484 79660
rect 158161 79600 158166 79656
rect 158222 79600 158227 79656
rect 158161 79595 158227 79600
rect 158392 79656 158484 79658
rect 158392 79600 158442 79656
rect 158392 79598 158484 79600
rect 158437 79596 158484 79598
rect 158548 79596 158554 79660
rect 158621 79656 158687 79661
rect 158621 79600 158626 79656
rect 158682 79600 158687 79656
rect 158437 79595 158503 79596
rect 158621 79595 158687 79600
rect 159222 79658 159282 79734
rect 159403 79792 159469 79797
rect 159403 79736 159408 79792
rect 159464 79736 159469 79792
rect 159403 79731 159469 79736
rect 159582 79732 159588 79796
rect 159652 79794 159658 79796
rect 159955 79794 160021 79797
rect 160185 79794 160251 79797
rect 159652 79792 160251 79794
rect 159652 79736 159960 79792
rect 160016 79736 160190 79792
rect 160246 79736 160251 79792
rect 159652 79734 160251 79736
rect 159652 79732 159658 79734
rect 159955 79731 160021 79734
rect 160185 79731 160251 79734
rect 160461 79792 160570 79797
rect 160461 79736 160466 79792
rect 160522 79736 160570 79792
rect 160461 79734 160570 79736
rect 160461 79731 160527 79734
rect 160686 79732 160692 79796
rect 160756 79794 160762 79796
rect 161059 79794 161125 79797
rect 160756 79792 161125 79794
rect 160756 79736 161064 79792
rect 161120 79736 161125 79792
rect 160756 79734 161125 79736
rect 160756 79732 160762 79734
rect 161059 79731 161125 79734
rect 160645 79658 160711 79661
rect 159222 79656 160711 79658
rect 159222 79600 160650 79656
rect 160706 79600 160711 79656
rect 159222 79598 160711 79600
rect 161246 79658 161306 79901
rect 161611 79872 161616 79928
rect 161672 79872 161812 79928
rect 161611 79870 161812 79872
rect 161611 79867 161677 79870
rect 161427 79794 161493 79797
rect 161606 79794 161612 79796
rect 161427 79792 161612 79794
rect 161427 79736 161432 79792
rect 161488 79736 161612 79792
rect 161427 79734 161612 79736
rect 161427 79731 161493 79734
rect 161606 79732 161612 79734
rect 161676 79732 161682 79796
rect 161752 79661 161812 79870
rect 161982 79797 162042 80414
rect 162710 80412 162716 80414
rect 162780 80474 162786 80476
rect 162780 80414 179430 80474
rect 162780 80412 162786 80414
rect 168284 80278 176532 80338
rect 167310 80140 167316 80204
rect 167380 80202 167386 80204
rect 167380 80142 168068 80202
rect 167380 80140 167386 80142
rect 163630 80004 163636 80068
rect 163700 80066 163706 80068
rect 163700 80004 163744 80066
rect 162715 79962 162781 79967
rect 162342 79868 162348 79932
rect 162412 79930 162418 79932
rect 162715 79930 162720 79962
rect 162412 79906 162720 79930
rect 162776 79906 162781 79962
rect 162412 79901 162781 79906
rect 163083 79928 163149 79933
rect 162412 79870 162778 79901
rect 163083 79872 163088 79928
rect 163144 79872 163149 79928
rect 162412 79868 162418 79870
rect 163083 79867 163149 79872
rect 163543 79930 163609 79933
rect 163684 79930 163744 80004
rect 166947 79962 167013 79967
rect 163543 79928 163744 79930
rect 163543 79872 163548 79928
rect 163604 79872 163744 79928
rect 163543 79870 163744 79872
rect 163543 79867 163609 79870
rect 163998 79868 164004 79932
rect 164068 79930 164074 79932
rect 164187 79930 164253 79933
rect 164068 79928 164253 79930
rect 164068 79872 164192 79928
rect 164248 79872 164253 79928
rect 164068 79870 164253 79872
rect 164068 79868 164074 79870
rect 164187 79867 164253 79870
rect 164923 79930 164989 79933
rect 165102 79930 165108 79932
rect 164923 79928 165108 79930
rect 164923 79872 164928 79928
rect 164984 79872 165108 79928
rect 164923 79870 165108 79872
rect 164923 79867 164989 79870
rect 165102 79868 165108 79870
rect 165172 79868 165178 79932
rect 165286 79868 165292 79932
rect 165356 79930 165362 79932
rect 165475 79930 165541 79933
rect 165356 79928 165541 79930
rect 165356 79872 165480 79928
rect 165536 79872 165541 79928
rect 165356 79870 165541 79872
rect 165356 79868 165362 79870
rect 165475 79867 165541 79870
rect 165843 79928 165909 79933
rect 165843 79872 165848 79928
rect 165904 79872 165909 79928
rect 165843 79867 165909 79872
rect 166022 79868 166028 79932
rect 166092 79930 166098 79932
rect 166579 79930 166645 79933
rect 166092 79928 166645 79930
rect 166092 79872 166584 79928
rect 166640 79872 166645 79928
rect 166092 79870 166645 79872
rect 166092 79868 166098 79870
rect 166579 79867 166645 79870
rect 166758 79868 166764 79932
rect 166828 79930 166834 79932
rect 166947 79930 166952 79962
rect 166828 79906 166952 79930
rect 167008 79906 167013 79962
rect 168008 79964 168068 80142
rect 168143 79964 168209 79967
rect 168008 79962 168209 79964
rect 166828 79901 167013 79906
rect 166828 79870 167010 79901
rect 166828 79868 166834 79870
rect 167494 79868 167500 79932
rect 167564 79930 167570 79932
rect 167683 79930 167749 79933
rect 167564 79928 167749 79930
rect 167564 79872 167688 79928
rect 167744 79872 167749 79928
rect 168008 79906 168148 79962
rect 168204 79906 168209 79962
rect 168008 79904 168209 79906
rect 168143 79901 168209 79904
rect 167564 79870 167749 79872
rect 167564 79868 167570 79870
rect 167683 79867 167749 79870
rect 161979 79792 162045 79797
rect 161979 79736 161984 79792
rect 162040 79736 162045 79792
rect 161979 79731 162045 79736
rect 163086 79794 163146 79867
rect 163313 79794 163379 79797
rect 163086 79792 163379 79794
rect 163086 79736 163318 79792
rect 163374 79736 163379 79792
rect 163086 79734 163379 79736
rect 163313 79731 163379 79734
rect 163446 79732 163452 79796
rect 163516 79794 163522 79796
rect 163911 79794 163977 79797
rect 164739 79796 164805 79797
rect 164734 79794 164740 79796
rect 163516 79792 163977 79794
rect 163516 79736 163916 79792
rect 163972 79736 163977 79792
rect 163516 79734 163977 79736
rect 164648 79734 164740 79794
rect 163516 79732 163522 79734
rect 163911 79731 163977 79734
rect 164734 79732 164740 79734
rect 164804 79732 164810 79796
rect 165846 79794 165906 79867
rect 166073 79794 166139 79797
rect 165846 79792 166139 79794
rect 165846 79736 166078 79792
rect 166134 79736 166139 79792
rect 165846 79734 166139 79736
rect 164739 79731 164805 79732
rect 166073 79731 166139 79734
rect 166303 79794 166369 79797
rect 166574 79794 166580 79796
rect 166303 79792 166580 79794
rect 166303 79736 166308 79792
rect 166364 79736 166580 79792
rect 166303 79734 166580 79736
rect 166303 79731 166369 79734
rect 166574 79732 166580 79734
rect 166644 79732 166650 79796
rect 168284 79794 168344 80278
rect 169702 80202 169708 80204
rect 169664 80140 169708 80202
rect 169772 80140 169778 80204
rect 170438 80202 170444 80204
rect 169848 80142 170444 80202
rect 168695 79964 168761 79967
rect 168695 79962 168804 79964
rect 168419 79932 168485 79933
rect 168414 79868 168420 79932
rect 168484 79930 168490 79932
rect 168484 79870 168576 79930
rect 168695 79906 168700 79962
rect 168756 79930 168804 79962
rect 169150 79930 169156 79932
rect 168756 79906 169156 79930
rect 168695 79901 169156 79906
rect 168744 79870 169156 79901
rect 168484 79868 168490 79870
rect 169150 79868 169156 79870
rect 169220 79868 169226 79932
rect 169431 79930 169497 79933
rect 169664 79930 169724 80140
rect 169848 79967 169908 80142
rect 170438 80140 170444 80142
rect 170508 80140 170514 80204
rect 174678 80142 175520 80202
rect 174118 80004 174124 80068
rect 174188 80066 174194 80068
rect 174188 80006 174370 80066
rect 174188 80004 174194 80006
rect 169431 79928 169724 79930
rect 169431 79872 169436 79928
rect 169492 79872 169724 79928
rect 169799 79962 169908 79967
rect 169799 79906 169804 79962
rect 169860 79906 169908 79962
rect 170075 79962 170141 79967
rect 170075 79932 170080 79962
rect 170136 79932 170141 79962
rect 172743 79962 172809 79967
rect 169799 79904 169908 79906
rect 169799 79901 169865 79904
rect 169431 79870 169724 79872
rect 168419 79867 168485 79868
rect 169431 79867 169497 79870
rect 170070 79868 170076 79932
rect 170140 79930 170146 79932
rect 170443 79930 170509 79933
rect 170806 79930 170812 79932
rect 170140 79870 170198 79930
rect 170443 79928 170812 79930
rect 170443 79872 170448 79928
rect 170504 79872 170812 79928
rect 170443 79870 170812 79872
rect 170140 79868 170146 79870
rect 170443 79867 170509 79870
rect 170806 79868 170812 79870
rect 170876 79868 170882 79932
rect 171363 79928 171429 79933
rect 171363 79872 171368 79928
rect 171424 79872 171429 79928
rect 171363 79867 171429 79872
rect 171547 79930 171613 79933
rect 171726 79930 171732 79932
rect 171547 79928 171732 79930
rect 171547 79872 171552 79928
rect 171608 79872 171732 79928
rect 171547 79870 171732 79872
rect 171547 79867 171613 79870
rect 171726 79868 171732 79870
rect 171796 79868 171802 79932
rect 172094 79868 172100 79932
rect 172164 79930 172170 79932
rect 172375 79930 172441 79933
rect 172164 79928 172441 79930
rect 172164 79872 172380 79928
rect 172436 79872 172441 79928
rect 172743 79906 172748 79962
rect 172804 79930 172809 79962
rect 173755 79962 173821 79967
rect 173382 79930 173388 79932
rect 172804 79906 173388 79930
rect 172743 79901 173388 79906
rect 172164 79870 172441 79872
rect 172746 79870 173388 79901
rect 172164 79868 172170 79870
rect 172375 79867 172441 79870
rect 173382 79868 173388 79870
rect 173452 79868 173458 79932
rect 173755 79906 173760 79962
rect 173816 79906 173821 79962
rect 173755 79901 173821 79906
rect 174310 79930 174370 80006
rect 174678 79967 174738 80142
rect 174491 79962 174557 79967
rect 174491 79930 174496 79962
rect 174310 79906 174496 79930
rect 174552 79906 174557 79962
rect 174310 79901 174557 79906
rect 174675 79962 174741 79967
rect 174675 79906 174680 79962
rect 174736 79906 174741 79962
rect 174859 79932 174925 79933
rect 174675 79901 174741 79906
rect 167134 79734 168344 79794
rect 168422 79797 168482 79867
rect 168422 79792 168531 79797
rect 169569 79796 169635 79797
rect 169518 79794 169524 79796
rect 168422 79736 168470 79792
rect 168526 79736 168531 79792
rect 168422 79734 168531 79736
rect 169478 79734 169524 79794
rect 169588 79792 169635 79796
rect 169630 79736 169635 79792
rect 161381 79658 161447 79661
rect 161246 79656 161447 79658
rect 161246 79600 161386 79656
rect 161442 79600 161447 79656
rect 161246 79598 161447 79600
rect 160645 79595 160711 79598
rect 161381 79595 161447 79598
rect 161749 79656 161815 79661
rect 161749 79600 161754 79656
rect 161810 79600 161815 79656
rect 161749 79595 161815 79600
rect 161974 79596 161980 79660
rect 162044 79658 162050 79660
rect 162209 79658 162275 79661
rect 162485 79658 162551 79661
rect 167134 79658 167194 79734
rect 168465 79731 168531 79734
rect 169518 79732 169524 79734
rect 169588 79732 169635 79736
rect 169886 79732 169892 79796
rect 169956 79794 169962 79796
rect 170121 79794 170187 79797
rect 169956 79792 170187 79794
rect 169956 79736 170126 79792
rect 170182 79736 170187 79792
rect 169956 79734 170187 79736
rect 169956 79732 169962 79734
rect 169569 79731 169635 79732
rect 170121 79731 170187 79734
rect 170254 79732 170260 79796
rect 170324 79794 170330 79796
rect 170995 79794 171061 79797
rect 170324 79792 171061 79794
rect 170324 79736 171000 79792
rect 171056 79736 171061 79792
rect 170324 79734 171061 79736
rect 170324 79732 170330 79734
rect 170995 79731 171061 79734
rect 171366 79661 171426 79867
rect 171726 79732 171732 79796
rect 171796 79794 171802 79796
rect 172007 79794 172073 79797
rect 171796 79792 172073 79794
rect 171796 79736 172012 79792
rect 172068 79736 172073 79792
rect 171796 79734 172073 79736
rect 171796 79732 171802 79734
rect 172007 79731 172073 79734
rect 172830 79732 172836 79796
rect 172900 79794 172906 79796
rect 173479 79794 173545 79797
rect 172900 79792 173545 79794
rect 172900 79736 173484 79792
rect 173540 79736 173545 79792
rect 172900 79734 173545 79736
rect 172900 79732 172906 79734
rect 173479 79731 173545 79734
rect 162044 79656 162551 79658
rect 162044 79600 162214 79656
rect 162270 79600 162490 79656
rect 162546 79600 162551 79656
rect 162044 79598 162551 79600
rect 162044 79596 162050 79598
rect 162209 79595 162275 79598
rect 162485 79595 162551 79598
rect 162902 79598 167194 79658
rect 157566 79525 157626 79595
rect 157425 79522 157491 79525
rect 157198 79520 157491 79522
rect 157198 79464 157430 79520
rect 157486 79464 157491 79520
rect 157198 79462 157491 79464
rect 157566 79520 157675 79525
rect 157566 79464 157614 79520
rect 157670 79464 157675 79520
rect 157566 79462 157675 79464
rect 154573 79459 154639 79462
rect 156505 79459 156571 79462
rect 157425 79459 157491 79462
rect 157609 79459 157675 79462
rect 157977 79520 158043 79525
rect 157977 79464 157982 79520
rect 158038 79464 158043 79520
rect 157977 79459 158043 79464
rect 158110 79460 158116 79524
rect 158180 79522 158186 79524
rect 158713 79522 158779 79525
rect 158180 79520 158779 79522
rect 158180 79464 158718 79520
rect 158774 79464 158779 79520
rect 158180 79462 158779 79464
rect 158180 79460 158186 79462
rect 158713 79459 158779 79462
rect 159030 79460 159036 79524
rect 159100 79522 159106 79524
rect 159817 79522 159883 79525
rect 159100 79520 159883 79522
rect 159100 79464 159822 79520
rect 159878 79464 159883 79520
rect 159100 79462 159883 79464
rect 159100 79460 159106 79462
rect 159817 79459 159883 79462
rect 160502 79460 160508 79524
rect 160572 79522 160578 79524
rect 160737 79522 160803 79525
rect 161105 79524 161171 79525
rect 161054 79522 161060 79524
rect 160572 79520 160803 79522
rect 160572 79464 160742 79520
rect 160798 79464 160803 79520
rect 160572 79462 160803 79464
rect 161014 79462 161060 79522
rect 161124 79520 161171 79524
rect 161166 79464 161171 79520
rect 160572 79460 160578 79462
rect 160737 79459 160803 79462
rect 161054 79460 161060 79462
rect 161124 79460 161171 79464
rect 161105 79459 161171 79460
rect 162393 79522 162459 79525
rect 162902 79522 162962 79598
rect 167494 79596 167500 79660
rect 167564 79658 167570 79660
rect 167729 79658 167795 79661
rect 167564 79656 167795 79658
rect 167564 79600 167734 79656
rect 167790 79600 167795 79656
rect 167564 79598 167795 79600
rect 167564 79596 167570 79598
rect 167729 79595 167795 79598
rect 167862 79596 167868 79660
rect 167932 79658 167938 79660
rect 168189 79658 168255 79661
rect 167932 79656 168255 79658
rect 167932 79600 168194 79656
rect 168250 79600 168255 79656
rect 167932 79598 168255 79600
rect 167932 79596 167938 79598
rect 168189 79595 168255 79598
rect 168782 79596 168788 79660
rect 168852 79658 168858 79660
rect 169017 79658 169083 79661
rect 169385 79660 169451 79661
rect 168852 79656 169083 79658
rect 168852 79600 169022 79656
rect 169078 79600 169083 79656
rect 168852 79598 169083 79600
rect 168852 79596 168858 79598
rect 169017 79595 169083 79598
rect 169334 79596 169340 79660
rect 169404 79658 169451 79660
rect 169661 79658 169727 79661
rect 169404 79656 169727 79658
rect 169446 79600 169666 79656
rect 169722 79600 169727 79656
rect 169404 79598 169727 79600
rect 169404 79596 169451 79598
rect 169385 79595 169451 79596
rect 169661 79595 169727 79598
rect 170397 79658 170463 79661
rect 170622 79658 170628 79660
rect 170397 79656 170628 79658
rect 170397 79600 170402 79656
rect 170458 79600 170628 79656
rect 170397 79598 170628 79600
rect 170397 79595 170463 79598
rect 170622 79596 170628 79598
rect 170692 79596 170698 79660
rect 171317 79656 171426 79661
rect 171317 79600 171322 79656
rect 171378 79600 171426 79656
rect 171317 79598 171426 79600
rect 171777 79658 171843 79661
rect 172605 79660 172671 79661
rect 171910 79658 171916 79660
rect 171777 79656 171916 79658
rect 171777 79600 171782 79656
rect 171838 79600 171916 79656
rect 171777 79598 171916 79600
rect 171317 79595 171383 79598
rect 171777 79595 171843 79598
rect 171910 79596 171916 79598
rect 171980 79596 171986 79660
rect 172605 79658 172652 79660
rect 172524 79656 172652 79658
rect 172716 79658 172722 79660
rect 173758 79658 173818 79901
rect 174123 79894 174189 79899
rect 174123 79838 174128 79894
rect 174184 79838 174189 79894
rect 174310 79870 174554 79901
rect 174854 79868 174860 79932
rect 174924 79930 174930 79932
rect 175135 79930 175201 79933
rect 174924 79870 175016 79930
rect 175092 79928 175201 79930
rect 175092 79872 175140 79928
rect 175196 79872 175201 79928
rect 174924 79868 174930 79870
rect 174859 79867 174925 79868
rect 175092 79867 175201 79872
rect 174123 79833 174189 79838
rect 174126 79661 174186 79833
rect 175092 79797 175152 79867
rect 174302 79732 174308 79796
rect 174372 79794 174378 79796
rect 175089 79794 175155 79797
rect 174372 79792 175155 79794
rect 174372 79736 175094 79792
rect 175150 79736 175155 79792
rect 174372 79734 175155 79736
rect 175460 79794 175520 80142
rect 176472 80066 176532 80278
rect 177246 80276 177252 80340
rect 177316 80338 177322 80340
rect 178493 80338 178559 80341
rect 177316 80336 178559 80338
rect 177316 80280 178498 80336
rect 178554 80280 178559 80336
rect 177316 80278 178559 80280
rect 177316 80276 177322 80278
rect 178493 80275 178559 80278
rect 179370 80202 179430 80414
rect 184974 80276 184980 80340
rect 185044 80338 185050 80340
rect 185209 80338 185275 80341
rect 185044 80336 185275 80338
rect 185044 80280 185214 80336
rect 185270 80280 185275 80336
rect 185044 80278 185275 80280
rect 185044 80276 185050 80278
rect 185209 80275 185275 80278
rect 382273 80202 382339 80205
rect 179370 80200 382339 80202
rect 179370 80144 382278 80200
rect 382334 80144 382339 80200
rect 179370 80142 382339 80144
rect 382273 80139 382339 80142
rect 176472 80006 183570 80066
rect 175963 79962 176029 79967
rect 175590 79868 175596 79932
rect 175660 79930 175666 79932
rect 175963 79930 175968 79962
rect 175660 79906 175968 79930
rect 176024 79906 176029 79962
rect 175660 79901 176029 79906
rect 176147 79928 176213 79933
rect 176694 79930 176700 79932
rect 175660 79870 176026 79901
rect 176147 79872 176152 79928
rect 176208 79872 176213 79928
rect 175660 79868 175666 79870
rect 176147 79867 176213 79872
rect 176656 79868 176700 79930
rect 176764 79930 176770 79932
rect 177343 79930 177409 79933
rect 177573 79932 177639 79933
rect 177573 79930 177620 79932
rect 176764 79928 177409 79930
rect 176764 79872 177348 79928
rect 177404 79872 177409 79928
rect 176764 79870 177409 79872
rect 177528 79928 177620 79930
rect 177528 79872 177578 79928
rect 177528 79870 177620 79872
rect 176764 79868 176770 79870
rect 176150 79797 176210 79867
rect 176009 79796 176075 79797
rect 175590 79794 175596 79796
rect 175460 79734 175596 79794
rect 174372 79732 174378 79734
rect 175089 79731 175155 79734
rect 175590 79732 175596 79734
rect 175660 79732 175666 79796
rect 175958 79794 175964 79796
rect 175918 79734 175964 79794
rect 176028 79792 176075 79796
rect 176070 79736 176075 79792
rect 175958 79732 175964 79734
rect 176028 79732 176075 79736
rect 176150 79792 176259 79797
rect 176331 79796 176397 79797
rect 176150 79736 176198 79792
rect 176254 79736 176259 79792
rect 176150 79734 176259 79736
rect 176009 79731 176075 79732
rect 176193 79731 176259 79734
rect 176326 79732 176332 79796
rect 176396 79794 176402 79796
rect 176396 79734 176488 79794
rect 176396 79732 176402 79734
rect 176331 79731 176397 79732
rect 176656 79661 176716 79868
rect 177343 79867 177409 79870
rect 177573 79868 177620 79870
rect 177684 79868 177690 79932
rect 177573 79867 177639 79868
rect 176878 79732 176884 79796
rect 176948 79794 176954 79796
rect 177481 79794 177547 79797
rect 177849 79794 177915 79797
rect 176948 79792 177915 79794
rect 176948 79736 177486 79792
rect 177542 79736 177854 79792
rect 177910 79736 177915 79792
rect 176948 79734 177915 79736
rect 183510 79794 183570 80006
rect 196566 80004 196572 80068
rect 196636 80066 196642 80068
rect 196801 80066 196867 80069
rect 196636 80064 196867 80066
rect 196636 80008 196806 80064
rect 196862 80008 196867 80064
rect 196636 80006 196867 80008
rect 196636 80004 196642 80006
rect 196801 80003 196867 80006
rect 306373 79794 306439 79797
rect 183510 79792 306439 79794
rect 183510 79736 306378 79792
rect 306434 79736 306439 79792
rect 183510 79734 306439 79736
rect 176948 79732 176954 79734
rect 177481 79731 177547 79734
rect 177849 79731 177915 79734
rect 306373 79731 306439 79734
rect 172524 79600 172610 79656
rect 172524 79598 172652 79600
rect 172605 79596 172652 79598
rect 172716 79598 173818 79658
rect 174077 79656 174186 79661
rect 174077 79600 174082 79656
rect 174138 79600 174186 79656
rect 174077 79598 174186 79600
rect 174353 79658 174419 79661
rect 174486 79658 174492 79660
rect 174353 79656 174492 79658
rect 174353 79600 174358 79656
rect 174414 79600 174492 79656
rect 174353 79598 174492 79600
rect 172716 79596 172722 79598
rect 172605 79595 172671 79596
rect 174077 79595 174143 79598
rect 174353 79595 174419 79598
rect 174486 79596 174492 79598
rect 174556 79596 174562 79660
rect 174905 79658 174971 79661
rect 175038 79658 175044 79660
rect 174905 79656 175044 79658
rect 174905 79600 174910 79656
rect 174966 79600 175044 79656
rect 174905 79598 175044 79600
rect 174905 79595 174971 79598
rect 175038 79596 175044 79598
rect 175108 79596 175114 79660
rect 175222 79596 175228 79660
rect 175292 79658 175298 79660
rect 176101 79658 176167 79661
rect 175292 79656 176167 79658
rect 175292 79600 176106 79656
rect 176162 79600 176167 79656
rect 175292 79598 176167 79600
rect 175292 79596 175298 79598
rect 176101 79595 176167 79598
rect 176377 79658 176443 79661
rect 176510 79658 176516 79660
rect 176377 79656 176516 79658
rect 176377 79600 176382 79656
rect 176438 79600 176516 79656
rect 176377 79598 176516 79600
rect 176377 79595 176443 79598
rect 176510 79596 176516 79598
rect 176580 79596 176586 79660
rect 176653 79656 176719 79661
rect 176653 79600 176658 79656
rect 176714 79600 176719 79656
rect 176653 79595 176719 79600
rect 162393 79520 162962 79522
rect 162393 79464 162398 79520
rect 162454 79464 162962 79520
rect 162393 79462 162962 79464
rect 162393 79459 162459 79462
rect 163262 79460 163268 79524
rect 163332 79522 163338 79524
rect 163497 79522 163563 79525
rect 164049 79522 164115 79525
rect 178677 79522 178743 79525
rect 163332 79520 163563 79522
rect 163332 79464 163502 79520
rect 163558 79464 163563 79520
rect 163332 79462 163563 79464
rect 163332 79460 163338 79462
rect 163497 79459 163563 79462
rect 163638 79520 178743 79522
rect 163638 79464 164054 79520
rect 164110 79464 178682 79520
rect 178738 79464 178743 79520
rect 163638 79462 178743 79464
rect 151077 79386 151143 79389
rect 155585 79388 155651 79389
rect 155534 79386 155540 79388
rect 148612 79384 149346 79386
rect 148612 79328 148690 79384
rect 148746 79328 149346 79384
rect 148612 79326 149346 79328
rect 149470 79384 151143 79386
rect 149470 79328 151082 79384
rect 151138 79328 151143 79384
rect 149470 79326 151143 79328
rect 155494 79326 155540 79386
rect 155604 79384 155651 79388
rect 155646 79328 155651 79384
rect 148612 79324 148618 79326
rect 148041 79323 148107 79324
rect 148685 79323 148751 79326
rect 125358 79188 125364 79252
rect 125428 79250 125434 79252
rect 146201 79250 146267 79253
rect 125428 79248 146267 79250
rect 125428 79192 146206 79248
rect 146262 79192 146267 79248
rect 125428 79190 146267 79192
rect 125428 79188 125434 79190
rect 146201 79187 146267 79190
rect 147070 79188 147076 79252
rect 147140 79250 147146 79252
rect 147213 79250 147279 79253
rect 147140 79248 147279 79250
rect 147140 79192 147218 79248
rect 147274 79192 147279 79248
rect 147140 79190 147279 79192
rect 147140 79188 147146 79190
rect 147213 79187 147279 79190
rect 147397 79250 147463 79253
rect 148685 79252 148751 79253
rect 148174 79250 148180 79252
rect 147397 79248 148180 79250
rect 147397 79192 147402 79248
rect 147458 79192 148180 79248
rect 147397 79190 148180 79192
rect 147397 79187 147463 79190
rect 148174 79188 148180 79190
rect 148244 79250 148250 79252
rect 148542 79250 148548 79252
rect 148244 79190 148548 79250
rect 148244 79188 148250 79190
rect 148542 79188 148548 79190
rect 148612 79188 148618 79252
rect 148685 79248 148732 79252
rect 148796 79250 148802 79252
rect 148961 79250 149027 79253
rect 149094 79250 149100 79252
rect 148685 79192 148690 79248
rect 148685 79188 148732 79192
rect 148796 79190 148842 79250
rect 148961 79248 149100 79250
rect 148961 79192 148966 79248
rect 149022 79192 149100 79248
rect 148961 79190 149100 79192
rect 148796 79188 148802 79190
rect 148685 79187 148751 79188
rect 148961 79187 149027 79190
rect 149094 79188 149100 79190
rect 149164 79188 149170 79252
rect 149286 79250 149346 79326
rect 151077 79323 151143 79326
rect 155534 79324 155540 79326
rect 155604 79324 155651 79328
rect 155585 79323 155651 79324
rect 149421 79250 149487 79253
rect 149286 79248 149487 79250
rect 149286 79192 149426 79248
rect 149482 79192 149487 79248
rect 149286 79190 149487 79192
rect 149421 79187 149487 79190
rect 149830 79188 149836 79252
rect 149900 79250 149906 79252
rect 150341 79250 150407 79253
rect 149900 79248 150407 79250
rect 149900 79192 150346 79248
rect 150402 79192 150407 79248
rect 149900 79190 150407 79192
rect 149900 79188 149906 79190
rect 150341 79187 150407 79190
rect 154614 79188 154620 79252
rect 154684 79250 154690 79252
rect 154757 79250 154823 79253
rect 155769 79250 155835 79253
rect 154684 79248 155835 79250
rect 154684 79192 154762 79248
rect 154818 79192 155774 79248
rect 155830 79192 155835 79248
rect 154684 79190 155835 79192
rect 154684 79188 154690 79190
rect 154757 79187 154823 79190
rect 155769 79187 155835 79190
rect 156965 79252 157031 79253
rect 156965 79248 157012 79252
rect 157076 79250 157082 79252
rect 157980 79250 158040 79459
rect 158161 79386 158227 79389
rect 158294 79386 158300 79388
rect 158161 79384 158300 79386
rect 158161 79328 158166 79384
rect 158222 79328 158300 79384
rect 158161 79326 158300 79328
rect 158161 79323 158227 79326
rect 158294 79324 158300 79326
rect 158364 79324 158370 79388
rect 162158 79324 162164 79388
rect 162228 79386 162234 79388
rect 162577 79386 162643 79389
rect 162228 79384 162643 79386
rect 162228 79328 162582 79384
rect 162638 79328 162643 79384
rect 162228 79326 162643 79328
rect 162228 79324 162234 79326
rect 162577 79323 162643 79326
rect 162894 79324 162900 79388
rect 162964 79386 162970 79388
rect 163638 79386 163698 79462
rect 164049 79459 164115 79462
rect 178677 79459 178743 79462
rect 164601 79388 164667 79389
rect 164550 79386 164556 79388
rect 162964 79326 163698 79386
rect 164510 79326 164556 79386
rect 164620 79384 164667 79388
rect 164662 79328 164667 79384
rect 162964 79324 162970 79326
rect 164550 79324 164556 79326
rect 164620 79324 164667 79328
rect 165838 79324 165844 79388
rect 165908 79386 165914 79388
rect 167177 79386 167243 79389
rect 165908 79384 167243 79386
rect 165908 79328 167182 79384
rect 167238 79328 167243 79384
rect 165908 79326 167243 79328
rect 165908 79324 165914 79326
rect 164601 79323 164667 79324
rect 167177 79323 167243 79326
rect 167453 79386 167519 79389
rect 168046 79386 168052 79388
rect 167453 79384 168052 79386
rect 167453 79328 167458 79384
rect 167514 79328 168052 79384
rect 167453 79326 168052 79328
rect 167453 79323 167519 79326
rect 168046 79324 168052 79326
rect 168116 79386 168122 79388
rect 168189 79386 168255 79389
rect 168116 79384 168255 79386
rect 168116 79328 168194 79384
rect 168250 79328 168255 79384
rect 168116 79326 168255 79328
rect 168116 79324 168122 79326
rect 168189 79323 168255 79326
rect 168966 79324 168972 79388
rect 169036 79386 169042 79388
rect 169385 79386 169451 79389
rect 169036 79384 169451 79386
rect 169036 79328 169390 79384
rect 169446 79328 169451 79384
rect 169036 79326 169451 79328
rect 169036 79324 169042 79326
rect 169385 79323 169451 79326
rect 170581 79386 170647 79389
rect 171358 79386 171364 79388
rect 170581 79384 171364 79386
rect 170581 79328 170586 79384
rect 170642 79328 171364 79384
rect 170581 79326 171364 79328
rect 170581 79323 170647 79326
rect 171358 79324 171364 79326
rect 171428 79324 171434 79388
rect 171542 79324 171548 79388
rect 171612 79386 171618 79388
rect 172237 79386 172303 79389
rect 171612 79384 172303 79386
rect 171612 79328 172242 79384
rect 172298 79328 172303 79384
rect 171612 79326 172303 79328
rect 171612 79324 171618 79326
rect 172237 79323 172303 79326
rect 172973 79388 173039 79389
rect 173249 79388 173315 79389
rect 172973 79384 173020 79388
rect 173084 79386 173090 79388
rect 172973 79328 172978 79384
rect 172973 79324 173020 79328
rect 173084 79326 173130 79386
rect 173084 79324 173090 79326
rect 173198 79324 173204 79388
rect 173268 79386 173315 79388
rect 173268 79384 173360 79386
rect 173310 79328 173360 79384
rect 173268 79326 173360 79328
rect 173268 79324 173315 79326
rect 173566 79324 173572 79388
rect 173636 79386 173642 79388
rect 173893 79386 173959 79389
rect 173636 79384 173959 79386
rect 173636 79328 173898 79384
rect 173954 79328 173959 79384
rect 173636 79326 173959 79328
rect 173636 79324 173642 79326
rect 172973 79323 173039 79324
rect 173249 79323 173315 79324
rect 173893 79323 173959 79326
rect 174537 79386 174603 79389
rect 174670 79386 174676 79388
rect 174537 79384 174676 79386
rect 174537 79328 174542 79384
rect 174598 79328 174676 79384
rect 174537 79326 174676 79328
rect 174537 79323 174603 79326
rect 174670 79324 174676 79326
rect 174740 79324 174746 79388
rect 175406 79324 175412 79388
rect 175476 79386 175482 79388
rect 175641 79386 175707 79389
rect 175476 79384 175707 79386
rect 175476 79328 175646 79384
rect 175702 79328 175707 79384
rect 175476 79326 175707 79328
rect 175476 79324 175482 79326
rect 175641 79323 175707 79326
rect 175774 79324 175780 79388
rect 175844 79386 175850 79388
rect 175917 79386 175983 79389
rect 187182 79386 187188 79388
rect 175844 79384 175983 79386
rect 175844 79328 175922 79384
rect 175978 79328 175983 79384
rect 175844 79326 175983 79328
rect 175844 79324 175850 79326
rect 175917 79323 175983 79326
rect 176150 79326 187188 79386
rect 158294 79250 158300 79252
rect 156965 79192 156970 79248
rect 156965 79188 157012 79192
rect 157076 79190 157122 79250
rect 157980 79190 158300 79250
rect 157076 79188 157082 79190
rect 158294 79188 158300 79190
rect 158364 79188 158370 79252
rect 164918 79188 164924 79252
rect 164988 79250 164994 79252
rect 165153 79250 165219 79253
rect 164988 79248 165219 79250
rect 164988 79192 165158 79248
rect 165214 79192 165219 79248
rect 164988 79190 165219 79192
rect 164988 79188 164994 79190
rect 156965 79187 157031 79188
rect 165153 79187 165219 79190
rect 166206 79188 166212 79252
rect 166276 79250 166282 79252
rect 166533 79250 166599 79253
rect 166276 79248 166599 79250
rect 166276 79192 166538 79248
rect 166594 79192 166599 79248
rect 166276 79190 166599 79192
rect 166276 79188 166282 79190
rect 166533 79187 166599 79190
rect 167678 79188 167684 79252
rect 167748 79250 167754 79252
rect 168281 79250 168347 79253
rect 167748 79248 168347 79250
rect 167748 79192 168286 79248
rect 168342 79192 168347 79248
rect 167748 79190 168347 79192
rect 167748 79188 167754 79190
rect 168281 79187 168347 79190
rect 169937 79250 170003 79253
rect 170949 79252 171015 79253
rect 171961 79252 172027 79253
rect 170806 79250 170812 79252
rect 169937 79248 170812 79250
rect 169937 79192 169942 79248
rect 169998 79192 170812 79248
rect 169937 79190 170812 79192
rect 169937 79187 170003 79190
rect 170806 79188 170812 79190
rect 170876 79188 170882 79252
rect 170949 79248 170996 79252
rect 171060 79250 171066 79252
rect 171910 79250 171916 79252
rect 170949 79192 170954 79248
rect 170949 79188 170996 79192
rect 171060 79190 171106 79250
rect 171870 79190 171916 79250
rect 171980 79248 172027 79252
rect 172022 79192 172027 79248
rect 171060 79188 171066 79190
rect 171910 79188 171916 79190
rect 171980 79188 172027 79192
rect 170949 79187 171015 79188
rect 171961 79187 172027 79188
rect 175181 79250 175247 79253
rect 176150 79250 176210 79326
rect 187182 79324 187188 79326
rect 187252 79324 187258 79388
rect 191598 79324 191604 79388
rect 191668 79386 191674 79388
rect 580257 79386 580323 79389
rect 191668 79384 580323 79386
rect 191668 79328 580262 79384
rect 580318 79328 580323 79384
rect 191668 79326 580323 79328
rect 191668 79324 191674 79326
rect 580257 79323 580323 79326
rect 175181 79248 176210 79250
rect 175181 79192 175186 79248
rect 175242 79192 176210 79248
rect 175181 79190 176210 79192
rect 176745 79250 176811 79253
rect 177062 79250 177068 79252
rect 176745 79248 177068 79250
rect 176745 79192 176750 79248
rect 176806 79192 177068 79248
rect 176745 79190 177068 79192
rect 175181 79187 175247 79190
rect 176745 79187 176811 79190
rect 177062 79188 177068 79190
rect 177132 79188 177138 79252
rect 177297 79250 177363 79253
rect 178033 79250 178099 79253
rect 187734 79250 187740 79252
rect 177297 79248 187740 79250
rect 177297 79192 177302 79248
rect 177358 79192 178038 79248
rect 178094 79192 187740 79248
rect 177297 79190 187740 79192
rect 177297 79187 177363 79190
rect 178033 79187 178099 79190
rect 187734 79188 187740 79190
rect 187804 79188 187810 79252
rect 119470 79052 119476 79116
rect 119540 79114 119546 79116
rect 151905 79114 151971 79117
rect 153009 79114 153075 79117
rect 119540 79112 153075 79114
rect 119540 79056 151910 79112
rect 151966 79056 153014 79112
rect 153070 79056 153075 79112
rect 119540 79054 153075 79056
rect 119540 79052 119546 79054
rect 151905 79051 151971 79054
rect 153009 79051 153075 79054
rect 156413 79114 156479 79117
rect 156638 79114 156644 79116
rect 156413 79112 156644 79114
rect 156413 79056 156418 79112
rect 156474 79056 156644 79112
rect 156413 79054 156644 79056
rect 156413 79051 156479 79054
rect 156638 79052 156644 79054
rect 156708 79114 156714 79116
rect 156965 79114 157031 79117
rect 156708 79112 157031 79114
rect 156708 79056 156970 79112
rect 157026 79056 157031 79112
rect 156708 79054 157031 79056
rect 156708 79052 156714 79054
rect 156965 79051 157031 79054
rect 157885 79114 157951 79117
rect 159398 79114 159404 79116
rect 157885 79112 159404 79114
rect 157885 79056 157890 79112
rect 157946 79056 159404 79112
rect 157885 79054 159404 79056
rect 157885 79051 157951 79054
rect 159398 79052 159404 79054
rect 159468 79052 159474 79116
rect 161238 79052 161244 79116
rect 161308 79114 161314 79116
rect 169753 79114 169819 79117
rect 161308 79112 169819 79114
rect 161308 79056 169758 79112
rect 169814 79056 169819 79112
rect 161308 79054 169819 79056
rect 161308 79052 161314 79054
rect 169753 79051 169819 79054
rect 171685 79114 171751 79117
rect 191966 79114 191972 79116
rect 171685 79112 191972 79114
rect 171685 79056 171690 79112
rect 171746 79056 191972 79112
rect 171685 79054 191972 79056
rect 171685 79051 171751 79054
rect 191966 79052 191972 79054
rect 192036 79052 192042 79116
rect 122598 78916 122604 78980
rect 122668 78978 122674 78980
rect 156137 78978 156203 78981
rect 158069 78978 158135 78981
rect 122668 78976 158135 78978
rect 122668 78920 156142 78976
rect 156198 78920 158074 78976
rect 158130 78920 158135 78976
rect 122668 78918 158135 78920
rect 122668 78916 122674 78918
rect 156137 78915 156203 78918
rect 158069 78915 158135 78918
rect 158662 78916 158668 78980
rect 158732 78978 158738 78980
rect 158897 78978 158963 78981
rect 158732 78976 158963 78978
rect 158732 78920 158902 78976
rect 158958 78920 158963 78976
rect 158732 78918 158963 78920
rect 158732 78916 158738 78918
rect 158897 78915 158963 78918
rect 163129 78978 163195 78981
rect 163814 78978 163820 78980
rect 163129 78976 163820 78978
rect 163129 78920 163134 78976
rect 163190 78920 163820 78976
rect 163129 78918 163820 78920
rect 163129 78915 163195 78918
rect 163814 78916 163820 78918
rect 163884 78916 163890 78980
rect 170489 78978 170555 78981
rect 190678 78978 190684 78980
rect 170489 78976 190684 78978
rect 170489 78920 170494 78976
rect 170550 78920 190684 78976
rect 170489 78918 190684 78920
rect 170489 78915 170555 78918
rect 190678 78916 190684 78918
rect 190748 78916 190754 78980
rect 122414 78780 122420 78844
rect 122484 78842 122490 78844
rect 156873 78842 156939 78845
rect 122484 78840 156939 78842
rect 122484 78784 156878 78840
rect 156934 78784 156939 78840
rect 122484 78782 156939 78784
rect 122484 78780 122490 78782
rect 156873 78779 156939 78782
rect 157701 78842 157767 78845
rect 157926 78842 157932 78844
rect 157701 78840 157932 78842
rect 157701 78784 157706 78840
rect 157762 78784 157932 78840
rect 157701 78782 157932 78784
rect 157701 78779 157767 78782
rect 157926 78780 157932 78782
rect 157996 78780 158002 78844
rect 165245 78842 165311 78845
rect 166625 78844 166691 78845
rect 165470 78842 165476 78844
rect 165245 78840 165476 78842
rect 165245 78784 165250 78840
rect 165306 78784 165476 78840
rect 165245 78782 165476 78784
rect 165245 78779 165311 78782
rect 165470 78780 165476 78782
rect 165540 78780 165546 78844
rect 166574 78842 166580 78844
rect 166534 78782 166580 78842
rect 166644 78840 166691 78844
rect 166686 78784 166691 78840
rect 166574 78780 166580 78782
rect 166644 78780 166691 78784
rect 166625 78779 166691 78780
rect 171317 78842 171383 78845
rect 176193 78842 176259 78845
rect 206277 78842 206343 78845
rect 171317 78840 174554 78842
rect 171317 78784 171322 78840
rect 171378 78784 174554 78840
rect 171317 78782 174554 78784
rect 171317 78779 171383 78782
rect 126462 78644 126468 78708
rect 126532 78706 126538 78708
rect 131021 78706 131087 78709
rect 126532 78704 131087 78706
rect 126532 78648 131026 78704
rect 131082 78648 131087 78704
rect 126532 78646 131087 78648
rect 126532 78644 126538 78646
rect 131021 78643 131087 78646
rect 132217 78706 132283 78709
rect 143533 78706 143599 78709
rect 132217 78704 143599 78706
rect 132217 78648 132222 78704
rect 132278 78648 143538 78704
rect 143594 78648 143599 78704
rect 132217 78646 143599 78648
rect 132217 78643 132283 78646
rect 143533 78643 143599 78646
rect 146702 78644 146708 78708
rect 146772 78706 146778 78708
rect 147305 78706 147371 78709
rect 146772 78704 147371 78706
rect 146772 78648 147310 78704
rect 147366 78648 147371 78704
rect 146772 78646 147371 78648
rect 146772 78644 146778 78646
rect 120022 78508 120028 78572
rect 120092 78570 120098 78572
rect 121310 78570 121316 78572
rect 120092 78510 121316 78570
rect 120092 78508 120098 78510
rect 121310 78508 121316 78510
rect 121380 78570 121386 78572
rect 132033 78570 132099 78573
rect 121380 78568 132099 78570
rect 121380 78512 132038 78568
rect 132094 78512 132099 78568
rect 121380 78510 132099 78512
rect 121380 78508 121386 78510
rect 132033 78507 132099 78510
rect 133965 78570 134031 78573
rect 134742 78570 134748 78572
rect 133965 78568 134748 78570
rect 133965 78512 133970 78568
rect 134026 78512 134748 78568
rect 133965 78510 134748 78512
rect 133965 78507 134031 78510
rect 134742 78508 134748 78510
rect 134812 78508 134818 78572
rect 135662 78508 135668 78572
rect 135732 78570 135738 78572
rect 135989 78570 136055 78573
rect 139894 78570 139900 78572
rect 135732 78568 136055 78570
rect 135732 78512 135994 78568
rect 136050 78512 136055 78568
rect 135732 78510 136055 78512
rect 135732 78508 135738 78510
rect 135989 78507 136055 78510
rect 138062 78510 139900 78570
rect 124029 78436 124095 78437
rect 124029 78434 124076 78436
rect 123984 78432 124076 78434
rect 123984 78376 124034 78432
rect 123984 78374 124076 78376
rect 124029 78372 124076 78374
rect 124140 78372 124146 78436
rect 124990 78372 124996 78436
rect 125060 78434 125066 78436
rect 138062 78434 138122 78510
rect 139894 78508 139900 78510
rect 139964 78508 139970 78572
rect 140773 78570 140839 78573
rect 141918 78570 141924 78572
rect 140773 78568 141924 78570
rect 140773 78512 140778 78568
rect 140834 78512 141924 78568
rect 140773 78510 141924 78512
rect 140773 78507 140839 78510
rect 141918 78508 141924 78510
rect 141988 78508 141994 78572
rect 144126 78508 144132 78572
rect 144196 78570 144202 78572
rect 144545 78570 144611 78573
rect 146385 78572 146451 78573
rect 144196 78568 144611 78570
rect 144196 78512 144550 78568
rect 144606 78512 144611 78568
rect 144196 78510 144611 78512
rect 144196 78508 144202 78510
rect 144545 78507 144611 78510
rect 146334 78508 146340 78572
rect 146404 78570 146451 78572
rect 146404 78568 146496 78570
rect 146446 78512 146496 78568
rect 146404 78510 146496 78512
rect 146404 78508 146451 78510
rect 146385 78507 146451 78508
rect 125060 78374 138122 78434
rect 138657 78434 138723 78437
rect 138790 78434 138796 78436
rect 138657 78432 138796 78434
rect 138657 78376 138662 78432
rect 138718 78376 138796 78432
rect 138657 78374 138796 78376
rect 125060 78372 125066 78374
rect 124029 78371 124095 78372
rect 138657 78371 138723 78374
rect 138790 78372 138796 78374
rect 138860 78372 138866 78436
rect 146710 78434 146770 78644
rect 147305 78643 147371 78646
rect 147806 78644 147812 78708
rect 147876 78706 147882 78708
rect 147876 78646 151922 78706
rect 147876 78644 147882 78646
rect 151445 78572 151511 78573
rect 149094 78508 149100 78572
rect 149164 78570 149170 78572
rect 150198 78570 150204 78572
rect 149164 78510 150204 78570
rect 149164 78508 149170 78510
rect 150198 78508 150204 78510
rect 150268 78508 150274 78572
rect 151445 78568 151492 78572
rect 151556 78570 151562 78572
rect 151445 78512 151450 78568
rect 151445 78508 151492 78512
rect 151556 78510 151602 78570
rect 151556 78508 151562 78510
rect 151445 78507 151511 78508
rect 150525 78434 150591 78437
rect 140730 78374 146770 78434
rect 147630 78432 150591 78434
rect 147630 78376 150530 78432
rect 150586 78376 150591 78432
rect 147630 78374 150591 78376
rect 151862 78434 151922 78646
rect 154062 78644 154068 78708
rect 154132 78706 154138 78708
rect 154205 78706 154271 78709
rect 154132 78704 154271 78706
rect 154132 78648 154210 78704
rect 154266 78648 154271 78704
rect 154132 78646 154271 78648
rect 154132 78644 154138 78646
rect 154205 78643 154271 78646
rect 159950 78644 159956 78708
rect 160020 78706 160026 78708
rect 171501 78706 171567 78709
rect 160020 78704 171567 78706
rect 160020 78648 171506 78704
rect 171562 78648 171567 78704
rect 160020 78646 171567 78648
rect 160020 78644 160026 78646
rect 171501 78643 171567 78646
rect 171726 78644 171732 78708
rect 171796 78706 171802 78708
rect 171961 78706 172027 78709
rect 171796 78704 172027 78706
rect 171796 78648 171966 78704
rect 172022 78648 172027 78704
rect 171796 78646 172027 78648
rect 171796 78644 171802 78646
rect 171961 78643 172027 78646
rect 172094 78644 172100 78708
rect 172164 78706 172170 78708
rect 174353 78706 174419 78709
rect 172164 78704 174419 78706
rect 172164 78648 174358 78704
rect 174414 78648 174419 78704
rect 172164 78646 174419 78648
rect 174494 78706 174554 78782
rect 176193 78840 206343 78842
rect 176193 78784 176198 78840
rect 176254 78784 206282 78840
rect 206338 78784 206343 78840
rect 176193 78782 206343 78784
rect 176193 78779 176259 78782
rect 206277 78779 206343 78782
rect 178217 78706 178283 78709
rect 174494 78704 178283 78706
rect 174494 78648 178222 78704
rect 178278 78648 178283 78704
rect 174494 78646 178283 78648
rect 172164 78644 172170 78646
rect 174353 78643 174419 78646
rect 178217 78643 178283 78646
rect 178350 78644 178356 78708
rect 178420 78706 178426 78708
rect 178861 78706 178927 78709
rect 178420 78704 178927 78706
rect 178420 78648 178866 78704
rect 178922 78648 178927 78704
rect 178420 78646 178927 78648
rect 178420 78644 178426 78646
rect 178861 78643 178927 78646
rect 158529 78570 158595 78573
rect 161197 78572 161263 78573
rect 163773 78572 163839 78573
rect 158662 78570 158668 78572
rect 158529 78568 158668 78570
rect 158529 78512 158534 78568
rect 158590 78512 158668 78568
rect 158529 78510 158668 78512
rect 158529 78507 158595 78510
rect 158662 78508 158668 78510
rect 158732 78508 158738 78572
rect 161197 78570 161244 78572
rect 161152 78568 161244 78570
rect 161152 78512 161202 78568
rect 161152 78510 161244 78512
rect 161197 78508 161244 78510
rect 161308 78508 161314 78572
rect 163773 78568 163820 78572
rect 163884 78570 163890 78572
rect 177573 78570 177639 78573
rect 581085 78570 581151 78573
rect 163773 78512 163778 78568
rect 163773 78508 163820 78512
rect 163884 78510 163930 78570
rect 177573 78568 581151 78570
rect 177573 78512 177578 78568
rect 177634 78512 581090 78568
rect 581146 78512 581151 78568
rect 177573 78510 581151 78512
rect 163884 78508 163890 78510
rect 161197 78507 161263 78508
rect 163773 78507 163839 78508
rect 177573 78507 177639 78510
rect 581085 78507 581151 78510
rect 159541 78434 159607 78437
rect 151862 78432 159607 78434
rect 151862 78376 159546 78432
rect 159602 78376 159607 78432
rect 151862 78374 159607 78376
rect 128118 78236 128124 78300
rect 128188 78298 128194 78300
rect 140730 78298 140790 78374
rect 147630 78298 147690 78374
rect 150525 78371 150591 78374
rect 159541 78371 159607 78374
rect 160686 78372 160692 78436
rect 160756 78434 160762 78436
rect 164969 78434 165035 78437
rect 165337 78436 165403 78437
rect 160756 78432 165035 78434
rect 160756 78376 164974 78432
rect 165030 78376 165035 78432
rect 160756 78374 165035 78376
rect 160756 78372 160762 78374
rect 164969 78371 165035 78374
rect 165286 78372 165292 78436
rect 165356 78434 165403 78436
rect 178033 78434 178099 78437
rect 178166 78434 178172 78436
rect 165356 78432 165448 78434
rect 165398 78376 165448 78432
rect 165356 78374 165448 78376
rect 178033 78432 178172 78434
rect 178033 78376 178038 78432
rect 178094 78376 178172 78432
rect 178033 78374 178172 78376
rect 165356 78372 165403 78374
rect 165337 78371 165403 78372
rect 178033 78371 178099 78374
rect 178166 78372 178172 78374
rect 178236 78372 178242 78436
rect 178309 78434 178375 78437
rect 198733 78434 198799 78437
rect 178309 78432 198799 78434
rect 178309 78376 178314 78432
rect 178370 78376 198738 78432
rect 198794 78376 198799 78432
rect 178309 78374 198799 78376
rect 178309 78371 178375 78374
rect 198733 78371 198799 78374
rect 160461 78298 160527 78301
rect 128188 78238 140790 78298
rect 142846 78238 147690 78298
rect 150206 78296 160527 78298
rect 150206 78240 160466 78296
rect 160522 78240 160527 78296
rect 150206 78238 160527 78240
rect 128188 78236 128194 78238
rect 132166 78100 132172 78164
rect 132236 78162 132242 78164
rect 142846 78162 142906 78238
rect 149513 78162 149579 78165
rect 132236 78102 142906 78162
rect 143490 78160 149579 78162
rect 143490 78104 149518 78160
rect 149574 78104 149579 78160
rect 143490 78102 149579 78104
rect 132236 78100 132242 78102
rect 130878 77964 130884 78028
rect 130948 78026 130954 78028
rect 137829 78026 137895 78029
rect 143490 78026 143550 78102
rect 149513 78099 149579 78102
rect 130948 78024 137895 78026
rect 130948 77968 137834 78024
rect 137890 77968 137895 78024
rect 130948 77966 137895 77968
rect 130948 77964 130954 77966
rect 137829 77963 137895 77966
rect 137970 77966 143550 78026
rect 131982 77828 131988 77892
rect 132052 77890 132058 77892
rect 137970 77890 138030 77966
rect 147990 77964 147996 78028
rect 148060 78026 148066 78028
rect 148501 78026 148567 78029
rect 148060 78024 148567 78026
rect 148060 77968 148506 78024
rect 148562 77968 148567 78024
rect 148060 77966 148567 77968
rect 148060 77964 148066 77966
rect 148501 77963 148567 77966
rect 148910 77964 148916 78028
rect 148980 78026 148986 78028
rect 150206 78026 150266 78238
rect 160461 78235 160527 78238
rect 160870 78236 160876 78300
rect 160940 78298 160946 78300
rect 161197 78298 161263 78301
rect 160940 78296 161263 78298
rect 160940 78240 161202 78296
rect 161258 78240 161263 78296
rect 160940 78238 161263 78240
rect 160940 78236 160946 78238
rect 161197 78235 161263 78238
rect 173382 78236 173388 78300
rect 173452 78298 173458 78300
rect 200665 78298 200731 78301
rect 173452 78296 209790 78298
rect 173452 78240 200670 78296
rect 200726 78240 209790 78296
rect 173452 78238 209790 78240
rect 173452 78236 173458 78238
rect 200665 78235 200731 78238
rect 154297 78164 154363 78165
rect 158529 78164 158595 78165
rect 154246 78162 154252 78164
rect 154206 78102 154252 78162
rect 154316 78160 154363 78164
rect 154358 78104 154363 78160
rect 154246 78100 154252 78102
rect 154316 78100 154363 78104
rect 158478 78100 158484 78164
rect 158548 78162 158595 78164
rect 164785 78162 164851 78165
rect 166390 78162 166396 78164
rect 158548 78160 158640 78162
rect 158590 78104 158640 78160
rect 158548 78102 158640 78104
rect 164785 78160 166396 78162
rect 164785 78104 164790 78160
rect 164846 78104 166396 78160
rect 164785 78102 166396 78104
rect 158548 78100 158595 78102
rect 154297 78099 154363 78100
rect 158529 78099 158595 78100
rect 164785 78099 164851 78102
rect 166390 78100 166396 78102
rect 166460 78100 166466 78164
rect 177021 78162 177087 78165
rect 204437 78162 204503 78165
rect 177021 78160 204503 78162
rect 177021 78104 177026 78160
rect 177082 78104 204442 78160
rect 204498 78104 204503 78160
rect 177021 78102 204503 78104
rect 177021 78099 177087 78102
rect 204437 78099 204503 78102
rect 148980 77966 150266 78026
rect 148980 77964 148986 77966
rect 164918 77964 164924 78028
rect 164988 78026 164994 78028
rect 165245 78026 165311 78029
rect 164988 78024 165311 78026
rect 164988 77968 165250 78024
rect 165306 77968 165311 78024
rect 164988 77966 165311 77968
rect 164988 77964 164994 77966
rect 165245 77963 165311 77966
rect 166441 78026 166507 78029
rect 166574 78026 166580 78028
rect 166441 78024 166580 78026
rect 166441 77968 166446 78024
rect 166502 77968 166580 78024
rect 166441 77966 166580 77968
rect 166441 77963 166507 77966
rect 166574 77964 166580 77966
rect 166644 77964 166650 78028
rect 171542 77964 171548 78028
rect 171612 78026 171618 78028
rect 172329 78026 172395 78029
rect 203190 78026 203196 78028
rect 171612 78024 172395 78026
rect 171612 77968 172334 78024
rect 172390 77968 172395 78024
rect 171612 77966 172395 77968
rect 171612 77964 171618 77966
rect 172329 77963 172395 77966
rect 186270 77966 203196 78026
rect 132052 77830 138030 77890
rect 138197 77892 138263 77893
rect 138197 77888 138244 77892
rect 138308 77890 138314 77892
rect 138749 77890 138815 77893
rect 148593 77890 148659 77893
rect 138197 77832 138202 77888
rect 132052 77828 132058 77830
rect 138197 77828 138244 77832
rect 138308 77830 138354 77890
rect 138749 77888 148659 77890
rect 138749 77832 138754 77888
rect 138810 77832 148598 77888
rect 148654 77832 148659 77888
rect 138749 77830 148659 77832
rect 138308 77828 138314 77830
rect 138197 77827 138263 77828
rect 138749 77827 138815 77830
rect 148593 77827 148659 77830
rect 153694 77828 153700 77892
rect 153764 77890 153770 77892
rect 154389 77890 154455 77893
rect 153764 77888 154455 77890
rect 153764 77832 154394 77888
rect 154450 77832 154455 77888
rect 153764 77830 154455 77832
rect 153764 77828 153770 77830
rect 154389 77827 154455 77830
rect 176837 77890 176903 77893
rect 177665 77890 177731 77893
rect 186270 77890 186330 77966
rect 203190 77964 203196 77966
rect 203260 77964 203266 78028
rect 176837 77888 186330 77890
rect 176837 77832 176842 77888
rect 176898 77832 177670 77888
rect 177726 77832 186330 77888
rect 176837 77830 186330 77832
rect 209730 77890 209790 78238
rect 264237 77890 264303 77893
rect 209730 77888 264303 77890
rect 209730 77832 264242 77888
rect 264298 77832 264303 77888
rect 209730 77830 264303 77832
rect 176837 77827 176903 77830
rect 177665 77827 177731 77830
rect 264237 77827 264303 77830
rect 134057 77756 134123 77757
rect 135161 77756 135227 77757
rect 134006 77754 134012 77756
rect 133966 77694 134012 77754
rect 134076 77752 134123 77756
rect 134118 77696 134123 77752
rect 134006 77692 134012 77694
rect 134076 77692 134123 77696
rect 135110 77692 135116 77756
rect 135180 77754 135227 77756
rect 135437 77754 135503 77757
rect 138105 77756 138171 77757
rect 135846 77754 135852 77756
rect 135180 77752 135272 77754
rect 135222 77696 135272 77752
rect 135180 77694 135272 77696
rect 135437 77752 135852 77754
rect 135437 77696 135442 77752
rect 135498 77696 135852 77752
rect 135437 77694 135852 77696
rect 135180 77692 135227 77694
rect 134057 77691 134123 77692
rect 135161 77691 135227 77692
rect 135437 77691 135503 77694
rect 135846 77692 135852 77694
rect 135916 77692 135922 77756
rect 138054 77754 138060 77756
rect 138014 77694 138060 77754
rect 138124 77752 138171 77756
rect 138166 77696 138171 77752
rect 138054 77692 138060 77694
rect 138124 77692 138171 77696
rect 138105 77691 138171 77692
rect 139485 77754 139551 77757
rect 139710 77754 139716 77756
rect 139485 77752 139716 77754
rect 139485 77696 139490 77752
rect 139546 77696 139716 77752
rect 139485 77694 139716 77696
rect 139485 77691 139551 77694
rect 139710 77692 139716 77694
rect 139780 77692 139786 77756
rect 141049 77754 141115 77757
rect 143758 77754 143764 77756
rect 141049 77752 143764 77754
rect 141049 77696 141054 77752
rect 141110 77696 143764 77752
rect 141049 77694 143764 77696
rect 141049 77691 141115 77694
rect 143758 77692 143764 77694
rect 143828 77692 143834 77756
rect 145230 77692 145236 77756
rect 145300 77754 145306 77756
rect 162945 77754 163011 77757
rect 145300 77752 163011 77754
rect 145300 77696 162950 77752
rect 163006 77696 163011 77752
rect 145300 77694 163011 77696
rect 145300 77692 145306 77694
rect 162945 77691 163011 77694
rect 135345 77618 135411 77621
rect 136398 77618 136404 77620
rect 135345 77616 136404 77618
rect 135345 77560 135350 77616
rect 135406 77560 136404 77616
rect 135345 77558 136404 77560
rect 135345 77555 135411 77558
rect 136398 77556 136404 77558
rect 136468 77556 136474 77620
rect 139577 77618 139643 77621
rect 140957 77620 141023 77621
rect 139894 77618 139900 77620
rect 139577 77616 139900 77618
rect 139577 77560 139582 77616
rect 139638 77560 139900 77616
rect 139577 77558 139900 77560
rect 139577 77555 139643 77558
rect 139894 77556 139900 77558
rect 139964 77556 139970 77620
rect 140957 77616 141004 77620
rect 141068 77618 141074 77620
rect 140957 77560 140962 77616
rect 140957 77556 141004 77560
rect 141068 77558 141114 77618
rect 141068 77556 141074 77558
rect 162710 77556 162716 77620
rect 162780 77618 162786 77620
rect 162853 77618 162919 77621
rect 162780 77616 162919 77618
rect 162780 77560 162858 77616
rect 162914 77560 162919 77616
rect 162780 77558 162919 77560
rect 162780 77556 162786 77558
rect 140957 77555 141023 77556
rect 162853 77555 162919 77558
rect 175825 77618 175891 77621
rect 176193 77618 176259 77621
rect 175825 77616 176259 77618
rect 175825 77560 175830 77616
rect 175886 77560 176198 77616
rect 176254 77560 176259 77616
rect 175825 77558 176259 77560
rect 175825 77555 175891 77558
rect 176193 77555 176259 77558
rect 177389 77618 177455 77621
rect 201718 77618 201724 77620
rect 177389 77616 201724 77618
rect 177389 77560 177394 77616
rect 177450 77560 201724 77616
rect 177389 77558 201724 77560
rect 177389 77555 177455 77558
rect 201718 77556 201724 77558
rect 201788 77556 201794 77620
rect 135294 77420 135300 77484
rect 135364 77482 135370 77484
rect 135805 77482 135871 77485
rect 135364 77480 135871 77482
rect 135364 77424 135810 77480
rect 135866 77424 135871 77480
rect 135364 77422 135871 77424
rect 135364 77420 135370 77422
rect 135805 77419 135871 77422
rect 140078 77420 140084 77484
rect 140148 77482 140154 77484
rect 178585 77482 178651 77485
rect 199101 77482 199167 77485
rect 140148 77422 140790 77482
rect 140148 77420 140154 77422
rect 127566 77284 127572 77348
rect 127636 77346 127642 77348
rect 138749 77346 138815 77349
rect 127636 77344 138815 77346
rect 127636 77288 138754 77344
rect 138810 77288 138815 77344
rect 127636 77286 138815 77288
rect 140730 77346 140790 77422
rect 178585 77480 199167 77482
rect 178585 77424 178590 77480
rect 178646 77424 199106 77480
rect 199162 77424 199167 77480
rect 178585 77422 199167 77424
rect 178585 77419 178651 77422
rect 199101 77419 199167 77422
rect 145649 77346 145715 77349
rect 140730 77344 145715 77346
rect 140730 77288 145654 77344
rect 145710 77288 145715 77344
rect 140730 77286 145715 77288
rect 127636 77284 127642 77286
rect 138749 77283 138815 77286
rect 145649 77283 145715 77286
rect 150525 77346 150591 77349
rect 150985 77346 151051 77349
rect 150525 77344 151051 77346
rect 150525 77288 150530 77344
rect 150586 77288 150990 77344
rect 151046 77288 151051 77344
rect 150525 77286 151051 77288
rect 150525 77283 150591 77286
rect 150985 77283 151051 77286
rect 175825 77346 175891 77349
rect 175958 77346 175964 77348
rect 175825 77344 175964 77346
rect 175825 77288 175830 77344
rect 175886 77288 175964 77344
rect 175825 77286 175964 77288
rect 175825 77283 175891 77286
rect 175958 77284 175964 77286
rect 176028 77284 176034 77348
rect 179413 77346 179479 77349
rect 179638 77346 179644 77348
rect 179413 77344 179644 77346
rect 179413 77288 179418 77344
rect 179474 77288 179644 77344
rect 179413 77286 179644 77288
rect 179413 77283 179479 77286
rect 179638 77284 179644 77286
rect 179708 77346 179714 77348
rect 180333 77346 180399 77349
rect 179708 77344 180399 77346
rect 179708 77288 180338 77344
rect 180394 77288 180399 77344
rect 179708 77286 180399 77288
rect 179708 77284 179714 77286
rect 180333 77283 180399 77286
rect 104157 77210 104223 77213
rect 138013 77210 138079 77213
rect 104157 77208 138079 77210
rect 104157 77152 104162 77208
rect 104218 77152 138018 77208
rect 138074 77152 138079 77208
rect 104157 77150 138079 77152
rect 104157 77147 104223 77150
rect 138013 77147 138079 77150
rect 163262 77148 163268 77212
rect 163332 77210 163338 77212
rect 164141 77210 164207 77213
rect 163332 77208 164207 77210
rect 163332 77152 164146 77208
rect 164202 77152 164207 77208
rect 163332 77150 164207 77152
rect 163332 77148 163338 77150
rect 164141 77147 164207 77150
rect 175958 77148 175964 77212
rect 176028 77210 176034 77212
rect 176561 77210 176627 77213
rect 179873 77212 179939 77213
rect 181345 77212 181411 77213
rect 179822 77210 179828 77212
rect 176028 77208 176627 77210
rect 176028 77152 176566 77208
rect 176622 77152 176627 77208
rect 176028 77150 176627 77152
rect 179782 77150 179828 77210
rect 179892 77208 179939 77212
rect 181294 77210 181300 77212
rect 179934 77152 179939 77208
rect 176028 77148 176034 77150
rect 176561 77147 176627 77150
rect 179822 77148 179828 77150
rect 179892 77148 179939 77152
rect 181254 77150 181300 77210
rect 181364 77208 181411 77212
rect 181406 77152 181411 77208
rect 181294 77148 181300 77150
rect 181364 77148 181411 77152
rect 179873 77147 179939 77148
rect 181345 77147 181411 77148
rect 115749 77074 115815 77077
rect 162485 77076 162551 77077
rect 147622 77074 147628 77076
rect 115749 77072 147628 77074
rect 115749 77016 115754 77072
rect 115810 77016 147628 77072
rect 115749 77014 147628 77016
rect 115749 77011 115815 77014
rect 147622 77012 147628 77014
rect 147692 77012 147698 77076
rect 162485 77074 162532 77076
rect 162440 77072 162532 77074
rect 162440 77016 162490 77072
rect 162440 77014 162532 77016
rect 162485 77012 162532 77014
rect 162596 77012 162602 77076
rect 174486 77012 174492 77076
rect 174556 77074 174562 77076
rect 175181 77074 175247 77077
rect 174556 77072 175247 77074
rect 174556 77016 175186 77072
rect 175242 77016 175247 77072
rect 174556 77014 175247 77016
rect 174556 77012 174562 77014
rect 162485 77011 162551 77012
rect 175181 77011 175247 77014
rect 176469 77076 176535 77077
rect 176469 77072 176516 77076
rect 176580 77074 176586 77076
rect 176837 77074 176903 77077
rect 204345 77074 204411 77077
rect 176469 77016 176474 77072
rect 176469 77012 176516 77016
rect 176580 77014 176626 77074
rect 176837 77072 204411 77074
rect 176837 77016 176842 77072
rect 176898 77016 204350 77072
rect 204406 77016 204411 77072
rect 176837 77014 204411 77016
rect 176580 77012 176586 77014
rect 176469 77011 176535 77012
rect 176837 77011 176903 77014
rect 204345 77011 204411 77014
rect 111793 76938 111859 76941
rect 112345 76938 112411 76941
rect 141233 76938 141299 76941
rect 111793 76936 141299 76938
rect 111793 76880 111798 76936
rect 111854 76880 112350 76936
rect 112406 76880 141238 76936
rect 141294 76880 141299 76936
rect 111793 76878 141299 76880
rect 111793 76875 111859 76878
rect 112345 76875 112411 76878
rect 141233 76875 141299 76878
rect 162342 76876 162348 76940
rect 162412 76938 162418 76940
rect 162485 76938 162551 76941
rect 162412 76936 162551 76938
rect 162412 76880 162490 76936
rect 162546 76880 162551 76936
rect 162412 76878 162551 76880
rect 162412 76876 162418 76878
rect 162485 76875 162551 76878
rect 162669 76938 162735 76941
rect 192109 76938 192175 76941
rect 162669 76936 192175 76938
rect 162669 76880 162674 76936
rect 162730 76880 192114 76936
rect 192170 76880 192175 76936
rect 162669 76878 192175 76880
rect 162669 76875 162735 76878
rect 192109 76875 192175 76878
rect 119889 76802 119955 76805
rect 142654 76802 142660 76804
rect 119889 76800 142660 76802
rect 119889 76744 119894 76800
rect 119950 76744 142660 76800
rect 119889 76742 142660 76744
rect 119889 76739 119955 76742
rect 142654 76740 142660 76742
rect 142724 76802 142730 76804
rect 145741 76802 145807 76805
rect 142724 76800 145807 76802
rect 142724 76744 145746 76800
rect 145802 76744 145807 76800
rect 142724 76742 145807 76744
rect 142724 76740 142730 76742
rect 145741 76739 145807 76742
rect 152958 76740 152964 76804
rect 153028 76802 153034 76804
rect 153285 76802 153351 76805
rect 153028 76800 153351 76802
rect 153028 76744 153290 76800
rect 153346 76744 153351 76800
rect 153028 76742 153351 76744
rect 153028 76740 153034 76742
rect 153285 76739 153351 76742
rect 174118 76740 174124 76804
rect 174188 76802 174194 76804
rect 175181 76802 175247 76805
rect 203609 76802 203675 76805
rect 174188 76800 203675 76802
rect 174188 76744 175186 76800
rect 175242 76744 203614 76800
rect 203670 76744 203675 76800
rect 174188 76742 203675 76744
rect 174188 76740 174194 76742
rect 175181 76739 175247 76742
rect 203609 76739 203675 76742
rect 109769 76666 109835 76669
rect 131113 76666 131179 76669
rect 131573 76666 131639 76669
rect 109769 76664 131639 76666
rect 109769 76608 109774 76664
rect 109830 76608 131118 76664
rect 131174 76608 131578 76664
rect 131634 76608 131639 76664
rect 109769 76606 131639 76608
rect 109769 76603 109835 76606
rect 131113 76603 131179 76606
rect 131573 76603 131639 76606
rect 135345 76666 135411 76669
rect 142889 76668 142955 76669
rect 136214 76666 136220 76668
rect 135345 76664 136220 76666
rect 135345 76608 135350 76664
rect 135406 76608 136220 76664
rect 135345 76606 136220 76608
rect 135345 76603 135411 76606
rect 136214 76604 136220 76606
rect 136284 76604 136290 76668
rect 142838 76604 142844 76668
rect 142908 76666 142955 76668
rect 146845 76668 146911 76669
rect 142908 76664 143000 76666
rect 142950 76608 143000 76664
rect 142908 76606 143000 76608
rect 146845 76664 146892 76668
rect 146956 76666 146962 76668
rect 154021 76666 154087 76669
rect 154246 76666 154252 76668
rect 146845 76608 146850 76664
rect 142908 76604 142955 76606
rect 142889 76603 142955 76604
rect 146845 76604 146892 76608
rect 146956 76606 147002 76666
rect 154021 76664 154252 76666
rect 154021 76608 154026 76664
rect 154082 76608 154252 76664
rect 154021 76606 154252 76608
rect 146956 76604 146962 76606
rect 146845 76603 146911 76604
rect 154021 76603 154087 76606
rect 154246 76604 154252 76606
rect 154316 76604 154322 76668
rect 173341 76666 173407 76669
rect 174077 76666 174143 76669
rect 195329 76666 195395 76669
rect 173341 76664 195395 76666
rect 173341 76608 173346 76664
rect 173402 76608 174082 76664
rect 174138 76608 195334 76664
rect 195390 76608 195395 76664
rect 173341 76606 195395 76608
rect 173341 76603 173407 76606
rect 174077 76603 174143 76606
rect 195329 76603 195395 76606
rect 167177 76530 167243 76533
rect 167310 76530 167316 76532
rect 167177 76528 167316 76530
rect 167177 76472 167182 76528
rect 167238 76472 167316 76528
rect 167177 76470 167316 76472
rect 167177 76467 167243 76470
rect 167310 76468 167316 76470
rect 167380 76468 167386 76532
rect 169845 76530 169911 76533
rect 186998 76530 187004 76532
rect 169845 76528 187004 76530
rect 169845 76472 169850 76528
rect 169906 76472 187004 76528
rect 169845 76470 187004 76472
rect 169845 76467 169911 76470
rect 186998 76468 187004 76470
rect 187068 76530 187074 76532
rect 187550 76530 187556 76532
rect 187068 76470 187556 76530
rect 187068 76468 187074 76470
rect 187550 76468 187556 76470
rect 187620 76468 187626 76532
rect 192109 76530 192175 76533
rect 192937 76530 193003 76533
rect 389173 76530 389239 76533
rect 192109 76528 389239 76530
rect 192109 76472 192114 76528
rect 192170 76472 192942 76528
rect 192998 76472 389178 76528
rect 389234 76472 389239 76528
rect 192109 76470 389239 76472
rect 192109 76467 192175 76470
rect 192937 76467 193003 76470
rect 389173 76467 389239 76470
rect 147438 76332 147444 76396
rect 147508 76394 147514 76396
rect 147806 76394 147812 76396
rect 147508 76334 147812 76394
rect 147508 76332 147514 76334
rect 147806 76332 147812 76334
rect 147876 76332 147882 76396
rect 149605 76394 149671 76397
rect 179454 76394 179460 76396
rect 149605 76392 179460 76394
rect 149605 76336 149610 76392
rect 149666 76336 179460 76392
rect 149605 76334 179460 76336
rect 149605 76331 149671 76334
rect 179454 76332 179460 76334
rect 179524 76332 179530 76396
rect 145230 76196 145236 76260
rect 145300 76258 145306 76260
rect 146017 76258 146083 76261
rect 145300 76256 146083 76258
rect 145300 76200 146022 76256
rect 146078 76200 146083 76256
rect 145300 76198 146083 76200
rect 145300 76196 145306 76198
rect 146017 76195 146083 76198
rect 149329 76258 149395 76261
rect 183686 76258 183692 76260
rect 149329 76256 183692 76258
rect 149329 76200 149334 76256
rect 149390 76200 183692 76256
rect 149329 76198 183692 76200
rect 149329 76195 149395 76198
rect 183686 76196 183692 76198
rect 183756 76196 183762 76260
rect 167310 76060 167316 76124
rect 167380 76122 167386 76124
rect 167821 76122 167887 76125
rect 167380 76120 167887 76122
rect 167380 76064 167826 76120
rect 167882 76064 167887 76120
rect 167380 76062 167887 76064
rect 167380 76060 167386 76062
rect 167821 76059 167887 76062
rect 170070 76060 170076 76124
rect 170140 76122 170146 76124
rect 170765 76122 170831 76125
rect 170140 76120 170831 76122
rect 170140 76064 170770 76120
rect 170826 76064 170831 76120
rect 170140 76062 170831 76064
rect 170140 76060 170146 76062
rect 170765 76059 170831 76062
rect 133822 75924 133828 75988
rect 133892 75986 133898 75988
rect 135069 75986 135135 75989
rect 133892 75984 135135 75986
rect 133892 75928 135074 75984
rect 135130 75928 135135 75984
rect 133892 75926 135135 75928
rect 133892 75924 133898 75926
rect 135069 75923 135135 75926
rect 142705 75986 142771 75989
rect 143165 75988 143231 75989
rect 143022 75986 143028 75988
rect 142705 75984 143028 75986
rect 142705 75928 142710 75984
rect 142766 75928 143028 75984
rect 142705 75926 143028 75928
rect 142705 75923 142771 75926
rect 143022 75924 143028 75926
rect 143092 75924 143098 75988
rect 143165 75984 143212 75988
rect 143276 75986 143282 75988
rect 152365 75986 152431 75989
rect 152590 75986 152596 75988
rect 143165 75928 143170 75984
rect 143165 75924 143212 75928
rect 143276 75926 143322 75986
rect 152365 75984 152596 75986
rect 152365 75928 152370 75984
rect 152426 75928 152596 75984
rect 152365 75926 152596 75928
rect 143276 75924 143282 75926
rect 143165 75923 143231 75924
rect 152365 75923 152431 75926
rect 152590 75924 152596 75926
rect 152660 75924 152666 75988
rect 159030 75924 159036 75988
rect 159100 75986 159106 75988
rect 160001 75986 160067 75989
rect 159100 75984 160067 75986
rect 159100 75928 160006 75984
rect 160062 75928 160067 75984
rect 159100 75926 160067 75928
rect 159100 75924 159106 75926
rect 160001 75923 160067 75926
rect 160829 75988 160895 75989
rect 160829 75984 160876 75988
rect 160940 75986 160946 75988
rect 160829 75928 160834 75984
rect 160829 75924 160876 75928
rect 160940 75926 160986 75986
rect 160940 75924 160946 75926
rect 166206 75924 166212 75988
rect 166276 75986 166282 75988
rect 166901 75986 166967 75989
rect 166276 75984 166967 75986
rect 166276 75928 166906 75984
rect 166962 75928 166967 75984
rect 166276 75926 166967 75928
rect 166276 75924 166282 75926
rect 160829 75923 160895 75924
rect 166901 75923 166967 75926
rect 167678 75924 167684 75988
rect 167748 75986 167754 75988
rect 168373 75986 168439 75989
rect 167748 75984 168439 75986
rect 167748 75928 168378 75984
rect 168434 75928 168439 75984
rect 167748 75926 168439 75928
rect 167748 75924 167754 75926
rect 168373 75923 168439 75926
rect 171225 75986 171291 75989
rect 172053 75988 172119 75989
rect 171726 75986 171732 75988
rect 171225 75984 171732 75986
rect 171225 75928 171230 75984
rect 171286 75928 171732 75984
rect 171225 75926 171732 75928
rect 171225 75923 171291 75926
rect 171726 75924 171732 75926
rect 171796 75924 171802 75988
rect 172053 75984 172100 75988
rect 172164 75986 172170 75988
rect 172053 75928 172058 75984
rect 172053 75924 172100 75928
rect 172164 75926 172210 75986
rect 172164 75924 172170 75926
rect 172053 75923 172119 75924
rect 112805 75850 112871 75853
rect 156781 75852 156847 75853
rect 147806 75850 147812 75852
rect 112805 75848 147812 75850
rect 112805 75792 112810 75848
rect 112866 75792 147812 75848
rect 112805 75790 147812 75792
rect 112805 75787 112871 75790
rect 147806 75788 147812 75790
rect 147876 75788 147882 75852
rect 156781 75848 156828 75852
rect 156892 75850 156898 75852
rect 156781 75792 156786 75848
rect 156781 75788 156828 75792
rect 156892 75790 156938 75850
rect 156892 75788 156898 75790
rect 167862 75788 167868 75852
rect 167932 75850 167938 75852
rect 168005 75850 168071 75853
rect 167932 75848 168071 75850
rect 167932 75792 168010 75848
rect 168066 75792 168071 75848
rect 167932 75790 168071 75792
rect 167932 75788 167938 75790
rect 156781 75787 156847 75788
rect 168005 75787 168071 75790
rect 172697 75850 172763 75853
rect 206001 75850 206067 75853
rect 172697 75848 209790 75850
rect 172697 75792 172702 75848
rect 172758 75792 206006 75848
rect 206062 75792 209790 75848
rect 172697 75790 209790 75792
rect 172697 75787 172763 75790
rect 206001 75787 206067 75790
rect 107101 75714 107167 75717
rect 138054 75714 138060 75716
rect 107101 75712 138060 75714
rect 107101 75656 107106 75712
rect 107162 75656 138060 75712
rect 107101 75654 138060 75656
rect 107101 75651 107167 75654
rect 138054 75652 138060 75654
rect 138124 75652 138130 75716
rect 160369 75714 160435 75717
rect 160686 75714 160692 75716
rect 160369 75712 160692 75714
rect 160369 75656 160374 75712
rect 160430 75656 160692 75712
rect 160369 75654 160692 75656
rect 160369 75651 160435 75654
rect 160686 75652 160692 75654
rect 160756 75652 160762 75716
rect 167269 75714 167335 75717
rect 168046 75714 168052 75716
rect 167269 75712 168052 75714
rect 167269 75656 167274 75712
rect 167330 75656 168052 75712
rect 167269 75654 168052 75656
rect 167269 75651 167335 75654
rect 168046 75652 168052 75654
rect 168116 75652 168122 75716
rect 175549 75714 175615 75717
rect 176561 75714 176627 75717
rect 206185 75714 206251 75717
rect 175549 75712 206251 75714
rect 175549 75656 175554 75712
rect 175610 75656 176566 75712
rect 176622 75656 206190 75712
rect 206246 75656 206251 75712
rect 175549 75654 206251 75656
rect 175549 75651 175615 75654
rect 176561 75651 176627 75654
rect 206185 75651 206251 75654
rect 114369 75578 114435 75581
rect 145230 75578 145236 75580
rect 114369 75576 145236 75578
rect 114369 75520 114374 75576
rect 114430 75520 145236 75576
rect 114369 75518 145236 75520
rect 114369 75515 114435 75518
rect 145230 75516 145236 75518
rect 145300 75516 145306 75580
rect 156873 75578 156939 75581
rect 185342 75578 185348 75580
rect 156873 75576 185348 75578
rect 156873 75520 156878 75576
rect 156934 75520 185348 75576
rect 156873 75518 185348 75520
rect 156873 75515 156939 75518
rect 185342 75516 185348 75518
rect 185412 75516 185418 75580
rect 108481 75442 108547 75445
rect 138422 75442 138428 75444
rect 108481 75440 138428 75442
rect 108481 75384 108486 75440
rect 108542 75384 138428 75440
rect 108481 75382 138428 75384
rect 108481 75379 108547 75382
rect 138422 75380 138428 75382
rect 138492 75380 138498 75444
rect 173709 75442 173775 75445
rect 189022 75442 189028 75444
rect 173709 75440 189028 75442
rect 173709 75384 173714 75440
rect 173770 75384 189028 75440
rect 173709 75382 189028 75384
rect 173709 75379 173775 75382
rect 189022 75380 189028 75382
rect 189092 75442 189098 75444
rect 190310 75442 190316 75444
rect 189092 75382 190316 75442
rect 189092 75380 189098 75382
rect 190310 75380 190316 75382
rect 190380 75380 190386 75444
rect 22737 75306 22803 75309
rect 134374 75306 134380 75308
rect 22737 75304 134380 75306
rect 22737 75248 22742 75304
rect 22798 75248 134380 75304
rect 22737 75246 134380 75248
rect 22737 75243 22803 75246
rect 134374 75244 134380 75246
rect 134444 75244 134450 75308
rect 173985 75306 174051 75309
rect 174721 75306 174787 75309
rect 188521 75306 188587 75309
rect 173985 75304 188587 75306
rect 173985 75248 173990 75304
rect 174046 75248 174726 75304
rect 174782 75248 188526 75304
rect 188582 75248 188587 75304
rect 173985 75246 188587 75248
rect 209730 75306 209790 75790
rect 475377 75306 475443 75309
rect 209730 75304 475443 75306
rect 209730 75248 475382 75304
rect 475438 75248 475443 75304
rect 209730 75246 475443 75248
rect 173985 75243 174051 75246
rect 174721 75243 174787 75246
rect 188521 75243 188587 75246
rect 475377 75243 475443 75246
rect 7557 75170 7623 75173
rect 120022 75170 120028 75172
rect 7557 75168 120028 75170
rect 7557 75112 7562 75168
rect 7618 75112 120028 75168
rect 7557 75110 120028 75112
rect 7557 75107 7623 75110
rect 120022 75108 120028 75110
rect 120092 75108 120098 75172
rect 173065 75170 173131 75173
rect 173750 75170 173756 75172
rect 173065 75168 173756 75170
rect 173065 75112 173070 75168
rect 173126 75112 173756 75168
rect 173065 75110 173756 75112
rect 173065 75107 173131 75110
rect 173750 75108 173756 75110
rect 173820 75108 173826 75172
rect 175457 75170 175523 75173
rect 176326 75170 176332 75172
rect 175457 75168 176332 75170
rect 175457 75112 175462 75168
rect 175518 75112 176332 75168
rect 175457 75110 176332 75112
rect 175457 75107 175523 75110
rect 176326 75108 176332 75110
rect 176396 75108 176402 75172
rect 177481 75170 177547 75173
rect 549253 75170 549319 75173
rect 177481 75168 549319 75170
rect 177481 75112 177486 75168
rect 177542 75112 549258 75168
rect 549314 75112 549319 75168
rect 177481 75110 549319 75112
rect 177481 75107 177547 75110
rect 549253 75107 549319 75110
rect 117129 75034 117195 75037
rect 144126 75034 144132 75036
rect 117129 75032 144132 75034
rect 117129 74976 117134 75032
rect 117190 74976 144132 75032
rect 117129 74974 144132 74976
rect 117129 74971 117195 74974
rect 144126 74972 144132 74974
rect 144196 74972 144202 75036
rect 157149 75034 157215 75037
rect 178718 75034 178724 75036
rect 157149 75032 178724 75034
rect 157149 74976 157154 75032
rect 157210 74976 178724 75032
rect 157149 74974 178724 74976
rect 157149 74971 157215 74974
rect 178718 74972 178724 74974
rect 178788 74972 178794 75036
rect 122373 74626 122439 74629
rect 122782 74626 122788 74628
rect 122373 74624 122788 74626
rect 122373 74568 122378 74624
rect 122434 74568 122788 74624
rect 122373 74566 122788 74568
rect 122373 74563 122439 74566
rect 122782 74564 122788 74566
rect 122852 74564 122858 74628
rect 152406 74564 152412 74628
rect 152476 74626 152482 74628
rect 152825 74626 152891 74629
rect 152476 74624 152891 74626
rect 152476 74568 152830 74624
rect 152886 74568 152891 74624
rect 152476 74566 152891 74568
rect 152476 74564 152482 74566
rect 152825 74563 152891 74566
rect 113081 74490 113147 74493
rect 144310 74490 144316 74492
rect 113081 74488 144316 74490
rect 113081 74432 113086 74488
rect 113142 74432 144316 74488
rect 113081 74430 144316 74432
rect 113081 74427 113147 74430
rect 144310 74428 144316 74430
rect 144380 74490 144386 74492
rect 144637 74490 144703 74493
rect 144380 74488 144703 74490
rect 144380 74432 144642 74488
rect 144698 74432 144703 74488
rect 144380 74430 144703 74432
rect 144380 74428 144386 74430
rect 144637 74427 144703 74430
rect 153377 74490 153443 74493
rect 205817 74490 205883 74493
rect 153377 74488 205883 74490
rect 153377 74432 153382 74488
rect 153438 74432 205822 74488
rect 205878 74432 205883 74488
rect 153377 74430 205883 74432
rect 153377 74427 153443 74430
rect 205817 74427 205883 74430
rect 124029 74354 124095 74357
rect 158069 74354 158135 74357
rect 158345 74354 158411 74357
rect 124029 74352 158411 74354
rect 124029 74296 124034 74352
rect 124090 74296 158074 74352
rect 158130 74296 158350 74352
rect 158406 74296 158411 74352
rect 124029 74294 158411 74296
rect 124029 74291 124095 74294
rect 158069 74291 158135 74294
rect 158345 74291 158411 74294
rect 172278 74292 172284 74356
rect 172348 74354 172354 74356
rect 172421 74354 172487 74357
rect 172348 74352 172487 74354
rect 172348 74296 172426 74352
rect 172482 74296 172487 74352
rect 172348 74294 172487 74296
rect 172348 74292 172354 74294
rect 172421 74291 172487 74294
rect 175089 74354 175155 74357
rect 201534 74354 201540 74356
rect 175089 74352 201540 74354
rect 175089 74296 175094 74352
rect 175150 74296 201540 74352
rect 175089 74294 201540 74296
rect 175089 74291 175155 74294
rect 201534 74292 201540 74294
rect 201604 74292 201610 74356
rect 134057 74218 134123 74221
rect 103470 74216 134123 74218
rect 103470 74160 134062 74216
rect 134118 74160 134123 74216
rect 103470 74158 134123 74160
rect 26233 73946 26299 73949
rect 103053 73946 103119 73949
rect 103470 73946 103530 74158
rect 134057 74155 134123 74158
rect 155677 74218 155743 74221
rect 184054 74218 184060 74220
rect 155677 74216 184060 74218
rect 155677 74160 155682 74216
rect 155738 74160 184060 74216
rect 155677 74158 184060 74160
rect 155677 74155 155743 74158
rect 184054 74156 184060 74158
rect 184124 74156 184130 74220
rect 118049 74082 118115 74085
rect 147990 74082 147996 74084
rect 118049 74080 147996 74082
rect 118049 74024 118054 74080
rect 118110 74024 147996 74080
rect 118049 74022 147996 74024
rect 118049 74019 118115 74022
rect 147990 74020 147996 74022
rect 148060 74020 148066 74084
rect 156781 74082 156847 74085
rect 182950 74082 182956 74084
rect 156781 74080 182956 74082
rect 156781 74024 156786 74080
rect 156842 74024 182956 74080
rect 156781 74022 182956 74024
rect 156781 74019 156847 74022
rect 182950 74020 182956 74022
rect 183020 74020 183026 74084
rect 26233 73944 103530 73946
rect 26233 73888 26238 73944
rect 26294 73888 103058 73944
rect 103114 73888 103530 73944
rect 26233 73886 103530 73888
rect 120717 73946 120783 73949
rect 147070 73946 147076 73948
rect 120717 73944 147076 73946
rect 120717 73888 120722 73944
rect 120778 73888 147076 73944
rect 120717 73886 147076 73888
rect 26233 73883 26299 73886
rect 103053 73883 103119 73886
rect 120717 73883 120783 73886
rect 147070 73884 147076 73886
rect 147140 73884 147146 73948
rect 158345 73946 158411 73949
rect 181110 73946 181116 73948
rect 158345 73944 181116 73946
rect 158345 73888 158350 73944
rect 158406 73888 181116 73944
rect 158345 73886 181116 73888
rect 158345 73883 158411 73886
rect 181110 73884 181116 73886
rect 181180 73884 181186 73948
rect 14457 73810 14523 73813
rect 108665 73810 108731 73813
rect 133229 73810 133295 73813
rect 14457 73808 133295 73810
rect 14457 73752 14462 73808
rect 14518 73752 108670 73808
rect 108726 73752 133234 73808
rect 133290 73752 133295 73808
rect 14457 73750 133295 73752
rect 14457 73747 14523 73750
rect 108665 73747 108731 73750
rect 133229 73747 133295 73750
rect 157926 73748 157932 73812
rect 157996 73810 158002 73812
rect 172421 73810 172487 73813
rect 157996 73808 172487 73810
rect 157996 73752 172426 73808
rect 172482 73752 172487 73808
rect 157996 73750 172487 73752
rect 157996 73748 158002 73750
rect 172421 73747 172487 73750
rect 205817 73810 205883 73813
rect 269113 73810 269179 73813
rect 205817 73808 269179 73810
rect 205817 73752 205822 73808
rect 205878 73752 269118 73808
rect 269174 73752 269179 73808
rect 205817 73750 269179 73752
rect 205817 73747 205883 73750
rect 269113 73747 269179 73750
rect 163262 73612 163268 73676
rect 163332 73674 163338 73676
rect 163589 73674 163655 73677
rect 163332 73672 163655 73674
rect 163332 73616 163594 73672
rect 163650 73616 163655 73672
rect 163332 73614 163655 73616
rect 163332 73612 163338 73614
rect 163589 73611 163655 73614
rect 165286 73612 165292 73676
rect 165356 73674 165362 73676
rect 165429 73674 165495 73677
rect 165356 73672 165495 73674
rect 165356 73616 165434 73672
rect 165490 73616 165495 73672
rect 165356 73614 165495 73616
rect 165356 73612 165362 73614
rect 165429 73611 165495 73614
rect 119654 73068 119660 73132
rect 119724 73130 119730 73132
rect 153469 73130 153535 73133
rect 154205 73130 154271 73133
rect 119724 73128 154271 73130
rect 119724 73072 153474 73128
rect 153530 73072 154210 73128
rect 154266 73072 154271 73128
rect 119724 73070 154271 73072
rect 119724 73068 119730 73070
rect 153469 73067 153535 73070
rect 154205 73067 154271 73070
rect 162117 73130 162183 73133
rect 183870 73130 183876 73132
rect 162117 73128 183876 73130
rect 162117 73072 162122 73128
rect 162178 73072 183876 73128
rect 162117 73070 183876 73072
rect 162117 73067 162183 73070
rect 183870 73068 183876 73070
rect 183940 73068 183946 73132
rect 115841 72994 115907 72997
rect 149278 72994 149284 72996
rect 115841 72992 149284 72994
rect 115841 72936 115846 72992
rect 115902 72936 149284 72992
rect 115841 72934 149284 72936
rect 115841 72931 115907 72934
rect 149278 72932 149284 72934
rect 149348 72994 149354 72996
rect 149830 72994 149836 72996
rect 149348 72934 149836 72994
rect 149348 72932 149354 72934
rect 149830 72932 149836 72934
rect 149900 72932 149906 72996
rect 159817 72994 159883 72997
rect 185158 72994 185164 72996
rect 159817 72992 185164 72994
rect 159817 72936 159822 72992
rect 159878 72936 185164 72992
rect 159817 72934 185164 72936
rect 159817 72931 159883 72934
rect 185158 72932 185164 72934
rect 185228 72932 185234 72996
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 124121 72858 124187 72861
rect 157977 72858 158043 72861
rect 124121 72856 158043 72858
rect 124121 72800 124126 72856
rect 124182 72800 157982 72856
rect 158038 72800 158043 72856
rect 583520 72844 584960 72934
rect 124121 72798 158043 72800
rect 124121 72795 124187 72798
rect 157977 72795 158043 72798
rect 106089 72722 106155 72725
rect 139894 72722 139900 72724
rect 106089 72720 139900 72722
rect 106089 72664 106094 72720
rect 106150 72664 139900 72720
rect 106089 72662 139900 72664
rect 106089 72659 106155 72662
rect 139894 72660 139900 72662
rect 139964 72660 139970 72724
rect 158662 72660 158668 72724
rect 158732 72722 158738 72724
rect 182766 72722 182772 72724
rect 158732 72662 182772 72722
rect 158732 72660 158738 72662
rect 182766 72660 182772 72662
rect 182836 72660 182842 72724
rect 118509 72586 118575 72589
rect 148358 72586 148364 72588
rect 118509 72584 148364 72586
rect 118509 72528 118514 72584
rect 118570 72528 148364 72584
rect 118509 72526 148364 72528
rect 118509 72523 118575 72526
rect 148358 72524 148364 72526
rect 148428 72524 148434 72588
rect 158437 72450 158503 72453
rect 162117 72450 162183 72453
rect 158437 72448 162183 72450
rect 158437 72392 158442 72448
rect 158498 72392 162122 72448
rect 162178 72392 162183 72448
rect 158437 72390 162183 72392
rect 158437 72387 158503 72390
rect 162117 72387 162183 72390
rect 105537 71906 105603 71909
rect 106089 71906 106155 71909
rect 105537 71904 106155 71906
rect 105537 71848 105542 71904
rect 105598 71848 106094 71904
rect 106150 71848 106155 71904
rect 105537 71846 106155 71848
rect 105537 71843 105603 71846
rect 106089 71843 106155 71846
rect 109861 71770 109927 71773
rect 144494 71770 144500 71772
rect 109861 71768 144500 71770
rect -960 71634 480 71724
rect 109861 71712 109866 71768
rect 109922 71712 144500 71768
rect 109861 71710 144500 71712
rect 109861 71707 109927 71710
rect 144494 71708 144500 71710
rect 144564 71770 144570 71772
rect 146753 71770 146819 71773
rect 144564 71768 146819 71770
rect 144564 71712 146758 71768
rect 146814 71712 146819 71768
rect 144564 71710 146819 71712
rect 144564 71708 144570 71710
rect 146753 71707 146819 71710
rect 146886 71708 146892 71772
rect 146956 71770 146962 71772
rect 180926 71770 180932 71772
rect 146956 71710 180932 71770
rect 146956 71708 146962 71710
rect 180926 71708 180932 71710
rect 180996 71770 181002 71772
rect 181529 71770 181595 71773
rect 187601 71772 187667 71773
rect 190361 71772 190427 71773
rect 187550 71770 187556 71772
rect 180996 71768 181595 71770
rect 180996 71712 181534 71768
rect 181590 71712 181595 71768
rect 180996 71710 181595 71712
rect 187510 71710 187556 71770
rect 187620 71768 187667 71772
rect 190310 71770 190316 71772
rect 187662 71712 187667 71768
rect 180996 71708 181002 71710
rect 181529 71707 181595 71710
rect 187550 71708 187556 71710
rect 187620 71708 187667 71712
rect 190270 71710 190316 71770
rect 190380 71768 190427 71772
rect 190422 71712 190427 71768
rect 190310 71708 190316 71710
rect 190380 71708 190427 71712
rect 187601 71707 187667 71708
rect 190361 71707 190427 71708
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 116209 71634 116275 71637
rect 151118 71634 151124 71636
rect 116209 71632 151124 71634
rect 116209 71576 116214 71632
rect 116270 71576 151124 71632
rect 116209 71574 151124 71576
rect 116209 71571 116275 71574
rect 151118 71572 151124 71574
rect 151188 71572 151194 71636
rect 175590 71572 175596 71636
rect 175660 71634 175666 71636
rect 200573 71634 200639 71637
rect 201401 71634 201467 71637
rect 175660 71632 201467 71634
rect 175660 71576 200578 71632
rect 200634 71576 201406 71632
rect 201462 71576 201467 71632
rect 175660 71574 201467 71576
rect 175660 71572 175666 71574
rect 200573 71571 200639 71574
rect 201401 71571 201467 71574
rect 121913 71498 121979 71501
rect 152406 71498 152412 71500
rect 121913 71496 152412 71498
rect 121913 71440 121918 71496
rect 121974 71440 152412 71496
rect 121913 71438 152412 71440
rect 121913 71435 121979 71438
rect 152406 71436 152412 71438
rect 152476 71436 152482 71500
rect 177205 71498 177271 71501
rect 182081 71498 182147 71501
rect 177205 71496 182147 71498
rect 177205 71440 177210 71496
rect 177266 71440 182086 71496
rect 182142 71440 182147 71496
rect 177205 71438 182147 71440
rect 177205 71435 177271 71438
rect 182081 71435 182147 71438
rect 121821 71362 121887 71365
rect 149094 71362 149100 71364
rect 121821 71360 149100 71362
rect 121821 71304 121826 71360
rect 121882 71304 149100 71360
rect 121821 71302 149100 71304
rect 121821 71299 121887 71302
rect 149094 71300 149100 71302
rect 149164 71300 149170 71364
rect 183686 71300 183692 71364
rect 183756 71362 183762 71364
rect 218053 71362 218119 71365
rect 183756 71360 218119 71362
rect 183756 71304 218058 71360
rect 218114 71304 218119 71360
rect 183756 71302 218119 71304
rect 183756 71300 183762 71302
rect 218053 71299 218119 71302
rect 112437 71226 112503 71229
rect 138238 71226 138244 71228
rect 112437 71224 138244 71226
rect 112437 71168 112442 71224
rect 112498 71168 138244 71224
rect 112437 71166 138244 71168
rect 112437 71163 112503 71166
rect 138238 71164 138244 71166
rect 138308 71164 138314 71228
rect 171133 71226 171199 71229
rect 190494 71226 190500 71228
rect 171133 71224 190500 71226
rect 171133 71168 171138 71224
rect 171194 71168 190500 71224
rect 171133 71166 190500 71168
rect 171133 71163 171199 71166
rect 190494 71164 190500 71166
rect 190564 71226 190570 71228
rect 494053 71226 494119 71229
rect 190564 71224 494119 71226
rect 190564 71168 494058 71224
rect 494114 71168 494119 71224
rect 190564 71166 494119 71168
rect 190564 71164 190570 71166
rect 494053 71163 494119 71166
rect 182081 71090 182147 71093
rect 189206 71090 189212 71092
rect 182081 71088 189212 71090
rect 182081 71032 182086 71088
rect 182142 71032 189212 71088
rect 182081 71030 189212 71032
rect 182081 71027 182147 71030
rect 189206 71028 189212 71030
rect 189276 71028 189282 71092
rect 201401 71090 201467 71093
rect 543733 71090 543799 71093
rect 201401 71088 543799 71090
rect 201401 71032 201406 71088
rect 201462 71032 543738 71088
rect 543794 71032 543799 71088
rect 201401 71030 543799 71032
rect 201401 71027 201467 71030
rect 543733 71027 543799 71030
rect 122966 70484 122972 70548
rect 123036 70484 123042 70548
rect 147990 70546 147996 70548
rect 147814 70486 147996 70546
rect 122974 70410 123034 70484
rect 142061 70412 142127 70413
rect 147814 70412 147874 70486
rect 147990 70484 147996 70486
rect 148060 70484 148066 70548
rect 124070 70410 124076 70412
rect 122974 70350 124076 70410
rect 124070 70348 124076 70350
rect 124140 70348 124146 70412
rect 142061 70408 142108 70412
rect 142172 70410 142178 70412
rect 142061 70352 142066 70408
rect 142061 70348 142108 70352
rect 142172 70350 142218 70410
rect 142172 70348 142178 70350
rect 147806 70348 147812 70412
rect 147876 70348 147882 70412
rect 199326 70348 199332 70412
rect 199396 70410 199402 70412
rect 199561 70410 199627 70413
rect 199396 70408 199627 70410
rect 199396 70352 199566 70408
rect 199622 70352 199627 70408
rect 199396 70350 199627 70352
rect 199396 70348 199402 70350
rect 142061 70347 142127 70348
rect 199561 70347 199627 70350
rect 119838 70212 119844 70276
rect 119908 70274 119914 70276
rect 153694 70274 153700 70276
rect 119908 70214 153700 70274
rect 119908 70212 119914 70214
rect 153694 70212 153700 70214
rect 153764 70212 153770 70276
rect 172145 70274 172211 70277
rect 172145 70272 180810 70274
rect 172145 70216 172150 70272
rect 172206 70216 180810 70272
rect 172145 70214 180810 70216
rect 172145 70211 172211 70214
rect 122966 70076 122972 70140
rect 123036 70138 123042 70140
rect 156597 70138 156663 70141
rect 123036 70136 156663 70138
rect 123036 70080 156602 70136
rect 156658 70080 156663 70136
rect 123036 70078 156663 70080
rect 123036 70076 123042 70078
rect 156597 70075 156663 70078
rect 124070 69940 124076 70004
rect 124140 70002 124146 70004
rect 153561 70002 153627 70005
rect 154113 70002 154179 70005
rect 124140 70000 154179 70002
rect 124140 69944 153566 70000
rect 153622 69944 154118 70000
rect 154174 69944 154179 70000
rect 124140 69942 154179 69944
rect 124140 69940 124146 69942
rect 153561 69939 153627 69942
rect 154113 69939 154179 69942
rect 180750 69594 180810 70214
rect 194542 69594 194548 69596
rect 180750 69534 194548 69594
rect 194542 69532 194548 69534
rect 194612 69594 194618 69596
rect 498193 69594 498259 69597
rect 194612 69592 498259 69594
rect 194612 69536 498198 69592
rect 498254 69536 498259 69592
rect 194612 69534 498259 69536
rect 194612 69532 194618 69534
rect 498193 69531 498259 69534
rect 196014 68852 196020 68916
rect 196084 68914 196090 68916
rect 196249 68914 196315 68917
rect 196084 68912 196315 68914
rect 196084 68856 196254 68912
rect 196310 68856 196315 68912
rect 196084 68854 196315 68856
rect 196084 68852 196090 68854
rect 196249 68851 196315 68854
rect 174445 68778 174511 68781
rect 201033 68778 201099 68781
rect 201401 68778 201467 68781
rect 174445 68776 201467 68778
rect 174445 68720 174450 68776
rect 174506 68720 201038 68776
rect 201094 68720 201406 68776
rect 201462 68720 201467 68776
rect 174445 68718 201467 68720
rect 174445 68715 174511 68718
rect 201033 68715 201099 68718
rect 201401 68715 201467 68718
rect 179454 68308 179460 68372
rect 179524 68370 179530 68372
rect 220813 68370 220879 68373
rect 179524 68368 220879 68370
rect 179524 68312 220818 68368
rect 220874 68312 220879 68368
rect 179524 68310 220879 68312
rect 179524 68308 179530 68310
rect 220813 68307 220879 68310
rect 8937 68234 9003 68237
rect 131246 68234 131252 68236
rect 8937 68232 131252 68234
rect 8937 68176 8942 68232
rect 8998 68176 131252 68232
rect 8937 68174 131252 68176
rect 8937 68171 9003 68174
rect 131246 68172 131252 68174
rect 131316 68172 131322 68236
rect 147622 68172 147628 68236
rect 147692 68234 147698 68236
rect 192477 68234 192543 68237
rect 147692 68232 192543 68234
rect 147692 68176 192482 68232
rect 192538 68176 192543 68232
rect 147692 68174 192543 68176
rect 147692 68172 147698 68174
rect 192477 68171 192543 68174
rect 201401 68234 201467 68237
rect 539685 68234 539751 68237
rect 201401 68232 539751 68234
rect 201401 68176 201406 68232
rect 201462 68176 539690 68232
rect 539746 68176 539751 68232
rect 201401 68174 539751 68176
rect 201401 68171 201467 68174
rect 539685 68171 539751 68174
rect 110137 67554 110203 67557
rect 143574 67554 143580 67556
rect 110137 67552 143580 67554
rect 110137 67496 110142 67552
rect 110198 67496 143580 67552
rect 110137 67494 143580 67496
rect 110137 67491 110203 67494
rect 143574 67492 143580 67494
rect 143644 67554 143650 67556
rect 144494 67554 144500 67556
rect 143644 67494 144500 67554
rect 143644 67492 143650 67494
rect 144494 67492 144500 67494
rect 144564 67492 144570 67556
rect 164918 67492 164924 67556
rect 164988 67554 164994 67556
rect 189073 67554 189139 67557
rect 189533 67554 189599 67557
rect 200849 67556 200915 67557
rect 200798 67554 200804 67556
rect 164988 67552 189599 67554
rect 164988 67496 189078 67552
rect 189134 67496 189538 67552
rect 189594 67496 189599 67552
rect 164988 67494 189599 67496
rect 200758 67494 200804 67554
rect 200868 67552 200915 67556
rect 200910 67496 200915 67552
rect 164988 67492 164994 67494
rect 189073 67491 189139 67494
rect 189533 67491 189599 67494
rect 200798 67492 200804 67494
rect 200868 67492 200915 67496
rect 200849 67491 200915 67492
rect 102133 67418 102199 67421
rect 103145 67418 103211 67421
rect 135846 67418 135852 67420
rect 102133 67416 135852 67418
rect 102133 67360 102138 67416
rect 102194 67360 103150 67416
rect 103206 67360 135852 67416
rect 102133 67358 135852 67360
rect 102133 67355 102199 67358
rect 103145 67355 103211 67358
rect 135846 67356 135852 67358
rect 135916 67356 135922 67420
rect 139710 67282 139716 67284
rect 113130 67222 139716 67282
rect 93853 67146 93919 67149
rect 108757 67146 108823 67149
rect 113130 67146 113190 67222
rect 139710 67220 139716 67222
rect 139780 67220 139786 67284
rect 147254 67220 147260 67284
rect 147324 67282 147330 67284
rect 193857 67282 193923 67285
rect 147324 67280 193923 67282
rect 147324 67224 193862 67280
rect 193918 67224 193923 67280
rect 147324 67222 193923 67224
rect 147324 67220 147330 67222
rect 193857 67219 193923 67222
rect 93853 67144 113190 67146
rect 93853 67088 93858 67144
rect 93914 67088 108762 67144
rect 108818 67088 113190 67144
rect 93853 67086 113190 67088
rect 114921 67146 114987 67149
rect 140998 67146 141004 67148
rect 114921 67144 141004 67146
rect 114921 67088 114926 67144
rect 114982 67088 141004 67144
rect 114921 67086 141004 67088
rect 93853 67083 93919 67086
rect 108757 67083 108823 67086
rect 114921 67083 114987 67086
rect 140998 67084 141004 67086
rect 141068 67084 141074 67148
rect 147990 67084 147996 67148
rect 148060 67146 148066 67148
rect 213913 67146 213979 67149
rect 148060 67144 213979 67146
rect 148060 67088 213918 67144
rect 213974 67088 213979 67144
rect 148060 67086 213979 67088
rect 148060 67084 148066 67086
rect 213913 67083 213979 67086
rect 40033 67010 40099 67013
rect 102133 67010 102199 67013
rect 40033 67008 102199 67010
rect 40033 66952 40038 67008
rect 40094 66952 102138 67008
rect 102194 66952 102199 67008
rect 40033 66950 102199 66952
rect 40033 66947 40099 66950
rect 102133 66947 102199 66950
rect 110413 67010 110479 67013
rect 142061 67010 142127 67013
rect 110413 67008 142127 67010
rect 110413 66952 110418 67008
rect 110474 66952 142066 67008
rect 142122 66952 142127 67008
rect 110413 66950 142127 66952
rect 110413 66947 110479 66950
rect 142061 66947 142127 66950
rect 189073 67010 189139 67013
rect 423673 67010 423739 67013
rect 189073 67008 423739 67010
rect 189073 66952 189078 67008
rect 189134 66952 423678 67008
rect 423734 66952 423739 67008
rect 189073 66950 423739 66952
rect 189073 66947 189139 66950
rect 423673 66947 423739 66950
rect 11053 66874 11119 66877
rect 133086 66874 133092 66876
rect 11053 66872 133092 66874
rect 11053 66816 11058 66872
rect 11114 66816 133092 66872
rect 11053 66814 133092 66816
rect 11053 66811 11119 66814
rect 133086 66812 133092 66814
rect 133156 66812 133162 66876
rect 170254 66812 170260 66876
rect 170324 66874 170330 66876
rect 496077 66874 496143 66877
rect 170324 66872 496143 66874
rect 170324 66816 496082 66872
rect 496138 66816 496143 66872
rect 170324 66814 496143 66816
rect 170324 66812 170330 66814
rect 496077 66811 496143 66814
rect 194041 66196 194107 66197
rect 171910 66132 171916 66196
rect 171980 66194 171986 66196
rect 193990 66194 193996 66196
rect 171980 66134 180810 66194
rect 193950 66134 193996 66194
rect 194060 66192 194107 66196
rect 194102 66136 194107 66192
rect 171980 66132 171986 66134
rect 180750 65514 180810 66134
rect 193990 66132 193996 66134
rect 194060 66132 194107 66136
rect 194041 66131 194107 66132
rect 193806 65514 193812 65516
rect 180750 65454 193812 65514
rect 193806 65452 193812 65454
rect 193876 65514 193882 65516
rect 507853 65514 507919 65517
rect 193876 65512 507919 65514
rect 193876 65456 507858 65512
rect 507914 65456 507919 65512
rect 193876 65454 507919 65456
rect 193876 65452 193882 65454
rect 507853 65451 507919 65454
rect 110873 64834 110939 64837
rect 139526 64834 139532 64836
rect 110873 64832 139532 64834
rect 110873 64776 110878 64832
rect 110934 64776 139532 64832
rect 110873 64774 139532 64776
rect 110873 64771 110939 64774
rect 139526 64772 139532 64774
rect 139596 64772 139602 64836
rect 152590 64772 152596 64836
rect 152660 64834 152666 64836
rect 186589 64834 186655 64837
rect 152660 64832 186655 64834
rect 152660 64776 186594 64832
rect 186650 64776 186655 64832
rect 152660 64774 186655 64776
rect 152660 64772 152666 64774
rect 186589 64771 186655 64774
rect 172094 64636 172100 64700
rect 172164 64698 172170 64700
rect 197721 64698 197787 64701
rect 172164 64696 197787 64698
rect 172164 64640 197726 64696
rect 197782 64640 197787 64696
rect 172164 64638 197787 64640
rect 172164 64636 172170 64638
rect 197721 64635 197787 64638
rect 174854 64500 174860 64564
rect 174924 64562 174930 64564
rect 174924 64502 180810 64562
rect 174924 64500 174930 64502
rect 92473 64154 92539 64157
rect 110873 64154 110939 64157
rect 92473 64152 110939 64154
rect 92473 64096 92478 64152
rect 92534 64096 110878 64152
rect 110934 64096 110939 64152
rect 92473 64094 110939 64096
rect 180750 64154 180810 64502
rect 186589 64426 186655 64429
rect 256693 64426 256759 64429
rect 186589 64424 256759 64426
rect 186589 64368 186594 64424
rect 186650 64368 256698 64424
rect 256754 64368 256759 64424
rect 186589 64366 256759 64368
rect 186589 64363 186655 64366
rect 256693 64363 256759 64366
rect 197721 64290 197787 64293
rect 511993 64290 512059 64293
rect 197721 64288 512059 64290
rect 197721 64232 197726 64288
rect 197782 64232 511998 64288
rect 512054 64232 512059 64288
rect 197721 64230 512059 64232
rect 197721 64227 197787 64230
rect 511993 64227 512059 64230
rect 191782 64154 191788 64156
rect 180750 64094 191788 64154
rect 92473 64091 92539 64094
rect 110873 64091 110939 64094
rect 191782 64092 191788 64094
rect 191852 64154 191858 64156
rect 547873 64154 547939 64157
rect 191852 64152 547939 64154
rect 191852 64096 547878 64152
rect 547934 64096 547939 64152
rect 191852 64094 547939 64096
rect 191852 64092 191858 64094
rect 547873 64091 547939 64094
rect 152774 63412 152780 63476
rect 152844 63474 152850 63476
rect 205725 63474 205791 63477
rect 152844 63472 209790 63474
rect 152844 63416 205730 63472
rect 205786 63416 209790 63472
rect 152844 63414 209790 63416
rect 152844 63412 152850 63414
rect 205725 63411 205791 63414
rect 165102 63276 165108 63340
rect 165172 63338 165178 63340
rect 199009 63338 199075 63341
rect 199377 63338 199443 63341
rect 165172 63336 199443 63338
rect 165172 63280 199014 63336
rect 199070 63280 199382 63336
rect 199438 63280 199443 63336
rect 165172 63278 199443 63280
rect 209730 63338 209790 63414
rect 259453 63338 259519 63341
rect 209730 63336 259519 63338
rect 209730 63280 259458 63336
rect 259514 63280 259519 63336
rect 209730 63278 259519 63280
rect 165172 63276 165178 63278
rect 199009 63275 199075 63278
rect 199377 63275 199443 63278
rect 259453 63275 259519 63278
rect 155534 63140 155540 63204
rect 155604 63202 155610 63204
rect 189165 63202 189231 63205
rect 292573 63202 292639 63205
rect 155604 63200 292639 63202
rect 155604 63144 189170 63200
rect 189226 63144 292578 63200
rect 292634 63144 292639 63200
rect 155604 63142 292639 63144
rect 155604 63140 155610 63142
rect 189165 63139 189231 63142
rect 292573 63139 292639 63142
rect 145414 63004 145420 63068
rect 145484 63066 145490 63068
rect 152457 63066 152523 63069
rect 145484 63064 152523 63066
rect 145484 63008 152462 63064
rect 152518 63008 152523 63064
rect 145484 63006 152523 63008
rect 145484 63004 145490 63006
rect 152457 63003 152523 63006
rect 172278 63004 172284 63068
rect 172348 63066 172354 63068
rect 199377 63066 199443 63069
rect 414657 63066 414723 63069
rect 172348 63006 180810 63066
rect 172348 63004 172354 63006
rect 180750 62930 180810 63006
rect 199377 63064 414723 63066
rect 199377 63008 199382 63064
rect 199438 63008 414662 63064
rect 414718 63008 414723 63064
rect 199377 63006 414723 63008
rect 199377 63003 199443 63006
rect 414657 63003 414723 63006
rect 197854 62930 197860 62932
rect 180750 62870 197860 62930
rect 197854 62868 197860 62870
rect 197924 62930 197930 62932
rect 514017 62930 514083 62933
rect 197924 62928 514083 62930
rect 197924 62872 514022 62928
rect 514078 62872 514083 62928
rect 197924 62870 514083 62872
rect 197924 62868 197930 62870
rect 514017 62867 514083 62870
rect 175958 62732 175964 62796
rect 176028 62794 176034 62796
rect 198774 62794 198780 62796
rect 176028 62734 198780 62794
rect 176028 62732 176034 62734
rect 198774 62732 198780 62734
rect 198844 62794 198850 62796
rect 567837 62794 567903 62797
rect 198844 62792 567903 62794
rect 198844 62736 567842 62792
rect 567898 62736 567903 62792
rect 198844 62734 567903 62736
rect 198844 62732 198850 62734
rect 567837 62731 567903 62734
rect 166206 62052 166212 62116
rect 166276 62114 166282 62116
rect 200481 62114 200547 62117
rect 201401 62114 201467 62117
rect 166276 62112 201467 62114
rect 166276 62056 200486 62112
rect 200542 62056 201406 62112
rect 201462 62056 201467 62112
rect 166276 62054 201467 62056
rect 166276 62052 166282 62054
rect 200481 62051 200547 62054
rect 201401 62051 201467 62054
rect 151486 61916 151492 61980
rect 151556 61978 151562 61980
rect 180558 61978 180564 61980
rect 151556 61918 180564 61978
rect 151556 61916 151562 61918
rect 180558 61916 180564 61918
rect 180628 61978 180634 61980
rect 245653 61978 245719 61981
rect 180628 61976 245719 61978
rect 180628 61920 245658 61976
rect 245714 61920 245719 61976
rect 180628 61918 245719 61920
rect 180628 61916 180634 61918
rect 245653 61915 245719 61918
rect 154246 61780 154252 61844
rect 154316 61842 154322 61844
rect 187785 61842 187851 61845
rect 277393 61842 277459 61845
rect 154316 61840 277459 61842
rect 154316 61784 187790 61840
rect 187846 61784 277398 61840
rect 277454 61784 277459 61840
rect 154316 61782 277459 61784
rect 154316 61780 154322 61782
rect 187785 61779 187851 61782
rect 277393 61779 277459 61782
rect 156638 61644 156644 61708
rect 156708 61706 156714 61708
rect 190729 61706 190795 61709
rect 309133 61706 309199 61709
rect 156708 61704 309199 61706
rect 156708 61648 190734 61704
rect 190790 61648 309138 61704
rect 309194 61648 309199 61704
rect 156708 61646 309199 61648
rect 156708 61644 156714 61646
rect 190729 61643 190795 61646
rect 309133 61643 309199 61646
rect 176142 61508 176148 61572
rect 176212 61570 176218 61572
rect 197302 61570 197308 61572
rect 176212 61510 197308 61570
rect 176212 61508 176218 61510
rect 197302 61508 197308 61510
rect 197372 61570 197378 61572
rect 201401 61570 201467 61573
rect 440233 61570 440299 61573
rect 197372 61510 200130 61570
rect 197372 61508 197378 61510
rect 200070 61434 200130 61510
rect 201401 61568 440299 61570
rect 201401 61512 201406 61568
rect 201462 61512 440238 61568
rect 440294 61512 440299 61568
rect 201401 61510 440299 61512
rect 201401 61507 201467 61510
rect 440233 61507 440299 61510
rect 563697 61434 563763 61437
rect 200070 61432 563763 61434
rect 200070 61376 563702 61432
rect 563758 61376 563763 61432
rect 200070 61374 563763 61376
rect 563697 61371 563763 61374
rect 152958 60556 152964 60620
rect 153028 60618 153034 60620
rect 186865 60618 186931 60621
rect 153028 60616 200130 60618
rect 153028 60560 186870 60616
rect 186926 60560 200130 60616
rect 153028 60558 200130 60560
rect 153028 60556 153034 60558
rect 186865 60555 186931 60558
rect 158110 60420 158116 60484
rect 158180 60482 158186 60484
rect 191925 60482 191991 60485
rect 193121 60482 193187 60485
rect 158180 60480 193187 60482
rect 158180 60424 191930 60480
rect 191986 60424 193126 60480
rect 193182 60424 193187 60480
rect 158180 60422 193187 60424
rect 158180 60420 158186 60422
rect 191925 60419 191991 60422
rect 193121 60419 193187 60422
rect 200070 60346 200130 60558
rect 263593 60346 263659 60349
rect 200070 60344 263659 60346
rect 200070 60288 263598 60344
rect 263654 60288 263659 60344
rect 200070 60286 263659 60288
rect 263593 60283 263659 60286
rect 155718 60148 155724 60212
rect 155788 60210 155794 60212
rect 189993 60210 190059 60213
rect 299473 60210 299539 60213
rect 155788 60208 299539 60210
rect 155788 60152 189998 60208
rect 190054 60152 299478 60208
rect 299534 60152 299539 60208
rect 155788 60150 299539 60152
rect 155788 60148 155794 60150
rect 189993 60147 190059 60150
rect 299473 60147 299539 60150
rect 193121 60074 193187 60077
rect 338113 60074 338179 60077
rect 193121 60072 338179 60074
rect 193121 60016 193126 60072
rect 193182 60016 338118 60072
rect 338174 60016 338179 60072
rect 193121 60014 338179 60016
rect 193121 60011 193187 60014
rect 338113 60011 338179 60014
rect 173566 59876 173572 59940
rect 173636 59938 173642 59940
rect 200389 59938 200455 59941
rect 525057 59938 525123 59941
rect 173636 59936 525123 59938
rect 173636 59880 200394 59936
rect 200450 59880 525062 59936
rect 525118 59880 525123 59936
rect 173636 59878 525123 59880
rect 173636 59876 173642 59878
rect 200389 59875 200455 59878
rect 525057 59875 525123 59878
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect 104801 59258 104867 59261
rect 135662 59258 135668 59260
rect 104801 59256 135668 59258
rect 104801 59200 104806 59256
rect 104862 59200 135668 59256
rect 104801 59198 135668 59200
rect 104801 59195 104867 59198
rect 135662 59196 135668 59198
rect 135732 59196 135738 59260
rect 160686 59196 160692 59260
rect 160756 59258 160762 59260
rect 194777 59258 194843 59261
rect 195053 59258 195119 59261
rect 160756 59256 195119 59258
rect 160756 59200 194782 59256
rect 194838 59200 195058 59256
rect 195114 59200 195119 59256
rect 160756 59198 195119 59200
rect 160756 59196 160762 59198
rect 194777 59195 194843 59198
rect 195053 59195 195119 59198
rect 154062 59060 154068 59124
rect 154132 59122 154138 59124
rect 187785 59122 187851 59125
rect 154132 59120 187851 59122
rect 154132 59064 187790 59120
rect 187846 59064 187851 59120
rect 154132 59062 187851 59064
rect 154132 59060 154138 59062
rect 187785 59059 187851 59062
rect 151670 58924 151676 58988
rect 151740 58986 151746 58988
rect 183686 58986 183692 58988
rect 151740 58926 183692 58986
rect 151740 58924 151746 58926
rect 183686 58924 183692 58926
rect 183756 58986 183762 58988
rect 249793 58986 249859 58989
rect 183756 58984 249859 58986
rect 183756 58928 249798 58984
rect 249854 58928 249859 58984
rect 183756 58926 249859 58928
rect 183756 58924 183762 58926
rect 249793 58923 249859 58926
rect 187785 58850 187851 58853
rect 188337 58850 188403 58853
rect 281533 58850 281599 58853
rect 187785 58848 281599 58850
rect 187785 58792 187790 58848
rect 187846 58792 188342 58848
rect 188398 58792 281538 58848
rect 281594 58792 281599 58848
rect 187785 58790 281599 58792
rect 187785 58787 187851 58790
rect 188337 58787 188403 58790
rect 281533 58787 281599 58790
rect -960 58578 480 58668
rect 158294 58652 158300 58716
rect 158364 58714 158370 58716
rect 191833 58714 191899 58717
rect 331213 58714 331279 58717
rect 158364 58712 331279 58714
rect 158364 58656 191838 58712
rect 191894 58656 331218 58712
rect 331274 58656 331279 58712
rect 158364 58654 331279 58656
rect 158364 58652 158370 58654
rect 191833 58651 191899 58654
rect 331213 58651 331279 58654
rect 49693 58578 49759 58581
rect 104065 58578 104131 58581
rect 104801 58578 104867 58581
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect 49693 58576 104867 58578
rect 49693 58520 49698 58576
rect 49754 58520 104070 58576
rect 104126 58520 104806 58576
rect 104862 58520 104867 58576
rect 49693 58518 104867 58520
rect 49693 58515 49759 58518
rect 104065 58515 104131 58518
rect 104801 58515 104867 58518
rect 195053 58578 195119 58581
rect 362953 58578 363019 58581
rect 195053 58576 363019 58578
rect 195053 58520 195058 58576
rect 195114 58520 362958 58576
rect 363014 58520 363019 58576
rect 195053 58518 363019 58520
rect 195053 58515 195119 58518
rect 362953 58515 363019 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 122046 58034 122052 58036
rect 246 57974 122052 58034
rect 122046 57972 122052 57974
rect 122116 57972 122122 58036
rect 100753 57898 100819 57901
rect 101673 57898 101739 57901
rect 134006 57898 134012 57900
rect 100753 57896 134012 57898
rect 100753 57840 100758 57896
rect 100814 57840 101678 57896
rect 101734 57840 134012 57896
rect 100753 57838 134012 57840
rect 100753 57835 100819 57838
rect 101673 57835 101739 57838
rect 134006 57836 134012 57838
rect 134076 57836 134082 57900
rect 156822 57836 156828 57900
rect 156892 57898 156898 57900
rect 190637 57898 190703 57901
rect 156892 57896 200130 57898
rect 156892 57840 190642 57896
rect 190698 57840 200130 57896
rect 156892 57838 200130 57840
rect 156892 57836 156898 57838
rect 190637 57835 190703 57838
rect 165286 57700 165292 57764
rect 165356 57762 165362 57764
rect 165356 57702 180810 57762
rect 165356 57700 165362 57702
rect 180750 57354 180810 57702
rect 200070 57490 200130 57838
rect 313273 57490 313339 57493
rect 200070 57488 313339 57490
rect 200070 57432 313278 57488
rect 313334 57432 313339 57488
rect 200070 57430 313339 57432
rect 313273 57427 313339 57430
rect 198917 57354 198983 57357
rect 418797 57354 418863 57357
rect 180750 57352 418863 57354
rect 180750 57296 198922 57352
rect 198978 57296 418802 57352
rect 418858 57296 418863 57352
rect 180750 57294 418863 57296
rect 198917 57291 198983 57294
rect 418797 57291 418863 57294
rect 25497 57218 25563 57221
rect 100753 57218 100819 57221
rect 25497 57216 100819 57218
rect 25497 57160 25502 57216
rect 25558 57160 100758 57216
rect 100814 57160 100819 57216
rect 25497 57158 100819 57160
rect 25497 57155 25563 57158
rect 100753 57155 100819 57158
rect 174486 57156 174492 57220
rect 174556 57218 174562 57220
rect 545757 57218 545823 57221
rect 174556 57216 545823 57218
rect 174556 57160 545762 57216
rect 545818 57160 545823 57216
rect 174556 57158 545823 57160
rect 174556 57156 174562 57158
rect 545757 57155 545823 57158
rect 162342 56476 162348 56540
rect 162412 56538 162418 56540
rect 196157 56538 196223 56541
rect 200665 56540 200731 56541
rect 200614 56538 200620 56540
rect 162412 56536 196223 56538
rect 162412 56480 196162 56536
rect 196218 56480 196223 56536
rect 162412 56478 196223 56480
rect 200574 56478 200620 56538
rect 200684 56536 200731 56540
rect 200726 56480 200731 56536
rect 162412 56476 162418 56478
rect 196157 56475 196223 56478
rect 200614 56476 200620 56478
rect 200684 56476 200731 56480
rect 200665 56475 200731 56476
rect 170438 56340 170444 56404
rect 170508 56402 170514 56404
rect 203149 56402 203215 56405
rect 204161 56402 204227 56405
rect 170508 56400 204227 56402
rect 170508 56344 203154 56400
rect 203210 56344 204166 56400
rect 204222 56344 204227 56400
rect 170508 56342 204227 56344
rect 170508 56340 170514 56342
rect 203149 56339 203215 56342
rect 204161 56339 204227 56342
rect 149830 56068 149836 56132
rect 149900 56130 149906 56132
rect 231853 56130 231919 56133
rect 149900 56128 231919 56130
rect 149900 56072 231858 56128
rect 231914 56072 231919 56128
rect 149900 56070 231919 56072
rect 149900 56068 149906 56070
rect 231853 56067 231919 56070
rect 196157 55994 196223 55997
rect 382917 55994 382983 55997
rect 196157 55992 382983 55994
rect 196157 55936 196162 55992
rect 196218 55936 382922 55992
rect 382978 55936 382983 55992
rect 196157 55934 382983 55936
rect 196157 55931 196223 55934
rect 382917 55931 382983 55934
rect 146886 55796 146892 55860
rect 146956 55858 146962 55860
rect 193305 55858 193371 55861
rect 146956 55856 193371 55858
rect 146956 55800 193310 55856
rect 193366 55800 193371 55856
rect 146956 55798 193371 55800
rect 146956 55796 146962 55798
rect 193305 55795 193371 55798
rect 204161 55858 204227 55861
rect 481633 55858 481699 55861
rect 204161 55856 481699 55858
rect 204161 55800 204166 55856
rect 204222 55800 481638 55856
rect 481694 55800 481699 55856
rect 204161 55798 481699 55800
rect 204161 55795 204227 55798
rect 481633 55795 481699 55798
rect 160870 55116 160876 55180
rect 160940 55178 160946 55180
rect 194685 55178 194751 55181
rect 160940 55176 200130 55178
rect 160940 55120 194690 55176
rect 194746 55120 200130 55176
rect 160940 55118 200130 55120
rect 160940 55116 160946 55118
rect 194685 55115 194751 55118
rect 165470 54980 165476 55044
rect 165540 55042 165546 55044
rect 198825 55042 198891 55045
rect 165540 55040 198891 55042
rect 165540 54984 198830 55040
rect 198886 54984 198891 55040
rect 165540 54982 198891 54984
rect 165540 54980 165546 54982
rect 198825 54979 198891 54982
rect 200070 54634 200130 55118
rect 364977 54634 365043 54637
rect 200070 54632 365043 54634
rect 200070 54576 364982 54632
rect 365038 54576 365043 54632
rect 200070 54574 365043 54576
rect 364977 54571 365043 54574
rect 198825 54498 198891 54501
rect 423765 54498 423831 54501
rect 198825 54496 423831 54498
rect 198825 54440 198830 54496
rect 198886 54440 423770 54496
rect 423826 54440 423831 54496
rect 198825 54438 423831 54440
rect 198825 54435 198891 54438
rect 423765 54435 423831 54438
rect 107561 53818 107627 53821
rect 139342 53818 139348 53820
rect 107561 53816 139348 53818
rect 107561 53760 107566 53816
rect 107622 53760 139348 53816
rect 107561 53758 139348 53760
rect 107561 53755 107627 53758
rect 139342 53756 139348 53758
rect 139412 53756 139418 53820
rect 157006 53756 157012 53820
rect 157076 53818 157082 53820
rect 190545 53818 190611 53821
rect 157076 53816 200130 53818
rect 157076 53760 190550 53816
rect 190606 53760 200130 53816
rect 157076 53758 200130 53760
rect 157076 53756 157082 53758
rect 190545 53755 190611 53758
rect 162526 53620 162532 53684
rect 162596 53682 162602 53684
rect 196065 53682 196131 53685
rect 162596 53680 196131 53682
rect 162596 53624 196070 53680
rect 196126 53624 196131 53680
rect 162596 53622 196131 53624
rect 162596 53620 162602 53622
rect 196065 53619 196131 53622
rect 158846 53484 158852 53548
rect 158916 53546 158922 53548
rect 189349 53546 189415 53549
rect 200070 53546 200130 53758
rect 320173 53546 320239 53549
rect 158916 53544 190470 53546
rect 158916 53488 189354 53544
rect 189410 53488 190470 53544
rect 158916 53486 190470 53488
rect 200070 53544 320239 53546
rect 200070 53488 320178 53544
rect 320234 53488 320239 53544
rect 200070 53486 320239 53488
rect 158916 53484 158922 53486
rect 189349 53483 189415 53486
rect 190410 53410 190470 53486
rect 320173 53483 320239 53486
rect 351913 53410 351979 53413
rect 190410 53408 351979 53410
rect 190410 53352 351918 53408
rect 351974 53352 351979 53408
rect 190410 53350 351979 53352
rect 351913 53347 351979 53350
rect 166390 53212 166396 53276
rect 166460 53274 166466 53276
rect 196065 53274 196131 53277
rect 387793 53274 387859 53277
rect 166460 53214 180810 53274
rect 166460 53212 166466 53214
rect 102133 53138 102199 53141
rect 107561 53138 107627 53141
rect 102133 53136 107627 53138
rect 102133 53080 102138 53136
rect 102194 53080 107566 53136
rect 107622 53080 107627 53136
rect 102133 53078 107627 53080
rect 180750 53138 180810 53214
rect 196065 53272 387859 53274
rect 196065 53216 196070 53272
rect 196126 53216 387798 53272
rect 387854 53216 387859 53272
rect 196065 53214 387859 53216
rect 196065 53211 196131 53214
rect 387793 53211 387859 53214
rect 190821 53138 190887 53141
rect 433333 53138 433399 53141
rect 180750 53136 433399 53138
rect 180750 53080 190826 53136
rect 190882 53080 433338 53136
rect 433394 53080 433399 53136
rect 180750 53078 433399 53080
rect 102133 53075 102199 53078
rect 107561 53075 107627 53078
rect 190821 53075 190887 53078
rect 433333 53075 433399 53078
rect 100753 52458 100819 52461
rect 101765 52458 101831 52461
rect 133822 52458 133828 52460
rect 100753 52456 133828 52458
rect 100753 52400 100758 52456
rect 100814 52400 101770 52456
rect 101826 52400 133828 52456
rect 100753 52398 133828 52400
rect 100753 52395 100819 52398
rect 101765 52395 101831 52398
rect 133822 52396 133828 52398
rect 133892 52396 133898 52460
rect 163262 52396 163268 52460
rect 163332 52458 163338 52460
rect 197537 52458 197603 52461
rect 197997 52458 198063 52461
rect 163332 52456 198063 52458
rect 163332 52400 197542 52456
rect 197598 52400 198002 52456
rect 198058 52400 198063 52456
rect 163332 52398 198063 52400
rect 163332 52396 163338 52398
rect 197537 52395 197603 52398
rect 197997 52395 198063 52398
rect 161238 52260 161244 52324
rect 161308 52322 161314 52324
rect 194593 52322 194659 52325
rect 161308 52320 194659 52322
rect 161308 52264 194598 52320
rect 194654 52264 194659 52320
rect 161308 52262 194659 52264
rect 161308 52260 161314 52262
rect 194593 52259 194659 52262
rect 161054 52124 161060 52188
rect 161124 52186 161130 52188
rect 188061 52186 188127 52189
rect 161124 52184 190470 52186
rect 161124 52128 188066 52184
rect 188122 52128 190470 52184
rect 161124 52126 190470 52128
rect 161124 52124 161130 52126
rect 188061 52123 188127 52126
rect 190410 51914 190470 52126
rect 194593 52050 194659 52053
rect 369853 52050 369919 52053
rect 194593 52048 369919 52050
rect 194593 51992 194598 52048
rect 194654 51992 369858 52048
rect 369914 51992 369919 52048
rect 194593 51990 369919 51992
rect 194593 51987 194659 51990
rect 369853 51987 369919 51990
rect 374085 51914 374151 51917
rect 190410 51912 374151 51914
rect 190410 51856 374090 51912
rect 374146 51856 374151 51912
rect 190410 51854 374151 51856
rect 374085 51851 374151 51854
rect 27705 51778 27771 51781
rect 100753 51778 100819 51781
rect 27705 51776 100819 51778
rect 27705 51720 27710 51776
rect 27766 51720 100758 51776
rect 100814 51720 100819 51776
rect 27705 51718 100819 51720
rect 27705 51715 27771 51718
rect 100753 51715 100819 51718
rect 197997 51778 198063 51781
rect 400949 51778 401015 51781
rect 197997 51776 401015 51778
rect 197997 51720 198002 51776
rect 198058 51720 400954 51776
rect 401010 51720 401015 51776
rect 197997 51718 401015 51720
rect 197997 51715 198063 51718
rect 400949 51715 401015 51718
rect 166574 50900 166580 50964
rect 166644 50962 166650 50964
rect 200205 50962 200271 50965
rect 201401 50962 201467 50965
rect 166644 50960 201467 50962
rect 166644 50904 200210 50960
rect 200266 50904 201406 50960
rect 201462 50904 201467 50960
rect 166644 50902 201467 50904
rect 166644 50900 166650 50902
rect 200205 50899 200271 50902
rect 201401 50899 201467 50902
rect 162710 50764 162716 50828
rect 162780 50826 162786 50828
rect 195973 50826 196039 50829
rect 196433 50826 196499 50829
rect 162780 50824 196499 50826
rect 162780 50768 195978 50824
rect 196034 50768 196438 50824
rect 196494 50768 196499 50824
rect 162780 50766 196499 50768
rect 162780 50764 162786 50766
rect 195973 50763 196039 50766
rect 196433 50763 196499 50766
rect 159030 50628 159036 50692
rect 159100 50690 159106 50692
rect 187969 50690 188035 50693
rect 356053 50690 356119 50693
rect 159100 50688 356119 50690
rect 159100 50632 187974 50688
rect 188030 50632 356058 50688
rect 356114 50632 356119 50688
rect 159100 50630 356119 50632
rect 159100 50628 159106 50630
rect 187969 50627 188035 50630
rect 356053 50627 356119 50630
rect 196433 50554 196499 50557
rect 390553 50554 390619 50557
rect 196433 50552 390619 50554
rect 196433 50496 196438 50552
rect 196494 50496 390558 50552
rect 390614 50496 390619 50552
rect 196433 50494 390619 50496
rect 196433 50491 196499 50494
rect 390553 50491 390619 50494
rect 201401 50418 201467 50421
rect 437473 50418 437539 50421
rect 201401 50416 437539 50418
rect 201401 50360 201406 50416
rect 201462 50360 437478 50416
rect 437534 50360 437539 50416
rect 201401 50358 437539 50360
rect 201401 50355 201467 50358
rect 437473 50355 437539 50358
rect 177062 50220 177068 50284
rect 177132 50282 177138 50284
rect 204713 50282 204779 50285
rect 569953 50282 570019 50285
rect 177132 50280 570019 50282
rect 177132 50224 204718 50280
rect 204774 50224 569958 50280
rect 570014 50224 570019 50280
rect 177132 50222 570019 50224
rect 177132 50220 177138 50222
rect 204713 50219 204779 50222
rect 569953 50219 570019 50222
rect 100753 49602 100819 49605
rect 101949 49602 102015 49605
rect 135478 49602 135484 49604
rect 100753 49600 135484 49602
rect 100753 49544 100758 49600
rect 100814 49544 101954 49600
rect 102010 49544 135484 49600
rect 100753 49542 135484 49544
rect 100753 49539 100819 49542
rect 101949 49539 102015 49542
rect 135478 49540 135484 49542
rect 135548 49540 135554 49604
rect 167494 49540 167500 49604
rect 167564 49602 167570 49604
rect 201769 49602 201835 49605
rect 202781 49602 202847 49605
rect 167564 49600 202847 49602
rect 167564 49544 201774 49600
rect 201830 49544 202786 49600
rect 202842 49544 202847 49600
rect 167564 49542 202847 49544
rect 167564 49540 167570 49542
rect 201769 49539 201835 49542
rect 202781 49539 202847 49542
rect 163446 49404 163452 49468
rect 163516 49466 163522 49468
rect 197353 49466 197419 49469
rect 198457 49466 198523 49469
rect 163516 49464 198523 49466
rect 163516 49408 197358 49464
rect 197414 49408 198462 49464
rect 198518 49408 198523 49464
rect 163516 49406 198523 49408
rect 163516 49404 163522 49406
rect 197353 49403 197419 49406
rect 198457 49403 198523 49406
rect 169334 49268 169340 49332
rect 169404 49330 169410 49332
rect 202965 49330 203031 49333
rect 204161 49330 204227 49333
rect 169404 49328 204227 49330
rect 169404 49272 202970 49328
rect 203026 49272 204166 49328
rect 204222 49272 204227 49328
rect 169404 49270 204227 49272
rect 169404 49268 169410 49270
rect 202965 49267 203031 49270
rect 204161 49267 204227 49270
rect 198457 49194 198523 49197
rect 405733 49194 405799 49197
rect 198457 49192 405799 49194
rect 198457 49136 198462 49192
rect 198518 49136 405738 49192
rect 405794 49136 405799 49192
rect 198457 49134 405799 49136
rect 198457 49131 198523 49134
rect 405733 49131 405799 49134
rect 202781 49058 202847 49061
rect 455413 49058 455479 49061
rect 202781 49056 455479 49058
rect 202781 49000 202786 49056
rect 202842 49000 455418 49056
rect 455474 49000 455479 49056
rect 202781 48998 455479 49000
rect 202781 48995 202847 48998
rect 455413 48995 455479 48998
rect 39297 48922 39363 48925
rect 100753 48922 100819 48925
rect 39297 48920 100819 48922
rect 39297 48864 39302 48920
rect 39358 48864 100758 48920
rect 100814 48864 100819 48920
rect 39297 48862 100819 48864
rect 39297 48859 39363 48862
rect 100753 48859 100819 48862
rect 204161 48922 204227 48925
rect 466453 48922 466519 48925
rect 204161 48920 466519 48922
rect 204161 48864 204166 48920
rect 204222 48864 466458 48920
rect 466514 48864 466519 48920
rect 204161 48862 466519 48864
rect 204161 48859 204227 48862
rect 466453 48859 466519 48862
rect 100753 48242 100819 48245
rect 102041 48242 102107 48245
rect 135294 48242 135300 48244
rect 100753 48240 135300 48242
rect 100753 48184 100758 48240
rect 100814 48184 102046 48240
rect 102102 48184 135300 48240
rect 100753 48182 135300 48184
rect 100753 48179 100819 48182
rect 102041 48179 102107 48182
rect 135294 48180 135300 48182
rect 135364 48180 135370 48244
rect 166758 48180 166764 48244
rect 166828 48242 166834 48244
rect 200297 48242 200363 48245
rect 201401 48242 201467 48245
rect 166828 48240 201467 48242
rect 166828 48184 200302 48240
rect 200358 48184 201406 48240
rect 201462 48184 201467 48240
rect 166828 48182 201467 48184
rect 166828 48180 166834 48182
rect 200297 48179 200363 48182
rect 201401 48179 201467 48182
rect 163630 48044 163636 48108
rect 163700 48106 163706 48108
rect 193213 48106 193279 48109
rect 194501 48106 194567 48109
rect 163700 48104 194567 48106
rect 163700 48048 193218 48104
rect 193274 48048 194506 48104
rect 194562 48048 194567 48104
rect 163700 48046 194567 48048
rect 163700 48044 163706 48046
rect 193213 48043 193279 48046
rect 194501 48043 194567 48046
rect 173750 47908 173756 47972
rect 173820 47970 173826 47972
rect 203006 47970 203012 47972
rect 173820 47910 203012 47970
rect 173820 47908 173826 47910
rect 203006 47908 203012 47910
rect 203076 47970 203082 47972
rect 204110 47970 204116 47972
rect 203076 47910 204116 47970
rect 203076 47908 203082 47910
rect 204110 47908 204116 47910
rect 204180 47908 204186 47972
rect 194501 47834 194567 47837
rect 408493 47834 408559 47837
rect 194501 47832 408559 47834
rect 194501 47776 194506 47832
rect 194562 47776 408498 47832
rect 408554 47776 408559 47832
rect 194501 47774 408559 47776
rect 194501 47771 194567 47774
rect 408493 47771 408559 47774
rect 201401 47698 201467 47701
rect 444373 47698 444439 47701
rect 201401 47696 444439 47698
rect 201401 47640 201406 47696
rect 201462 47640 444378 47696
rect 444434 47640 444439 47696
rect 201401 47638 444439 47640
rect 201401 47635 201467 47638
rect 444373 47635 444439 47638
rect 44173 47562 44239 47565
rect 100753 47562 100819 47565
rect 44173 47560 100819 47562
rect 44173 47504 44178 47560
rect 44234 47504 100758 47560
rect 100814 47504 100819 47560
rect 44173 47502 100819 47504
rect 44173 47499 44239 47502
rect 100753 47499 100819 47502
rect 204110 47500 204116 47564
rect 204180 47562 204186 47564
rect 520917 47562 520983 47565
rect 204180 47560 520983 47562
rect 204180 47504 520922 47560
rect 520978 47504 520983 47560
rect 204180 47502 520983 47504
rect 204180 47500 204186 47502
rect 520917 47499 520983 47502
rect 102225 46882 102291 46885
rect 102685 46882 102751 46885
rect 136582 46882 136588 46884
rect 102225 46880 136588 46882
rect 102225 46824 102230 46880
rect 102286 46824 102690 46880
rect 102746 46824 136588 46880
rect 102225 46822 136588 46824
rect 102225 46819 102291 46822
rect 102685 46819 102751 46822
rect 136582 46820 136588 46822
rect 136652 46820 136658 46884
rect 167678 46820 167684 46884
rect 167748 46882 167754 46884
rect 201677 46882 201743 46885
rect 202781 46882 202847 46885
rect 167748 46880 202847 46882
rect 167748 46824 201682 46880
rect 201738 46824 202786 46880
rect 202842 46824 202847 46880
rect 167748 46822 202847 46824
rect 167748 46820 167754 46822
rect 201677 46819 201743 46822
rect 202781 46819 202847 46822
rect 148174 46276 148180 46340
rect 148244 46338 148250 46340
rect 208393 46338 208459 46341
rect 583520 46338 584960 46428
rect 148244 46336 208459 46338
rect 148244 46280 208398 46336
rect 208454 46280 208459 46336
rect 148244 46278 208459 46280
rect 148244 46276 148250 46278
rect 208393 46275 208459 46278
rect 583342 46278 584960 46338
rect 56593 46202 56659 46205
rect 102225 46202 102291 46205
rect 56593 46200 102291 46202
rect 56593 46144 56598 46200
rect 56654 46144 102230 46200
rect 102286 46144 102291 46200
rect 56593 46142 102291 46144
rect 56593 46139 56659 46142
rect 102225 46139 102291 46142
rect 202781 46202 202847 46205
rect 462313 46202 462379 46205
rect 202781 46200 462379 46202
rect 202781 46144 202786 46200
rect 202842 46144 462318 46200
rect 462374 46144 462379 46200
rect 202781 46142 462379 46144
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect 202781 46139 202847 46142
rect 462313 46139 462379 46142
rect -960 45522 480 45612
rect 192334 45596 192340 45660
rect 192404 45658 192410 45660
rect 583526 45658 583586 46142
rect 192404 45598 583586 45658
rect 192404 45596 192410 45598
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 167862 45460 167868 45524
rect 167932 45522 167938 45524
rect 201585 45522 201651 45525
rect 167932 45520 201651 45522
rect 167932 45464 201590 45520
rect 201646 45464 201651 45520
rect 167932 45462 201651 45464
rect 167932 45460 167938 45462
rect 201585 45459 201651 45462
rect 157190 45324 157196 45388
rect 157260 45386 157266 45388
rect 190453 45386 190519 45389
rect 157260 45384 190519 45386
rect 157260 45328 190458 45384
rect 190514 45328 190519 45384
rect 157260 45326 190519 45328
rect 157260 45324 157266 45326
rect 190410 45323 190519 45326
rect 190410 45250 190470 45323
rect 315297 45250 315363 45253
rect 190410 45248 315363 45250
rect 190410 45192 315302 45248
rect 315358 45192 315363 45248
rect 190410 45190 315363 45192
rect 315297 45187 315363 45190
rect 201585 45114 201651 45117
rect 458173 45114 458239 45117
rect 201585 45112 458239 45114
rect 201585 45056 201590 45112
rect 201646 45056 458178 45112
rect 458234 45056 458239 45112
rect 201585 45054 458239 45056
rect 201585 45051 201651 45054
rect 458173 45051 458239 45054
rect 176326 44916 176332 44980
rect 176396 44978 176402 44980
rect 205633 44978 205699 44981
rect 553393 44978 553459 44981
rect 176396 44976 553459 44978
rect 176396 44920 205638 44976
rect 205694 44920 553398 44976
rect 553454 44920 553459 44976
rect 176396 44918 553459 44920
rect 176396 44916 176402 44918
rect 205633 44915 205699 44918
rect 553393 44915 553459 44918
rect 176510 44780 176516 44844
rect 176580 44842 176586 44844
rect 204529 44842 204595 44845
rect 565813 44842 565879 44845
rect 176580 44840 565879 44842
rect 176580 44784 204534 44840
rect 204590 44784 565818 44840
rect 565874 44784 565879 44840
rect 176580 44782 565879 44784
rect 176580 44780 176586 44782
rect 204529 44779 204595 44782
rect 565813 44779 565879 44782
rect 168046 44100 168052 44164
rect 168116 44162 168122 44164
rect 202321 44162 202387 44165
rect 168116 44160 202387 44162
rect 168116 44104 202326 44160
rect 202382 44104 202387 44160
rect 168116 44102 202387 44104
rect 168116 44100 168122 44102
rect 202321 44099 202387 44102
rect 169518 43964 169524 44028
rect 169588 44026 169594 44028
rect 202873 44026 202939 44029
rect 169588 44024 202939 44026
rect 169588 43968 202878 44024
rect 202934 43968 202939 44024
rect 169588 43966 202939 43968
rect 169588 43964 169594 43966
rect 202873 43963 202939 43966
rect 202321 43618 202387 43621
rect 448605 43618 448671 43621
rect 202321 43616 448671 43618
rect 202321 43560 202326 43616
rect 202382 43560 448610 43616
rect 448666 43560 448671 43616
rect 202321 43558 448671 43560
rect 202321 43555 202387 43558
rect 448605 43555 448671 43558
rect 202873 43482 202939 43485
rect 476113 43482 476179 43485
rect 202873 43480 476179 43482
rect 202873 43424 202878 43480
rect 202934 43424 476118 43480
rect 476174 43424 476179 43480
rect 202873 43422 476179 43424
rect 202873 43419 202939 43422
rect 476113 43419 476179 43422
rect 149646 42060 149652 42124
rect 149716 42122 149722 42124
rect 229093 42122 229159 42125
rect 149716 42120 229159 42122
rect 149716 42064 229098 42120
rect 229154 42064 229159 42120
rect 149716 42062 229159 42064
rect 149716 42060 149722 42062
rect 229093 42059 229159 42062
rect 17217 36546 17283 36549
rect 133638 36546 133644 36548
rect 17217 36544 133644 36546
rect 17217 36488 17222 36544
rect 17278 36488 133644 36544
rect 17217 36486 133644 36488
rect 17217 36483 17283 36486
rect 133638 36484 133644 36486
rect 133708 36484 133714 36548
rect 24853 33826 24919 33829
rect 134558 33826 134564 33828
rect 24853 33824 134564 33826
rect 24853 33768 24858 33824
rect 24914 33768 134564 33824
rect 24853 33766 134564 33768
rect 24853 33763 24919 33766
rect 134558 33764 134564 33766
rect 134628 33764 134634 33828
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31786 306 32270
rect 120758 31786 120764 31788
rect 246 31726 120764 31786
rect 120758 31724 120764 31726
rect 120828 31724 120834 31788
rect 189758 31724 189764 31788
rect 189828 31786 189834 31788
rect 583526 31786 583586 32950
rect 189828 31726 583586 31786
rect 189828 31724 189834 31726
rect 144494 30908 144500 30972
rect 144564 30970 144570 30972
rect 160093 30970 160159 30973
rect 144564 30968 160159 30970
rect 144564 30912 160098 30968
rect 160154 30912 160159 30968
rect 144564 30910 160159 30912
rect 144564 30908 144570 30910
rect 160093 30907 160159 30910
rect 151118 29548 151124 29612
rect 151188 29610 151194 29612
rect 242985 29610 243051 29613
rect 151188 29608 243051 29610
rect 151188 29552 242990 29608
rect 243046 29552 243051 29608
rect 151188 29550 243051 29552
rect 151188 29548 151194 29550
rect 242985 29547 243051 29550
rect 153694 26828 153700 26892
rect 153764 26890 153770 26892
rect 282913 26890 282979 26893
rect 153764 26888 282979 26890
rect 153764 26832 282918 26888
rect 282974 26832 282979 26888
rect 153764 26830 282979 26832
rect 153764 26828 153770 26830
rect 282913 26827 282979 26830
rect 144310 21252 144316 21316
rect 144380 21314 144386 21316
rect 157333 21314 157399 21317
rect 144380 21312 157399 21314
rect 144380 21256 157338 21312
rect 157394 21256 157399 21312
rect 144380 21254 157399 21256
rect 144380 21252 144386 21254
rect 157333 21251 157399 21254
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 145598 18532 145604 18596
rect 145668 18594 145674 18596
rect 175917 18594 175983 18597
rect 145668 18592 175983 18594
rect 145668 18536 175922 18592
rect 175978 18536 175983 18592
rect 145668 18534 175983 18536
rect 145668 18532 145674 18534
rect 175917 18531 175983 18534
rect 152406 12956 152412 13020
rect 152476 13018 152482 13020
rect 264973 13018 265039 13021
rect 152476 13016 265039 13018
rect 152476 12960 264978 13016
rect 265034 12960 265039 13016
rect 152476 12958 265039 12960
rect 152476 12956 152482 12958
rect 264973 12955 265039 12958
rect 144126 8876 144132 8940
rect 144196 8938 144202 8940
rect 161289 8938 161355 8941
rect 144196 8936 161355 8938
rect 144196 8880 161294 8936
rect 161350 8880 161355 8936
rect 144196 8878 161355 8880
rect 144196 8876 144202 8878
rect 161289 8875 161355 8878
rect 148542 7516 148548 7580
rect 148612 7578 148618 7580
rect 213361 7578 213427 7581
rect 148612 7576 213427 7578
rect 148612 7520 213366 7576
rect 213422 7520 213427 7576
rect 148612 7518 213427 7520
rect 148612 7516 148618 7518
rect 213361 7515 213427 7518
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 158478 6156 158484 6220
rect 158548 6218 158554 6220
rect 336273 6218 336339 6221
rect 158548 6216 336339 6218
rect 158548 6160 336278 6216
rect 336334 6160 336339 6216
rect 158548 6158 336339 6160
rect 158548 6156 158554 6158
rect 336273 6155 336339 6158
rect 142654 3300 142660 3364
rect 142724 3362 142730 3364
rect 171961 3362 172027 3365
rect 142724 3360 172027 3362
rect 142724 3304 171966 3360
rect 172022 3304 172027 3360
rect 142724 3302 172027 3304
rect 142724 3300 142730 3302
rect 171961 3299 172027 3302
<< via3 >>
rect 187372 284276 187436 284340
rect 189028 278020 189092 278084
rect 189028 277476 189092 277540
rect 187740 275980 187804 276044
rect 196204 265372 196268 265436
rect 193260 265236 193324 265300
rect 112852 265100 112916 265164
rect 194732 265100 194796 265164
rect 113036 264964 113100 265028
rect 197492 264964 197556 265028
rect 122604 263876 122668 263940
rect 115796 263740 115860 263804
rect 118372 263604 118436 263668
rect 116900 263196 116964 263260
rect 119844 263060 119908 263124
rect 113772 262924 113836 262988
rect 113956 262788 114020 262852
rect 118188 262652 118252 262716
rect 193444 262652 193508 262716
rect 115428 262516 115492 262580
rect 192156 262516 192220 262580
rect 114140 262380 114204 262444
rect 191972 262380 192036 262444
rect 187924 262304 187988 262308
rect 187924 262248 187974 262304
rect 187974 262248 187988 262304
rect 187924 262244 187988 262248
rect 192340 262304 192404 262308
rect 192340 262248 192354 262304
rect 192354 262248 192404 262304
rect 192340 262244 192404 262248
rect 111564 261020 111628 261084
rect 111380 260884 111444 260948
rect 193628 260884 193692 260948
rect 115612 260476 115676 260540
rect 117084 260340 117148 260404
rect 120948 260204 121012 260268
rect 118556 260068 118620 260132
rect 189396 260068 189460 260132
rect 119660 259932 119724 259996
rect 188108 259932 188172 259996
rect 122236 259796 122300 259860
rect 188292 259796 188356 259860
rect 116716 259660 116780 259724
rect 121132 259584 121196 259588
rect 121132 259528 121182 259584
rect 121182 259528 121196 259584
rect 121132 259524 121196 259528
rect 123156 259524 123220 259588
rect 124076 259524 124140 259588
rect 189580 259660 189644 259724
rect 186084 259524 186148 259588
rect 122972 259388 123036 259452
rect 186084 213828 186148 213892
rect 122788 209612 122852 209676
rect 122788 205532 122852 205596
rect 123892 200908 123956 200972
rect 153516 200908 153580 200972
rect 170996 200908 171060 200972
rect 158116 200772 158180 200836
rect 124076 200696 124140 200700
rect 124076 200640 124090 200696
rect 124090 200640 124140 200696
rect 124076 200636 124140 200640
rect 156276 200636 156340 200700
rect 173756 200636 173820 200700
rect 122972 200500 123036 200564
rect 142844 200500 142908 200564
rect 138980 200364 139044 200428
rect 132540 199820 132604 199884
rect 133092 199820 133156 199884
rect 134012 199820 134076 199884
rect 134564 199820 134628 199884
rect 135852 199820 135916 199884
rect 136220 199880 136284 199884
rect 136220 199824 136224 199880
rect 136224 199824 136280 199880
rect 136280 199824 136284 199880
rect 136220 199820 136284 199824
rect 137140 199880 137204 199884
rect 137140 199824 137144 199880
rect 137144 199824 137200 199880
rect 137200 199824 137204 199880
rect 137140 199820 137204 199824
rect 137508 199880 137572 199884
rect 137508 199824 137512 199880
rect 137512 199824 137568 199880
rect 137568 199824 137572 199880
rect 137508 199820 137572 199824
rect 137692 199820 137756 199884
rect 138428 199820 138492 199884
rect 141924 199820 141988 199884
rect 140452 199684 140516 199748
rect 142660 199820 142724 199884
rect 142844 199820 142908 199884
rect 144132 199858 144136 199884
rect 144136 199858 144192 199884
rect 144192 199858 144196 199884
rect 144132 199820 144196 199858
rect 138428 199412 138492 199476
rect 138796 199472 138860 199476
rect 138796 199416 138846 199472
rect 138846 199416 138860 199472
rect 138796 199412 138860 199416
rect 138980 199412 139044 199476
rect 146892 199684 146956 199748
rect 148916 199956 148980 200020
rect 148364 199820 148428 199884
rect 149652 199880 149716 199884
rect 149652 199824 149656 199880
rect 149656 199824 149712 199880
rect 149712 199824 149716 199880
rect 149652 199820 149716 199824
rect 150020 199880 150084 199884
rect 150020 199824 150024 199880
rect 150024 199824 150080 199880
rect 150080 199824 150084 199880
rect 150020 199820 150084 199824
rect 180748 200500 180812 200564
rect 151308 199820 151372 199884
rect 168604 200228 168668 200292
rect 161428 200092 161492 200156
rect 165660 199956 165724 200020
rect 152596 199880 152660 199884
rect 152596 199824 152600 199880
rect 152600 199824 152656 199880
rect 152656 199824 152660 199880
rect 152596 199820 152660 199824
rect 153700 199820 153764 199884
rect 154436 199820 154500 199884
rect 155540 199820 155604 199884
rect 155724 199820 155788 199884
rect 153516 199548 153580 199612
rect 153884 199548 153948 199612
rect 155724 199744 155788 199748
rect 155724 199688 155774 199744
rect 155774 199688 155788 199744
rect 155724 199684 155788 199688
rect 156828 199858 156832 199884
rect 156832 199858 156888 199884
rect 156888 199858 156892 199884
rect 156828 199820 156892 199858
rect 157932 199820 157996 199884
rect 158300 199858 158304 199884
rect 158304 199858 158360 199884
rect 158360 199858 158364 199884
rect 158300 199820 158364 199858
rect 158668 199820 158732 199884
rect 158116 199684 158180 199748
rect 159036 199684 159100 199748
rect 160876 199820 160940 199884
rect 163084 199880 163148 199884
rect 163084 199824 163088 199880
rect 163088 199824 163144 199880
rect 163144 199824 163148 199880
rect 163084 199820 163148 199824
rect 163268 199820 163332 199884
rect 164372 199880 164436 199884
rect 164372 199824 164376 199880
rect 164376 199824 164432 199880
rect 164432 199824 164436 199880
rect 164372 199820 164436 199824
rect 164556 199820 164620 199884
rect 159772 199684 159836 199748
rect 160324 199744 160388 199748
rect 160324 199688 160374 199744
rect 160374 199688 160388 199744
rect 160324 199684 160388 199688
rect 162900 199684 162964 199748
rect 163820 199684 163884 199748
rect 165844 199858 165848 199884
rect 165848 199858 165904 199884
rect 165904 199858 165908 199884
rect 165844 199820 165908 199858
rect 166580 199820 166644 199884
rect 168604 199880 168668 199884
rect 168604 199824 168608 199880
rect 168608 199824 168664 199880
rect 168664 199824 168668 199880
rect 168604 199820 168668 199824
rect 168788 199820 168852 199884
rect 166764 199744 166828 199748
rect 166764 199688 166814 199744
rect 166814 199688 166828 199744
rect 166764 199684 166828 199688
rect 167868 199684 167932 199748
rect 169156 199684 169220 199748
rect 169524 199548 169588 199612
rect 169892 200092 169956 200156
rect 170812 199956 170876 200020
rect 178356 199956 178420 200020
rect 170444 199880 170508 199884
rect 170444 199824 170448 199880
rect 170448 199824 170504 199880
rect 170504 199824 170508 199880
rect 170444 199820 170508 199824
rect 170076 199684 170140 199748
rect 171364 199858 171368 199884
rect 171368 199858 171424 199884
rect 171424 199858 171428 199884
rect 171364 199820 171428 199858
rect 171916 199820 171980 199884
rect 172100 199820 172164 199884
rect 172652 199820 172716 199884
rect 170812 199744 170876 199748
rect 170812 199688 170826 199744
rect 170826 199688 170876 199744
rect 170812 199684 170876 199688
rect 170996 199744 171060 199748
rect 170996 199688 171046 199744
rect 171046 199688 171060 199744
rect 170996 199684 171060 199688
rect 172284 199744 172348 199748
rect 172284 199688 172334 199744
rect 172334 199688 172348 199744
rect 172284 199684 172348 199688
rect 174492 199820 174556 199884
rect 176148 199820 176212 199884
rect 174492 199684 174556 199748
rect 175596 199684 175660 199748
rect 200620 199684 200684 199748
rect 180932 199548 180996 199612
rect 154620 199472 154684 199476
rect 154620 199416 154670 199472
rect 154670 199416 154684 199472
rect 154620 199412 154684 199416
rect 156276 199412 156340 199476
rect 156460 199412 156524 199476
rect 158852 199412 158916 199476
rect 161428 199412 161492 199476
rect 162900 199472 162964 199476
rect 162900 199416 162950 199472
rect 162950 199416 162964 199472
rect 162900 199412 162964 199416
rect 163268 199472 163332 199476
rect 163268 199416 163282 199472
rect 163282 199416 163332 199472
rect 163268 199412 163332 199416
rect 169892 199412 169956 199476
rect 170444 199472 170508 199476
rect 170444 199416 170458 199472
rect 170458 199416 170508 199472
rect 170444 199412 170508 199416
rect 170996 199412 171060 199476
rect 171364 199412 171428 199476
rect 173756 199472 173820 199476
rect 173756 199416 173806 199472
rect 173806 199416 173820 199472
rect 173756 199412 173820 199416
rect 133092 199336 133156 199340
rect 133092 199280 133142 199336
rect 133142 199280 133156 199336
rect 133092 199276 133156 199280
rect 139164 199276 139228 199340
rect 137508 198868 137572 198932
rect 140636 199336 140700 199340
rect 140636 199280 140650 199336
rect 140650 199280 140700 199336
rect 140636 199276 140700 199280
rect 141924 199276 141988 199340
rect 156828 199336 156892 199340
rect 156828 199280 156878 199336
rect 156878 199280 156892 199336
rect 156828 199276 156892 199280
rect 182588 199276 182652 199340
rect 140452 199140 140516 199204
rect 183508 199140 183572 199204
rect 178172 199004 178236 199068
rect 148180 198732 148244 198796
rect 183692 198868 183756 198932
rect 155908 198792 155972 198796
rect 155908 198736 155958 198792
rect 155958 198736 155972 198792
rect 155908 198732 155972 198736
rect 184980 198732 185044 198796
rect 167500 198596 167564 198660
rect 171732 198596 171796 198660
rect 171916 198596 171980 198660
rect 189212 198596 189276 198660
rect 196572 198596 196636 198660
rect 133644 198520 133708 198524
rect 133644 198464 133658 198520
rect 133658 198464 133708 198520
rect 133644 198460 133708 198464
rect 153700 198460 153764 198524
rect 187004 198460 187068 198524
rect 126836 198324 126900 198388
rect 156276 198324 156340 198388
rect 159772 198324 159836 198388
rect 190500 198324 190564 198388
rect 125364 198052 125428 198116
rect 163636 198248 163700 198252
rect 163636 198192 163650 198248
rect 163650 198192 163700 198248
rect 163636 198188 163700 198192
rect 126652 197916 126716 197980
rect 169524 198052 169588 198116
rect 171916 198112 171980 198116
rect 171916 198056 171930 198112
rect 171930 198056 171980 198112
rect 171916 198052 171980 198056
rect 174124 198052 174188 198116
rect 194548 198188 194612 198252
rect 145604 197644 145668 197708
rect 179460 197780 179524 197844
rect 179644 197508 179708 197572
rect 133460 197372 133524 197436
rect 134196 197372 134260 197436
rect 140084 197432 140148 197436
rect 140084 197376 140098 197432
rect 140098 197376 140148 197432
rect 140084 197372 140148 197376
rect 156644 197432 156708 197436
rect 156644 197376 156658 197432
rect 156658 197376 156708 197432
rect 156644 197372 156708 197376
rect 154068 197236 154132 197300
rect 166028 197236 166092 197300
rect 165844 197100 165908 197164
rect 161244 196964 161308 197028
rect 197308 196964 197372 197028
rect 163084 196828 163148 196892
rect 174676 196480 174740 196484
rect 174676 196424 174690 196480
rect 174690 196424 174740 196480
rect 174676 196420 174740 196424
rect 135852 196284 135916 196348
rect 135852 196148 135916 196212
rect 122788 196012 122852 196076
rect 136220 196072 136284 196076
rect 136220 196016 136270 196072
rect 136270 196016 136284 196072
rect 136220 196012 136284 196016
rect 139164 196072 139228 196076
rect 139164 196016 139214 196072
rect 139214 196016 139228 196072
rect 139164 196012 139228 196016
rect 158668 196012 158732 196076
rect 151492 195936 151556 195940
rect 151492 195880 151542 195936
rect 151542 195880 151556 195936
rect 151492 195876 151556 195880
rect 156092 195876 156156 195940
rect 160324 195936 160388 195940
rect 160324 195880 160338 195936
rect 160338 195880 160388 195936
rect 160324 195876 160388 195880
rect 162716 195876 162780 195940
rect 131988 195740 132052 195804
rect 128124 195604 128188 195668
rect 187188 195604 187252 195668
rect 127940 195468 128004 195532
rect 149652 195528 149716 195532
rect 149652 195472 149702 195528
rect 149702 195472 149716 195528
rect 149652 195468 149716 195472
rect 150020 195528 150084 195532
rect 150020 195472 150034 195528
rect 150034 195472 150084 195528
rect 150020 195468 150084 195472
rect 153884 195468 153948 195532
rect 168052 195468 168116 195532
rect 169156 195468 169220 195532
rect 172100 195468 172164 195532
rect 191788 195468 191852 195532
rect 145236 195332 145300 195396
rect 167684 195332 167748 195396
rect 121316 195196 121380 195260
rect 132172 195196 132236 195260
rect 148916 195196 148980 195260
rect 151124 195196 151188 195260
rect 153516 195196 153580 195260
rect 154436 195196 154500 195260
rect 162900 195196 162964 195260
rect 164740 195256 164804 195260
rect 164740 195200 164754 195256
rect 164754 195200 164804 195256
rect 164740 195196 164804 195200
rect 166580 195196 166644 195260
rect 130884 195060 130948 195124
rect 149652 195060 149716 195124
rect 152596 195060 152660 195124
rect 164372 195060 164436 195124
rect 136220 194924 136284 194988
rect 137140 194984 137204 194988
rect 137140 194928 137190 194984
rect 137190 194928 137204 194984
rect 137140 194924 137204 194928
rect 138060 194924 138124 194988
rect 139164 194984 139228 194988
rect 139164 194928 139178 194984
rect 139178 194928 139228 194984
rect 139164 194924 139228 194928
rect 148732 194924 148796 194988
rect 164556 194984 164620 194988
rect 164556 194928 164570 194984
rect 164570 194928 164620 194984
rect 164556 194924 164620 194928
rect 165660 194924 165724 194988
rect 138428 194788 138492 194852
rect 175412 194788 175476 194852
rect 187372 194788 187436 194852
rect 152228 194168 152292 194172
rect 152228 194112 152278 194168
rect 152278 194112 152292 194168
rect 152228 194108 152292 194112
rect 124996 193972 125060 194036
rect 158484 193972 158548 194036
rect 133276 193836 133340 193900
rect 151860 191524 151924 191588
rect 148916 191388 148980 191452
rect 149468 191252 149532 191316
rect 173388 191252 173452 191316
rect 141004 191116 141068 191180
rect 145420 191116 145484 191180
rect 147076 191116 147140 191180
rect 156092 191116 156156 191180
rect 158116 191116 158180 191180
rect 161060 191116 161124 191180
rect 162164 191116 162228 191180
rect 165844 191116 165908 191180
rect 169340 191176 169404 191180
rect 169340 191120 169354 191176
rect 169354 191120 169404 191176
rect 169340 191116 169404 191120
rect 171548 191116 171612 191180
rect 173020 191176 173084 191180
rect 173020 191120 173034 191176
rect 173034 191120 173084 191176
rect 173020 191116 173084 191120
rect 175780 191116 175844 191180
rect 142476 190980 142540 191044
rect 150020 190980 150084 191044
rect 160876 190980 160940 191044
rect 172836 190980 172900 191044
rect 122788 190436 122852 190500
rect 122788 190300 122852 190364
rect 140820 190300 140884 190364
rect 166212 190028 166276 190092
rect 155724 189892 155788 189956
rect 157012 189212 157076 189276
rect 170812 189212 170876 189276
rect 134380 189076 134444 189140
rect 138428 188804 138492 188868
rect 143580 188804 143644 188868
rect 152596 188864 152660 188868
rect 152596 188808 152610 188864
rect 152610 188808 152660 188864
rect 152596 188804 152660 188808
rect 138796 188532 138860 188596
rect 140452 188532 140516 188596
rect 165108 188532 165172 188596
rect 131620 188396 131684 188460
rect 136036 188396 136100 188460
rect 136588 188396 136652 188460
rect 137508 188396 137572 188460
rect 138428 188396 138492 188460
rect 140268 188396 140332 188460
rect 149836 188396 149900 188460
rect 176516 188396 176580 188460
rect 176884 188396 176948 188460
rect 130516 188260 130580 188324
rect 176700 188260 176764 188324
rect 130700 188124 130764 188188
rect 144132 188124 144196 188188
rect 138612 187988 138676 188052
rect 198780 187988 198844 188052
rect 176148 187716 176212 187780
rect 142292 187580 142356 187644
rect 161980 187444 162044 187508
rect 152780 187368 152844 187372
rect 152780 187312 152794 187368
rect 152794 187312 152844 187368
rect 152780 187308 152844 187312
rect 163268 187308 163332 187372
rect 136404 187036 136468 187100
rect 178540 187036 178604 187100
rect 137692 186220 137756 186284
rect 165292 185812 165356 185876
rect 168972 185812 169036 185876
rect 147444 184044 147508 184108
rect 125180 183772 125244 183836
rect 164924 182548 164988 182612
rect 142108 180916 142172 180980
rect 122972 180780 123036 180844
rect 142108 180704 142172 180708
rect 142108 180648 142122 180704
rect 142122 180648 142172 180704
rect 142108 180644 142172 180648
rect 196020 179284 196084 179348
rect 142108 171260 142172 171324
rect 142108 170852 142172 170916
rect 142108 161528 142172 161532
rect 142108 161472 142122 161528
rect 142122 161472 142172 161528
rect 142108 161468 142172 161472
rect 142108 161392 142172 161396
rect 142108 161336 142122 161392
rect 142122 161336 142172 161392
rect 142108 161332 142172 161336
rect 162348 154396 162412 154460
rect 186084 152492 186148 152556
rect 142108 151948 142172 152012
rect 142108 151540 142172 151604
rect 142660 151132 142724 151196
rect 142476 150996 142540 151060
rect 182772 150316 182836 150380
rect 201724 150316 201788 150380
rect 203012 150316 203076 150380
rect 183876 150180 183940 150244
rect 201540 150044 201604 150108
rect 185164 149908 185228 149972
rect 184060 149772 184124 149836
rect 185348 149636 185412 149700
rect 181116 149500 181180 149564
rect 122788 149016 122852 149020
rect 122788 148960 122838 149016
rect 122838 148960 122852 149016
rect 122788 148956 122852 148960
rect 122972 148412 123036 148476
rect 197860 147732 197924 147796
rect 182956 147324 183020 147388
rect 181300 147188 181364 147252
rect 202828 147052 202892 147116
rect 143580 146916 143644 146980
rect 179828 146916 179892 146980
rect 116900 146236 116964 146300
rect 193996 146236 194060 146300
rect 199332 146236 199396 146300
rect 112852 146100 112916 146164
rect 193812 146100 193876 146164
rect 111564 145964 111628 146028
rect 111380 145828 111444 145892
rect 194732 145828 194796 145892
rect 116716 145692 116780 145756
rect 118372 145692 118436 145756
rect 193260 145692 193324 145756
rect 118188 145556 118252 145620
rect 119660 144740 119724 144804
rect 196204 144740 196268 144804
rect 113956 144604 114020 144668
rect 197492 144604 197556 144668
rect 114140 144468 114204 144532
rect 193444 144468 193508 144532
rect 115428 144332 115492 144396
rect 187924 144332 187988 144396
rect 115796 144196 115860 144260
rect 193628 144196 193692 144260
rect 119844 144060 119908 144124
rect 192340 144060 192404 144124
rect 113772 143924 113836 143988
rect 192156 143924 192220 143988
rect 113036 143788 113100 143852
rect 188108 143244 188172 143308
rect 122420 143108 122484 143172
rect 188292 143108 188356 143172
rect 120948 142972 121012 143036
rect 121132 142836 121196 142900
rect 187740 142836 187804 142900
rect 122236 142700 122300 142764
rect 189028 142700 189092 142764
rect 142108 142352 142172 142356
rect 142108 142296 142122 142352
rect 142122 142296 142172 142352
rect 142108 142292 142172 142296
rect 191604 142156 191668 142220
rect 189580 142020 189644 142084
rect 115612 141612 115676 141676
rect 118556 141476 118620 141540
rect 177620 141612 177684 141676
rect 141740 141476 141804 141540
rect 191972 141476 192036 141540
rect 117084 141340 117148 141404
rect 189396 141340 189460 141404
rect 141372 141204 141436 141268
rect 177436 141204 177500 141268
rect 188292 141068 188356 141132
rect 189764 140932 189828 140996
rect 192340 140796 192404 140860
rect 120580 140524 120644 140588
rect 190684 140388 190748 140452
rect 126284 140252 126348 140316
rect 122604 139980 122668 140044
rect 178724 140116 178788 140180
rect 185900 140176 185964 140180
rect 185900 140120 185914 140176
rect 185914 140120 185964 140176
rect 123524 139980 123588 140044
rect 180012 139980 180076 140044
rect 119844 139844 119908 139908
rect 185900 140116 185964 140120
rect 189028 140116 189092 140180
rect 181668 140040 181732 140044
rect 181668 139984 181682 140040
rect 181682 139984 181732 140040
rect 181668 139980 181732 139984
rect 188660 139980 188724 140044
rect 191972 139844 192036 139908
rect 187740 139708 187804 139772
rect 122052 139572 122116 139636
rect 120764 139436 120828 139500
rect 122420 139300 122484 139364
rect 124812 139300 124876 139364
rect 126468 139300 126532 139364
rect 130332 139300 130396 139364
rect 131804 139300 131868 139364
rect 150940 139360 151004 139364
rect 150940 139304 150990 139360
rect 150990 139304 151004 139360
rect 119660 138620 119724 138684
rect 150940 139300 151004 139304
rect 154804 139300 154868 139364
rect 155356 139300 155420 139364
rect 159220 139300 159284 139364
rect 159956 139300 160020 139364
rect 185900 138892 185964 138956
rect 181668 138756 181732 138820
rect 119476 138076 119540 138140
rect 200804 138076 200868 138140
rect 186084 137940 186148 138004
rect 122788 132500 122852 132564
rect 122788 132364 122852 132428
rect 188660 125564 188724 125628
rect 122788 122844 122852 122908
rect 122788 122708 122852 122772
rect 122788 113188 122852 113252
rect 122788 113052 122852 113116
rect 188292 111828 188356 111892
rect 122788 103532 122852 103596
rect 122788 103396 122852 103460
rect 120580 96596 120644 96660
rect 122788 93876 122852 93940
rect 122788 93740 122852 93804
rect 122788 84220 122852 84284
rect 122788 84084 122852 84148
rect 137140 81636 137204 81700
rect 142292 81636 142356 81700
rect 138244 81500 138308 81564
rect 130516 81228 130580 81292
rect 144684 81228 144748 81292
rect 174124 81228 174188 81292
rect 174860 81228 174924 81292
rect 126836 81092 126900 81156
rect 145052 81092 145116 81156
rect 150020 81092 150084 81156
rect 158668 81092 158732 81156
rect 171364 81092 171428 81156
rect 125180 80956 125244 81020
rect 144500 80956 144564 81020
rect 159404 80956 159468 81020
rect 180012 80956 180076 81020
rect 126652 80820 126716 80884
rect 146340 80820 146404 80884
rect 162532 80820 162596 80884
rect 168420 80820 168484 80884
rect 170628 80820 170692 80884
rect 126284 80412 126348 80476
rect 145972 80684 146036 80748
rect 167684 80684 167748 80748
rect 177252 80684 177316 80748
rect 177436 80684 177500 80748
rect 178540 80684 178604 80748
rect 182588 80744 182652 80748
rect 182588 80688 182602 80744
rect 182602 80688 182652 80744
rect 182588 80684 182652 80688
rect 130700 80548 130764 80612
rect 143580 80548 143644 80612
rect 175228 80548 175292 80612
rect 131804 80472 131868 80476
rect 131804 80416 131854 80472
rect 131854 80416 131868 80472
rect 131804 80412 131868 80416
rect 135668 80412 135732 80476
rect 123524 80276 123588 80340
rect 148548 80412 148612 80476
rect 149468 80276 149532 80340
rect 160508 80276 160572 80340
rect 132908 79868 132972 79932
rect 133276 79868 133340 79932
rect 134380 80004 134444 80068
rect 135116 80004 135180 80068
rect 135668 80004 135732 80068
rect 139900 80140 139964 80204
rect 133644 79868 133708 79932
rect 134564 79868 134628 79932
rect 136220 79868 136284 79932
rect 140084 80004 140148 80068
rect 140820 80004 140884 80068
rect 136772 79928 136836 79932
rect 136772 79872 136776 79928
rect 136776 79872 136832 79928
rect 136832 79872 136836 79928
rect 136772 79868 136836 79872
rect 137140 79906 137144 79932
rect 137144 79906 137200 79932
rect 137200 79906 137204 79932
rect 137140 79868 137204 79906
rect 137692 79868 137756 79932
rect 138244 79868 138308 79932
rect 138796 79868 138860 79932
rect 138980 79868 139044 79932
rect 140268 79868 140332 79932
rect 131252 79596 131316 79660
rect 131620 79596 131684 79660
rect 133460 79596 133524 79660
rect 134196 79656 134260 79660
rect 134196 79600 134246 79656
rect 134246 79600 134260 79656
rect 134196 79596 134260 79600
rect 136036 79596 136100 79660
rect 136588 79596 136652 79660
rect 137140 79596 137204 79660
rect 124812 79460 124876 79524
rect 134748 79460 134812 79524
rect 135484 79520 135548 79524
rect 135484 79464 135534 79520
rect 135534 79464 135548 79520
rect 135484 79460 135548 79464
rect 135852 79460 135916 79524
rect 137324 79460 137388 79524
rect 137508 79460 137572 79524
rect 138244 79732 138308 79796
rect 139532 79792 139596 79796
rect 139532 79736 139536 79792
rect 139536 79736 139592 79792
rect 139592 79736 139596 79792
rect 139532 79732 139596 79736
rect 140636 79792 140700 79796
rect 140636 79736 140650 79792
rect 140650 79736 140700 79792
rect 140636 79732 140700 79736
rect 138612 79596 138676 79660
rect 139348 79596 139412 79660
rect 144500 80004 144564 80068
rect 141188 79868 141252 79932
rect 142844 79868 142908 79932
rect 146708 80004 146772 80068
rect 148364 80140 148428 80204
rect 149100 80140 149164 80204
rect 149284 80140 149348 80204
rect 143212 79868 143276 79932
rect 143764 79928 143828 79932
rect 143764 79872 143768 79928
rect 143768 79872 143824 79928
rect 143824 79872 143828 79928
rect 143764 79868 143828 79872
rect 144500 79928 144564 79932
rect 144500 79872 144504 79928
rect 144504 79872 144560 79928
rect 144560 79872 144564 79928
rect 144500 79868 144564 79872
rect 145420 79868 145484 79932
rect 146340 79868 146404 79932
rect 143028 79732 143092 79796
rect 144684 79732 144748 79796
rect 143580 79596 143644 79660
rect 147444 79868 147508 79932
rect 147628 79928 147692 79932
rect 147628 79872 147632 79928
rect 147632 79872 147688 79928
rect 147688 79872 147692 79928
rect 147628 79868 147692 79872
rect 147996 79928 148060 79932
rect 147996 79872 148000 79928
rect 148000 79872 148056 79928
rect 148056 79872 148060 79928
rect 147996 79868 148060 79872
rect 148364 79868 148428 79932
rect 146892 79732 146956 79796
rect 145604 79596 145668 79660
rect 148364 79596 148428 79660
rect 150204 80004 150268 80068
rect 149836 79868 149900 79932
rect 151124 80140 151188 80204
rect 156460 80140 156524 80204
rect 151124 80004 151188 80068
rect 151676 80004 151740 80068
rect 155356 80004 155420 80068
rect 152412 79868 152476 79932
rect 152780 79894 152844 79932
rect 152780 79868 152784 79894
rect 152784 79868 152840 79894
rect 152840 79868 152844 79894
rect 154252 79868 154316 79932
rect 151308 79792 151372 79796
rect 151308 79736 151322 79792
rect 151322 79736 151372 79792
rect 151308 79732 151372 79736
rect 151860 79732 151924 79796
rect 150940 79596 151004 79660
rect 152596 79596 152660 79660
rect 153884 79732 153948 79796
rect 155356 79868 155420 79932
rect 155540 79732 155604 79796
rect 155724 79732 155788 79796
rect 154804 79656 154868 79660
rect 154804 79600 154854 79656
rect 154854 79600 154868 79656
rect 154804 79596 154868 79600
rect 130332 79324 130396 79388
rect 139900 79324 139964 79388
rect 140452 79324 140516 79388
rect 141004 79324 141068 79388
rect 141372 79384 141436 79388
rect 141372 79328 141386 79384
rect 141386 79328 141436 79384
rect 141372 79324 141436 79328
rect 141740 79324 141804 79388
rect 143580 79324 143644 79388
rect 145052 79324 145116 79388
rect 145972 79324 146036 79388
rect 147076 79324 147140 79388
rect 147996 79384 148060 79388
rect 147996 79328 148046 79384
rect 148046 79328 148060 79384
rect 147996 79324 148060 79328
rect 148548 79324 148612 79388
rect 149652 79460 149716 79524
rect 151492 79460 151556 79524
rect 152228 79460 152292 79524
rect 153516 79520 153580 79524
rect 153516 79464 153530 79520
rect 153530 79464 153580 79520
rect 153516 79460 153580 79464
rect 153700 79460 153764 79524
rect 156460 79906 156464 79932
rect 156464 79906 156520 79932
rect 156520 79906 156524 79932
rect 157196 80004 157260 80068
rect 156460 79868 156524 79906
rect 157702 79868 157766 79932
rect 158116 79868 158180 79932
rect 157012 79792 157076 79796
rect 157012 79736 157016 79792
rect 157016 79736 157072 79792
rect 157072 79736 157076 79792
rect 157012 79732 157076 79736
rect 156276 79596 156340 79660
rect 158300 79792 158364 79796
rect 158300 79736 158304 79792
rect 158304 79736 158360 79792
rect 158360 79736 158364 79792
rect 158300 79732 158364 79736
rect 159220 80004 159284 80068
rect 161060 80004 161124 80068
rect 158852 79868 158916 79932
rect 158484 79656 158548 79660
rect 158484 79600 158498 79656
rect 158498 79600 158548 79656
rect 158484 79596 158548 79600
rect 159588 79732 159652 79796
rect 160692 79732 160756 79796
rect 161612 79732 161676 79796
rect 162716 80412 162780 80476
rect 167316 80140 167380 80204
rect 163636 80004 163700 80068
rect 162348 79868 162412 79932
rect 164004 79868 164068 79932
rect 165108 79868 165172 79932
rect 165292 79868 165356 79932
rect 166028 79868 166092 79932
rect 166764 79868 166828 79932
rect 167500 79868 167564 79932
rect 163452 79732 163516 79796
rect 164740 79792 164804 79796
rect 164740 79736 164744 79792
rect 164744 79736 164800 79792
rect 164800 79736 164804 79792
rect 164740 79732 164804 79736
rect 166580 79732 166644 79796
rect 169708 80140 169772 80204
rect 168420 79928 168484 79932
rect 168420 79872 168424 79928
rect 168424 79872 168480 79928
rect 168480 79872 168484 79928
rect 168420 79868 168484 79872
rect 169156 79868 169220 79932
rect 170444 80140 170508 80204
rect 174124 80004 174188 80068
rect 170076 79906 170080 79932
rect 170080 79906 170136 79932
rect 170136 79906 170140 79932
rect 170076 79868 170140 79906
rect 170812 79868 170876 79932
rect 171732 79868 171796 79932
rect 172100 79868 172164 79932
rect 173388 79868 173452 79932
rect 169524 79792 169588 79796
rect 169524 79736 169574 79792
rect 169574 79736 169588 79792
rect 161980 79596 162044 79660
rect 169524 79732 169588 79736
rect 169892 79732 169956 79796
rect 170260 79732 170324 79796
rect 171732 79732 171796 79796
rect 172836 79732 172900 79796
rect 158116 79460 158180 79524
rect 159036 79460 159100 79524
rect 160508 79460 160572 79524
rect 161060 79520 161124 79524
rect 161060 79464 161110 79520
rect 161110 79464 161124 79520
rect 161060 79460 161124 79464
rect 167500 79596 167564 79660
rect 167868 79596 167932 79660
rect 168788 79596 168852 79660
rect 169340 79656 169404 79660
rect 169340 79600 169390 79656
rect 169390 79600 169404 79656
rect 169340 79596 169404 79600
rect 170628 79596 170692 79660
rect 171916 79596 171980 79660
rect 172652 79656 172716 79660
rect 174860 79928 174924 79932
rect 174860 79872 174864 79928
rect 174864 79872 174920 79928
rect 174920 79872 174924 79928
rect 174860 79868 174924 79872
rect 174308 79732 174372 79796
rect 177252 80276 177316 80340
rect 184980 80276 185044 80340
rect 175596 79868 175660 79932
rect 176700 79868 176764 79932
rect 177620 79928 177684 79932
rect 177620 79872 177634 79928
rect 177634 79872 177684 79928
rect 175596 79732 175660 79796
rect 175964 79792 176028 79796
rect 175964 79736 176014 79792
rect 176014 79736 176028 79792
rect 175964 79732 176028 79736
rect 176332 79792 176396 79796
rect 176332 79736 176336 79792
rect 176336 79736 176392 79792
rect 176392 79736 176396 79792
rect 176332 79732 176396 79736
rect 177620 79868 177684 79872
rect 176884 79732 176948 79796
rect 196572 80004 196636 80068
rect 172652 79600 172666 79656
rect 172666 79600 172716 79656
rect 172652 79596 172716 79600
rect 174492 79596 174556 79660
rect 175044 79596 175108 79660
rect 175228 79596 175292 79660
rect 176516 79596 176580 79660
rect 163268 79460 163332 79524
rect 155540 79384 155604 79388
rect 155540 79328 155590 79384
rect 155590 79328 155604 79384
rect 125364 79188 125428 79252
rect 147076 79188 147140 79252
rect 148180 79188 148244 79252
rect 148548 79188 148612 79252
rect 148732 79248 148796 79252
rect 148732 79192 148746 79248
rect 148746 79192 148796 79248
rect 148732 79188 148796 79192
rect 149100 79188 149164 79252
rect 155540 79324 155604 79328
rect 149836 79188 149900 79252
rect 154620 79188 154684 79252
rect 157012 79248 157076 79252
rect 158300 79324 158364 79388
rect 162164 79324 162228 79388
rect 162900 79324 162964 79388
rect 164556 79384 164620 79388
rect 164556 79328 164606 79384
rect 164606 79328 164620 79384
rect 164556 79324 164620 79328
rect 165844 79324 165908 79388
rect 168052 79324 168116 79388
rect 168972 79324 169036 79388
rect 171364 79324 171428 79388
rect 171548 79324 171612 79388
rect 173020 79384 173084 79388
rect 173020 79328 173034 79384
rect 173034 79328 173084 79384
rect 173020 79324 173084 79328
rect 173204 79384 173268 79388
rect 173204 79328 173254 79384
rect 173254 79328 173268 79384
rect 173204 79324 173268 79328
rect 173572 79324 173636 79388
rect 174676 79324 174740 79388
rect 175412 79324 175476 79388
rect 175780 79324 175844 79388
rect 157012 79192 157026 79248
rect 157026 79192 157076 79248
rect 157012 79188 157076 79192
rect 158300 79188 158364 79252
rect 164924 79188 164988 79252
rect 166212 79188 166276 79252
rect 167684 79188 167748 79252
rect 170812 79188 170876 79252
rect 170996 79248 171060 79252
rect 170996 79192 171010 79248
rect 171010 79192 171060 79248
rect 170996 79188 171060 79192
rect 171916 79248 171980 79252
rect 171916 79192 171966 79248
rect 171966 79192 171980 79248
rect 171916 79188 171980 79192
rect 187188 79324 187252 79388
rect 191604 79324 191668 79388
rect 177068 79188 177132 79252
rect 187740 79188 187804 79252
rect 119476 79052 119540 79116
rect 156644 79052 156708 79116
rect 159404 79052 159468 79116
rect 161244 79052 161308 79116
rect 191972 79052 192036 79116
rect 122604 78916 122668 78980
rect 158668 78916 158732 78980
rect 163820 78916 163884 78980
rect 190684 78916 190748 78980
rect 122420 78780 122484 78844
rect 157932 78780 157996 78844
rect 165476 78780 165540 78844
rect 166580 78840 166644 78844
rect 166580 78784 166630 78840
rect 166630 78784 166644 78840
rect 166580 78780 166644 78784
rect 126468 78644 126532 78708
rect 146708 78644 146772 78708
rect 120028 78508 120092 78572
rect 121316 78508 121380 78572
rect 134748 78508 134812 78572
rect 135668 78508 135732 78572
rect 124076 78432 124140 78436
rect 124076 78376 124090 78432
rect 124090 78376 124140 78432
rect 124076 78372 124140 78376
rect 124996 78372 125060 78436
rect 139900 78508 139964 78572
rect 141924 78508 141988 78572
rect 144132 78508 144196 78572
rect 146340 78568 146404 78572
rect 146340 78512 146390 78568
rect 146390 78512 146404 78568
rect 146340 78508 146404 78512
rect 138796 78372 138860 78436
rect 147812 78644 147876 78708
rect 149100 78508 149164 78572
rect 150204 78508 150268 78572
rect 151492 78568 151556 78572
rect 151492 78512 151506 78568
rect 151506 78512 151556 78568
rect 151492 78508 151556 78512
rect 154068 78644 154132 78708
rect 159956 78644 160020 78708
rect 171732 78644 171796 78708
rect 172100 78644 172164 78708
rect 178356 78644 178420 78708
rect 158668 78508 158732 78572
rect 161244 78568 161308 78572
rect 161244 78512 161258 78568
rect 161258 78512 161308 78568
rect 161244 78508 161308 78512
rect 163820 78568 163884 78572
rect 163820 78512 163834 78568
rect 163834 78512 163884 78568
rect 163820 78508 163884 78512
rect 128124 78236 128188 78300
rect 160692 78372 160756 78436
rect 165292 78432 165356 78436
rect 165292 78376 165342 78432
rect 165342 78376 165356 78432
rect 165292 78372 165356 78376
rect 178172 78372 178236 78436
rect 132172 78100 132236 78164
rect 130884 77964 130948 78028
rect 131988 77828 132052 77892
rect 147996 77964 148060 78028
rect 148916 77964 148980 78028
rect 160876 78236 160940 78300
rect 173388 78236 173452 78300
rect 154252 78160 154316 78164
rect 154252 78104 154302 78160
rect 154302 78104 154316 78160
rect 154252 78100 154316 78104
rect 158484 78160 158548 78164
rect 158484 78104 158534 78160
rect 158534 78104 158548 78160
rect 158484 78100 158548 78104
rect 166396 78100 166460 78164
rect 164924 77964 164988 78028
rect 166580 77964 166644 78028
rect 171548 77964 171612 78028
rect 138244 77888 138308 77892
rect 138244 77832 138258 77888
rect 138258 77832 138308 77888
rect 138244 77828 138308 77832
rect 153700 77828 153764 77892
rect 203196 77964 203260 78028
rect 134012 77752 134076 77756
rect 134012 77696 134062 77752
rect 134062 77696 134076 77752
rect 134012 77692 134076 77696
rect 135116 77752 135180 77756
rect 135116 77696 135166 77752
rect 135166 77696 135180 77752
rect 135116 77692 135180 77696
rect 135852 77692 135916 77756
rect 138060 77752 138124 77756
rect 138060 77696 138110 77752
rect 138110 77696 138124 77752
rect 138060 77692 138124 77696
rect 139716 77692 139780 77756
rect 143764 77692 143828 77756
rect 145236 77692 145300 77756
rect 136404 77556 136468 77620
rect 139900 77556 139964 77620
rect 141004 77616 141068 77620
rect 141004 77560 141018 77616
rect 141018 77560 141068 77616
rect 141004 77556 141068 77560
rect 162716 77556 162780 77620
rect 201724 77556 201788 77620
rect 135300 77420 135364 77484
rect 140084 77420 140148 77484
rect 127572 77284 127636 77348
rect 175964 77284 176028 77348
rect 179644 77284 179708 77348
rect 163268 77148 163332 77212
rect 175964 77148 176028 77212
rect 179828 77208 179892 77212
rect 179828 77152 179878 77208
rect 179878 77152 179892 77208
rect 179828 77148 179892 77152
rect 181300 77208 181364 77212
rect 181300 77152 181350 77208
rect 181350 77152 181364 77208
rect 181300 77148 181364 77152
rect 147628 77012 147692 77076
rect 162532 77072 162596 77076
rect 162532 77016 162546 77072
rect 162546 77016 162596 77072
rect 162532 77012 162596 77016
rect 174492 77012 174556 77076
rect 176516 77072 176580 77076
rect 176516 77016 176530 77072
rect 176530 77016 176580 77072
rect 176516 77012 176580 77016
rect 162348 76876 162412 76940
rect 142660 76740 142724 76804
rect 152964 76740 153028 76804
rect 174124 76740 174188 76804
rect 136220 76604 136284 76668
rect 142844 76664 142908 76668
rect 142844 76608 142894 76664
rect 142894 76608 142908 76664
rect 142844 76604 142908 76608
rect 146892 76664 146956 76668
rect 146892 76608 146906 76664
rect 146906 76608 146956 76664
rect 146892 76604 146956 76608
rect 154252 76604 154316 76668
rect 167316 76468 167380 76532
rect 187004 76468 187068 76532
rect 187556 76468 187620 76532
rect 147444 76332 147508 76396
rect 147812 76332 147876 76396
rect 179460 76332 179524 76396
rect 145236 76196 145300 76260
rect 183692 76196 183756 76260
rect 167316 76060 167380 76124
rect 170076 76060 170140 76124
rect 133828 75924 133892 75988
rect 143028 75924 143092 75988
rect 143212 75984 143276 75988
rect 143212 75928 143226 75984
rect 143226 75928 143276 75984
rect 143212 75924 143276 75928
rect 152596 75924 152660 75988
rect 159036 75924 159100 75988
rect 160876 75984 160940 75988
rect 160876 75928 160890 75984
rect 160890 75928 160940 75984
rect 160876 75924 160940 75928
rect 166212 75924 166276 75988
rect 167684 75924 167748 75988
rect 171732 75924 171796 75988
rect 172100 75984 172164 75988
rect 172100 75928 172114 75984
rect 172114 75928 172164 75984
rect 172100 75924 172164 75928
rect 147812 75788 147876 75852
rect 156828 75848 156892 75852
rect 156828 75792 156842 75848
rect 156842 75792 156892 75848
rect 156828 75788 156892 75792
rect 167868 75788 167932 75852
rect 138060 75652 138124 75716
rect 160692 75652 160756 75716
rect 168052 75652 168116 75716
rect 145236 75516 145300 75580
rect 185348 75516 185412 75580
rect 138428 75380 138492 75444
rect 189028 75380 189092 75444
rect 190316 75380 190380 75444
rect 134380 75244 134444 75308
rect 120028 75108 120092 75172
rect 173756 75108 173820 75172
rect 176332 75108 176396 75172
rect 144132 74972 144196 75036
rect 178724 74972 178788 75036
rect 122788 74564 122852 74628
rect 152412 74564 152476 74628
rect 144316 74428 144380 74492
rect 172284 74292 172348 74356
rect 201540 74292 201604 74356
rect 184060 74156 184124 74220
rect 147996 74020 148060 74084
rect 182956 74020 183020 74084
rect 147076 73884 147140 73948
rect 181116 73884 181180 73948
rect 157932 73748 157996 73812
rect 163268 73612 163332 73676
rect 165292 73612 165356 73676
rect 119660 73068 119724 73132
rect 183876 73068 183940 73132
rect 149284 72932 149348 72996
rect 149836 72932 149900 72996
rect 185164 72932 185228 72996
rect 139900 72660 139964 72724
rect 158668 72660 158732 72724
rect 182772 72660 182836 72724
rect 148364 72524 148428 72588
rect 144500 71708 144564 71772
rect 146892 71708 146956 71772
rect 180932 71708 180996 71772
rect 187556 71768 187620 71772
rect 187556 71712 187606 71768
rect 187606 71712 187620 71768
rect 187556 71708 187620 71712
rect 190316 71768 190380 71772
rect 190316 71712 190366 71768
rect 190366 71712 190380 71768
rect 190316 71708 190380 71712
rect 151124 71572 151188 71636
rect 175596 71572 175660 71636
rect 152412 71436 152476 71500
rect 149100 71300 149164 71364
rect 183692 71300 183756 71364
rect 138244 71164 138308 71228
rect 190500 71164 190564 71228
rect 189212 71028 189276 71092
rect 122972 70484 123036 70548
rect 147996 70484 148060 70548
rect 124076 70348 124140 70412
rect 142108 70408 142172 70412
rect 142108 70352 142122 70408
rect 142122 70352 142172 70408
rect 142108 70348 142172 70352
rect 147812 70348 147876 70412
rect 199332 70348 199396 70412
rect 119844 70212 119908 70276
rect 153700 70212 153764 70276
rect 122972 70076 123036 70140
rect 124076 69940 124140 70004
rect 194548 69532 194612 69596
rect 196020 68852 196084 68916
rect 179460 68308 179524 68372
rect 131252 68172 131316 68236
rect 147628 68172 147692 68236
rect 143580 67492 143644 67556
rect 144500 67492 144564 67556
rect 164924 67492 164988 67556
rect 200804 67552 200868 67556
rect 200804 67496 200854 67552
rect 200854 67496 200868 67552
rect 200804 67492 200868 67496
rect 135852 67356 135916 67420
rect 139716 67220 139780 67284
rect 147260 67220 147324 67284
rect 141004 67084 141068 67148
rect 147996 67084 148060 67148
rect 133092 66812 133156 66876
rect 170260 66812 170324 66876
rect 171916 66132 171980 66196
rect 193996 66192 194060 66196
rect 193996 66136 194046 66192
rect 194046 66136 194060 66192
rect 193996 66132 194060 66136
rect 193812 65452 193876 65516
rect 139532 64772 139596 64836
rect 152596 64772 152660 64836
rect 172100 64636 172164 64700
rect 174860 64500 174924 64564
rect 191788 64092 191852 64156
rect 152780 63412 152844 63476
rect 165108 63276 165172 63340
rect 155540 63140 155604 63204
rect 145420 63004 145484 63068
rect 172284 63004 172348 63068
rect 197860 62868 197924 62932
rect 175964 62732 176028 62796
rect 198780 62732 198844 62796
rect 166212 62052 166276 62116
rect 151492 61916 151556 61980
rect 180564 61916 180628 61980
rect 154252 61780 154316 61844
rect 156644 61644 156708 61708
rect 176148 61508 176212 61572
rect 197308 61508 197372 61572
rect 152964 60556 153028 60620
rect 158116 60420 158180 60484
rect 155724 60148 155788 60212
rect 173572 59876 173636 59940
rect 135668 59196 135732 59260
rect 160692 59196 160756 59260
rect 154068 59060 154132 59124
rect 151676 58924 151740 58988
rect 183692 58924 183756 58988
rect 158300 58652 158364 58716
rect 122052 57972 122116 58036
rect 134012 57836 134076 57900
rect 156828 57836 156892 57900
rect 165292 57700 165356 57764
rect 174492 57156 174556 57220
rect 162348 56476 162412 56540
rect 200620 56536 200684 56540
rect 200620 56480 200670 56536
rect 200670 56480 200684 56536
rect 200620 56476 200684 56480
rect 170444 56340 170508 56404
rect 149836 56068 149900 56132
rect 146892 55796 146956 55860
rect 160876 55116 160940 55180
rect 165476 54980 165540 55044
rect 139348 53756 139412 53820
rect 157012 53756 157076 53820
rect 162532 53620 162596 53684
rect 158852 53484 158916 53548
rect 166396 53212 166460 53276
rect 133828 52396 133892 52460
rect 163268 52396 163332 52460
rect 161244 52260 161308 52324
rect 161060 52124 161124 52188
rect 166580 50900 166644 50964
rect 162716 50764 162780 50828
rect 159036 50628 159100 50692
rect 177068 50220 177132 50284
rect 135484 49540 135548 49604
rect 167500 49540 167564 49604
rect 163452 49404 163516 49468
rect 169340 49268 169404 49332
rect 135300 48180 135364 48244
rect 166764 48180 166828 48244
rect 163636 48044 163700 48108
rect 173756 47908 173820 47972
rect 203012 47908 203076 47972
rect 204116 47908 204180 47972
rect 204116 47500 204180 47564
rect 136588 46820 136652 46884
rect 167684 46820 167748 46884
rect 148180 46276 148244 46340
rect 192340 45596 192404 45660
rect 167868 45460 167932 45524
rect 157196 45324 157260 45388
rect 176332 44916 176396 44980
rect 176516 44780 176580 44844
rect 168052 44100 168116 44164
rect 169524 43964 169588 44028
rect 149652 42060 149716 42124
rect 133644 36484 133708 36548
rect 134564 33764 134628 33828
rect 120764 31724 120828 31788
rect 189764 31724 189828 31788
rect 144500 30908 144564 30972
rect 151124 29548 151188 29612
rect 153700 26828 153764 26892
rect 144316 21252 144380 21316
rect 145604 18532 145668 18596
rect 152412 12956 152476 13020
rect 144132 8876 144196 8940
rect 148548 7516 148612 7580
rect 158484 6156 158548 6220
rect 142660 3300 142724 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 112851 265164 112917 265165
rect 112851 265100 112852 265164
rect 112916 265100 112917 265164
rect 112851 265099 112917 265100
rect 111563 261084 111629 261085
rect 111563 261020 111564 261084
rect 111628 261020 111629 261084
rect 111563 261019 111629 261020
rect 111379 260948 111445 260949
rect 111379 260884 111380 260948
rect 111444 260884 111445 260948
rect 111379 260883 111445 260884
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 111382 145893 111442 260883
rect 111566 146029 111626 261019
rect 112854 146165 112914 265099
rect 113035 265028 113101 265029
rect 113035 264964 113036 265028
rect 113100 264964 113101 265028
rect 113035 264963 113101 264964
rect 112851 146164 112917 146165
rect 112851 146100 112852 146164
rect 112916 146100 112917 146164
rect 112851 146099 112917 146100
rect 111563 146028 111629 146029
rect 111563 145964 111564 146028
rect 111628 145964 111629 146028
rect 111563 145963 111629 145964
rect 111379 145892 111445 145893
rect 111379 145828 111380 145892
rect 111444 145828 111445 145892
rect 111379 145827 111445 145828
rect 113038 143853 113098 264963
rect 113771 262988 113837 262989
rect 113771 262924 113772 262988
rect 113836 262924 113837 262988
rect 113771 262923 113837 262924
rect 113774 143989 113834 262923
rect 113955 262852 114021 262853
rect 113955 262788 113956 262852
rect 114020 262788 114021 262852
rect 113955 262787 114021 262788
rect 113958 144669 114018 262787
rect 114139 262444 114205 262445
rect 114139 262380 114140 262444
rect 114204 262380 114205 262444
rect 114139 262379 114205 262380
rect 113955 144668 114021 144669
rect 113955 144604 113956 144668
rect 114020 144604 114021 144668
rect 113955 144603 114021 144604
rect 114142 144533 114202 262379
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 115795 263804 115861 263805
rect 115795 263740 115796 263804
rect 115860 263740 115861 263804
rect 115795 263739 115861 263740
rect 115427 262580 115493 262581
rect 115427 262516 115428 262580
rect 115492 262516 115493 262580
rect 115427 262515 115493 262516
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114139 144532 114205 144533
rect 114139 144468 114140 144532
rect 114204 144468 114205 144532
rect 114139 144467 114205 144468
rect 113771 143988 113837 143989
rect 113771 143924 113772 143988
rect 113836 143924 113837 143988
rect 113771 143923 113837 143924
rect 113035 143852 113101 143853
rect 113035 143788 113036 143852
rect 113100 143788 113101 143852
rect 113035 143787 113101 143788
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 115954 114914 151398
rect 115430 144397 115490 262515
rect 115611 260540 115677 260541
rect 115611 260476 115612 260540
rect 115676 260476 115677 260540
rect 115611 260475 115677 260476
rect 115427 144396 115493 144397
rect 115427 144332 115428 144396
rect 115492 144332 115493 144396
rect 115427 144331 115493 144332
rect 115614 141677 115674 260475
rect 115798 144261 115858 263739
rect 118371 263668 118437 263669
rect 118371 263604 118372 263668
rect 118436 263604 118437 263668
rect 118371 263603 118437 263604
rect 116899 263260 116965 263261
rect 116899 263196 116900 263260
rect 116964 263196 116965 263260
rect 116899 263195 116965 263196
rect 116715 259724 116781 259725
rect 116715 259660 116716 259724
rect 116780 259660 116781 259724
rect 116715 259659 116781 259660
rect 116718 145757 116778 259659
rect 116902 146301 116962 263195
rect 118187 262716 118253 262717
rect 118187 262652 118188 262716
rect 118252 262652 118253 262716
rect 118187 262651 118253 262652
rect 117083 260404 117149 260405
rect 117083 260340 117084 260404
rect 117148 260340 117149 260404
rect 117083 260339 117149 260340
rect 116899 146300 116965 146301
rect 116899 146236 116900 146300
rect 116964 146236 116965 146300
rect 116899 146235 116965 146236
rect 116715 145756 116781 145757
rect 116715 145692 116716 145756
rect 116780 145692 116781 145756
rect 116715 145691 116781 145692
rect 115795 144260 115861 144261
rect 115795 144196 115796 144260
rect 115860 144196 115861 144260
rect 115795 144195 115861 144196
rect 115611 141676 115677 141677
rect 115611 141612 115612 141676
rect 115676 141612 115677 141676
rect 115611 141611 115677 141612
rect 117086 141405 117146 260339
rect 118190 145621 118250 262651
rect 118374 145757 118434 263603
rect 118794 262000 119414 263898
rect 122603 263940 122669 263941
rect 122603 263876 122604 263940
rect 122668 263876 122669 263940
rect 122603 263875 122669 263876
rect 119843 263124 119909 263125
rect 119843 263060 119844 263124
rect 119908 263060 119909 263124
rect 119843 263059 119909 263060
rect 118555 260132 118621 260133
rect 118555 260068 118556 260132
rect 118620 260068 118621 260132
rect 118555 260067 118621 260068
rect 118371 145756 118437 145757
rect 118371 145692 118372 145756
rect 118436 145692 118437 145756
rect 118371 145691 118437 145692
rect 118187 145620 118253 145621
rect 118187 145556 118188 145620
rect 118252 145556 118253 145620
rect 118187 145555 118253 145556
rect 118558 141541 118618 260067
rect 119659 259996 119725 259997
rect 119659 259932 119660 259996
rect 119724 259932 119725 259996
rect 119659 259931 119725 259932
rect 118794 192454 119414 198000
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 119662 144805 119722 259931
rect 119659 144804 119725 144805
rect 119659 144740 119660 144804
rect 119724 144740 119725 144804
rect 119659 144739 119725 144740
rect 119846 144125 119906 263059
rect 120947 260268 121013 260269
rect 120947 260204 120948 260268
rect 121012 260204 121013 260268
rect 120947 260203 121013 260204
rect 119843 144124 119909 144125
rect 119843 144060 119844 144124
rect 119908 144060 119909 144124
rect 119843 144059 119909 144060
rect 120950 143037 121010 260203
rect 122235 259860 122301 259861
rect 122235 259796 122236 259860
rect 122300 259796 122301 259860
rect 122235 259795 122301 259796
rect 121131 259588 121197 259589
rect 121131 259524 121132 259588
rect 121196 259524 121197 259588
rect 121131 259523 121197 259524
rect 120947 143036 121013 143037
rect 120947 142972 120948 143036
rect 121012 142972 121013 143036
rect 120947 142971 121013 142972
rect 121134 142901 121194 259523
rect 122238 209810 122298 259795
rect 122606 257410 122666 263875
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 187371 284340 187437 284341
rect 187371 284276 187372 284340
rect 187436 284276 187437 284340
rect 187371 284275 187437 284276
rect 123155 259588 123221 259589
rect 123155 259524 123156 259588
rect 123220 259524 123221 259588
rect 123155 259523 123221 259524
rect 124075 259588 124141 259589
rect 124075 259524 124076 259588
rect 124140 259524 124141 259588
rect 124075 259523 124141 259524
rect 186083 259588 186149 259589
rect 186083 259524 186084 259588
rect 186148 259524 186149 259588
rect 186083 259523 186149 259524
rect 122971 259452 123037 259453
rect 122971 259388 122972 259452
rect 123036 259388 123037 259452
rect 122971 259387 123037 259388
rect 122974 258090 123034 259387
rect 122422 257350 122666 257410
rect 122790 258030 123034 258090
rect 122790 257410 122850 258030
rect 122790 257350 123034 257410
rect 122422 248570 122482 257350
rect 122974 256730 123034 257350
rect 122606 256670 123034 256730
rect 122606 249250 122666 256670
rect 122606 249190 123034 249250
rect 122974 248570 123034 249190
rect 122422 248510 122666 248570
rect 122606 248430 122666 248510
rect 122422 248370 122666 248430
rect 122790 248510 123034 248570
rect 122422 238770 122482 248370
rect 122790 247890 122850 248510
rect 122606 247830 122850 247890
rect 122606 239050 122666 247830
rect 122606 238990 122850 239050
rect 122422 238710 122666 238770
rect 122606 238370 122666 238710
rect 122422 238310 122666 238370
rect 122790 238370 122850 238990
rect 122790 238310 123034 238370
rect 122422 229530 122482 238310
rect 122974 237690 123034 238310
rect 122606 237630 123034 237690
rect 122606 230210 122666 237630
rect 122606 230150 123034 230210
rect 122974 229530 123034 230150
rect 122422 229470 122666 229530
rect 122606 229110 122666 229470
rect 122422 229050 122666 229110
rect 122790 229470 123034 229530
rect 122422 219450 122482 229050
rect 122790 228850 122850 229470
rect 122606 228790 122850 228850
rect 122606 220010 122666 228790
rect 122606 219950 123034 220010
rect 122974 219450 123034 219950
rect 122422 219390 122666 219450
rect 122606 219330 122666 219390
rect 122422 219270 122666 219330
rect 122790 219390 123034 219450
rect 122790 219330 122850 219390
rect 122790 219270 123034 219330
rect 122422 210490 122482 219270
rect 122974 218650 123034 219270
rect 122606 218590 123034 218650
rect 122606 211170 122666 218590
rect 122606 211110 123034 211170
rect 122974 210490 123034 211110
rect 122422 210430 122666 210490
rect 122238 209750 122482 209810
rect 121315 195260 121381 195261
rect 121315 195196 121316 195260
rect 121380 195196 121381 195260
rect 121315 195195 121381 195196
rect 121131 142900 121197 142901
rect 121131 142836 121132 142900
rect 121196 142836 121197 142900
rect 121131 142835 121197 142836
rect 118555 141540 118621 141541
rect 118555 141476 118556 141540
rect 118620 141476 118621 141540
rect 118555 141475 118621 141476
rect 117083 141404 117149 141405
rect 117083 141340 117084 141404
rect 117148 141340 117149 141404
rect 117083 141339 117149 141340
rect 120579 140588 120645 140589
rect 120579 140524 120580 140588
rect 120644 140524 120645 140588
rect 120579 140523 120645 140524
rect 119843 139908 119909 139909
rect 119843 139844 119844 139908
rect 119908 139844 119909 139908
rect 119843 139843 119909 139844
rect 119659 138684 119725 138685
rect 119659 138620 119660 138684
rect 119724 138620 119725 138684
rect 119659 138619 119725 138620
rect 119475 138140 119541 138141
rect 119475 138076 119476 138140
rect 119540 138076 119541 138140
rect 119475 138075 119541 138076
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 119478 79117 119538 138075
rect 119475 79116 119541 79117
rect 119475 79052 119476 79116
rect 119540 79052 119541 79116
rect 119475 79051 119541 79052
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 119662 73133 119722 138619
rect 119659 73132 119725 73133
rect 119659 73068 119660 73132
rect 119724 73068 119725 73132
rect 119659 73067 119725 73068
rect 119846 70277 119906 139843
rect 120582 96661 120642 140523
rect 120763 139500 120829 139501
rect 120763 139436 120764 139500
rect 120828 139436 120829 139500
rect 120763 139435 120829 139436
rect 120579 96660 120645 96661
rect 120579 96596 120580 96660
rect 120644 96596 120645 96660
rect 120579 96595 120645 96596
rect 120027 78572 120093 78573
rect 120027 78508 120028 78572
rect 120092 78508 120093 78572
rect 120027 78507 120093 78508
rect 120030 75173 120090 78507
rect 120027 75172 120093 75173
rect 120027 75108 120028 75172
rect 120092 75108 120093 75172
rect 120027 75107 120093 75108
rect 119843 70276 119909 70277
rect 119843 70212 119844 70276
rect 119908 70212 119909 70276
rect 119843 70211 119909 70212
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 120766 31789 120826 139435
rect 121318 78573 121378 195195
rect 122422 180810 122482 209750
rect 122238 180750 122482 180810
rect 122238 142765 122298 180750
rect 122606 180570 122666 210430
rect 122790 210430 123034 210490
rect 122790 209677 122850 210430
rect 123158 209810 123218 259523
rect 122974 209750 123218 209810
rect 122787 209676 122853 209677
rect 122787 209612 122788 209676
rect 122852 209612 122853 209676
rect 122787 209611 122853 209612
rect 122787 205596 122853 205597
rect 122787 205532 122788 205596
rect 122852 205532 122853 205596
rect 122787 205531 122853 205532
rect 122790 196077 122850 205531
rect 122974 200565 123034 209750
rect 123891 200972 123957 200973
rect 123891 200908 123892 200972
rect 123956 200908 123957 200972
rect 123891 200907 123957 200908
rect 122971 200564 123037 200565
rect 122971 200500 122972 200564
rect 123036 200500 123037 200564
rect 122971 200499 123037 200500
rect 123894 198250 123954 200907
rect 124078 200701 124138 259523
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 186086 213893 186146 259523
rect 186083 213892 186149 213893
rect 186083 213828 186084 213892
rect 186148 213828 186149 213892
rect 186083 213827 186149 213828
rect 153515 200972 153581 200973
rect 153515 200908 153516 200972
rect 153580 200908 153581 200972
rect 153515 200907 153581 200908
rect 170995 200972 171061 200973
rect 170995 200908 170996 200972
rect 171060 200908 171061 200972
rect 170995 200907 171061 200908
rect 124075 200700 124141 200701
rect 124075 200636 124076 200700
rect 124140 200636 124141 200700
rect 124075 200635 124141 200636
rect 142843 200564 142909 200565
rect 142843 200500 142844 200564
rect 142908 200500 142909 200564
rect 142843 200499 142909 200500
rect 138979 200428 139045 200429
rect 138979 200364 138980 200428
rect 139044 200364 139045 200428
rect 138979 200363 139045 200364
rect 132539 199884 132605 199885
rect 132539 199820 132540 199884
rect 132604 199820 132605 199884
rect 132539 199819 132605 199820
rect 133091 199884 133157 199885
rect 133091 199820 133092 199884
rect 133156 199882 133157 199884
rect 134011 199884 134077 199885
rect 133156 199822 133338 199882
rect 133156 199820 133157 199822
rect 133091 199819 133157 199820
rect 126835 198388 126901 198389
rect 126835 198324 126836 198388
rect 126900 198324 126901 198388
rect 126835 198323 126901 198324
rect 123894 198190 124138 198250
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 122787 196076 122853 196077
rect 122787 196012 122788 196076
rect 122852 196012 122853 196076
rect 122787 196011 122853 196012
rect 122787 190500 122853 190501
rect 122787 190436 122788 190500
rect 122852 190436 122853 190500
rect 122787 190435 122853 190436
rect 122790 190365 122850 190435
rect 122787 190364 122853 190365
rect 122787 190300 122788 190364
rect 122852 190300 122853 190364
rect 122787 190299 122853 190300
rect 122971 180844 123037 180845
rect 122971 180780 122972 180844
rect 123036 180780 123037 180844
rect 122971 180779 123037 180780
rect 122422 180510 122666 180570
rect 122422 171730 122482 180510
rect 122974 179890 123034 180779
rect 122606 179830 123034 179890
rect 122606 172410 122666 179830
rect 122606 172350 123034 172410
rect 122422 171670 122666 171730
rect 122606 171150 122666 171670
rect 122422 171090 122666 171150
rect 122422 161490 122482 171090
rect 122974 170370 123034 172350
rect 122606 170310 123034 170370
rect 122606 162210 122666 170310
rect 122606 162150 123034 162210
rect 122422 161430 122666 161490
rect 122606 160850 122666 161430
rect 122422 160790 122666 160850
rect 122422 152010 122482 160790
rect 122974 160170 123034 162150
rect 122606 160110 123034 160170
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 122606 152690 122666 160110
rect 122606 152630 123034 152690
rect 122422 151950 122666 152010
rect 122606 151830 122666 151950
rect 122422 151770 122666 151830
rect 122422 143173 122482 151770
rect 122974 151330 123034 152630
rect 122606 151270 123034 151330
rect 122606 149290 122666 151270
rect 122606 149230 122850 149290
rect 122790 149021 122850 149230
rect 122787 149020 122853 149021
rect 122787 148956 122788 149020
rect 122852 148956 122853 149020
rect 122787 148955 122853 148956
rect 122971 148476 123037 148477
rect 122971 148412 122972 148476
rect 123036 148412 123037 148476
rect 122971 148411 123037 148412
rect 122419 143172 122485 143173
rect 122419 143108 122420 143172
rect 122484 143108 122485 143172
rect 122419 143107 122485 143108
rect 122235 142764 122301 142765
rect 122235 142700 122236 142764
rect 122300 142700 122301 142764
rect 122235 142699 122301 142700
rect 122603 140044 122669 140045
rect 122603 139980 122604 140044
rect 122668 139980 122669 140044
rect 122603 139979 122669 139980
rect 122051 139636 122117 139637
rect 122051 139572 122052 139636
rect 122116 139572 122117 139636
rect 122051 139571 122117 139572
rect 121315 78572 121381 78573
rect 121315 78508 121316 78572
rect 121380 78508 121381 78572
rect 121315 78507 121381 78508
rect 122054 58037 122114 139571
rect 122419 139364 122485 139365
rect 122419 139300 122420 139364
rect 122484 139300 122485 139364
rect 122419 139299 122485 139300
rect 122422 78845 122482 139299
rect 122606 78981 122666 139979
rect 122787 132564 122853 132565
rect 122787 132500 122788 132564
rect 122852 132500 122853 132564
rect 122787 132499 122853 132500
rect 122790 132429 122850 132499
rect 122787 132428 122853 132429
rect 122787 132364 122788 132428
rect 122852 132364 122853 132428
rect 122787 132363 122853 132364
rect 122787 122908 122853 122909
rect 122787 122844 122788 122908
rect 122852 122844 122853 122908
rect 122787 122843 122853 122844
rect 122790 122773 122850 122843
rect 122787 122772 122853 122773
rect 122787 122708 122788 122772
rect 122852 122708 122853 122772
rect 122787 122707 122853 122708
rect 122787 113252 122853 113253
rect 122787 113188 122788 113252
rect 122852 113188 122853 113252
rect 122787 113187 122853 113188
rect 122790 113117 122850 113187
rect 122787 113116 122853 113117
rect 122787 113052 122788 113116
rect 122852 113052 122853 113116
rect 122787 113051 122853 113052
rect 122787 103596 122853 103597
rect 122787 103532 122788 103596
rect 122852 103532 122853 103596
rect 122787 103531 122853 103532
rect 122790 103461 122850 103531
rect 122787 103460 122853 103461
rect 122787 103396 122788 103460
rect 122852 103396 122853 103460
rect 122787 103395 122853 103396
rect 122787 93940 122853 93941
rect 122787 93876 122788 93940
rect 122852 93876 122853 93940
rect 122787 93875 122853 93876
rect 122790 93805 122850 93875
rect 122787 93804 122853 93805
rect 122787 93740 122788 93804
rect 122852 93740 122853 93804
rect 122787 93739 122853 93740
rect 122787 84284 122853 84285
rect 122787 84220 122788 84284
rect 122852 84220 122853 84284
rect 122787 84219 122853 84220
rect 122790 84149 122850 84219
rect 122787 84148 122853 84149
rect 122787 84084 122788 84148
rect 122852 84084 122853 84148
rect 122787 84083 122853 84084
rect 122603 78980 122669 78981
rect 122603 78916 122604 78980
rect 122668 78916 122669 78980
rect 122603 78915 122669 78916
rect 122419 78844 122485 78845
rect 122419 78780 122420 78844
rect 122484 78780 122485 78844
rect 122419 78779 122485 78780
rect 122787 74628 122853 74629
rect 122787 74564 122788 74628
rect 122852 74564 122853 74628
rect 122787 74563 122853 74564
rect 122790 74490 122850 74563
rect 122606 74430 122850 74490
rect 122606 70410 122666 74430
rect 122974 70549 123034 148411
rect 123294 142000 123914 160398
rect 123523 140044 123589 140045
rect 123523 139980 123524 140044
rect 123588 139980 123589 140044
rect 123523 139979 123589 139980
rect 123526 80341 123586 139979
rect 123523 80340 123589 80341
rect 123523 80276 123524 80340
rect 123588 80276 123589 80340
rect 123523 80275 123589 80276
rect 124078 78437 124138 198190
rect 125363 198116 125429 198117
rect 125363 198052 125364 198116
rect 125428 198052 125429 198116
rect 125363 198051 125429 198052
rect 124995 194036 125061 194037
rect 124995 193972 124996 194036
rect 125060 193972 125061 194036
rect 124995 193971 125061 193972
rect 124811 139364 124877 139365
rect 124811 139300 124812 139364
rect 124876 139300 124877 139364
rect 124811 139299 124877 139300
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 124814 79525 124874 139299
rect 124811 79524 124877 79525
rect 124811 79460 124812 79524
rect 124876 79460 124877 79524
rect 124811 79459 124877 79460
rect 124998 78437 125058 193971
rect 125179 183836 125245 183837
rect 125179 183772 125180 183836
rect 125244 183772 125245 183836
rect 125179 183771 125245 183772
rect 125182 81021 125242 183771
rect 125179 81020 125245 81021
rect 125179 80956 125180 81020
rect 125244 80956 125245 81020
rect 125179 80955 125245 80956
rect 125366 79253 125426 198051
rect 126651 197980 126717 197981
rect 126651 197916 126652 197980
rect 126716 197916 126717 197980
rect 126651 197915 126717 197916
rect 126283 140316 126349 140317
rect 126283 140252 126284 140316
rect 126348 140252 126349 140316
rect 126283 140251 126349 140252
rect 126286 80477 126346 140251
rect 126467 139364 126533 139365
rect 126467 139300 126468 139364
rect 126532 139300 126533 139364
rect 126467 139299 126533 139300
rect 126283 80476 126349 80477
rect 126283 80412 126284 80476
rect 126348 80412 126349 80476
rect 126283 80411 126349 80412
rect 125363 79252 125429 79253
rect 125363 79188 125364 79252
rect 125428 79188 125429 79252
rect 125363 79187 125429 79188
rect 126470 78709 126530 139299
rect 126654 80885 126714 197915
rect 126838 81157 126898 198323
rect 131987 195804 132053 195805
rect 131987 195740 131988 195804
rect 132052 195740 132053 195804
rect 131987 195739 132053 195740
rect 128123 195668 128189 195669
rect 128123 195604 128124 195668
rect 128188 195604 128189 195668
rect 128123 195603 128189 195604
rect 127939 195532 128005 195533
rect 127939 195468 127940 195532
rect 128004 195468 128005 195532
rect 127939 195467 128005 195468
rect 127942 84210 128002 195467
rect 127574 84150 128002 84210
rect 126835 81156 126901 81157
rect 126835 81092 126836 81156
rect 126900 81092 126901 81156
rect 126835 81091 126901 81092
rect 126651 80884 126717 80885
rect 126651 80820 126652 80884
rect 126716 80820 126717 80884
rect 126651 80819 126717 80820
rect 126467 78708 126533 78709
rect 126467 78644 126468 78708
rect 126532 78644 126533 78708
rect 126467 78643 126533 78644
rect 124075 78436 124141 78437
rect 124075 78372 124076 78436
rect 124140 78372 124141 78436
rect 124075 78371 124141 78372
rect 124995 78436 125061 78437
rect 124995 78372 124996 78436
rect 125060 78372 125061 78436
rect 124995 78371 125061 78372
rect 122971 70548 123037 70549
rect 122971 70484 122972 70548
rect 123036 70484 123037 70548
rect 122971 70483 123037 70484
rect 122606 70350 123034 70410
rect 122974 70141 123034 70350
rect 122971 70140 123037 70141
rect 122971 70076 122972 70140
rect 123036 70076 123037 70140
rect 122971 70075 123037 70076
rect 122051 58036 122117 58037
rect 122051 57972 122052 58036
rect 122116 57972 122117 58036
rect 122051 57971 122117 57972
rect 123294 52954 123914 78000
rect 127574 77349 127634 84150
rect 128126 78301 128186 195603
rect 130883 195124 130949 195125
rect 130883 195060 130884 195124
rect 130948 195060 130949 195124
rect 130883 195059 130949 195060
rect 130515 188324 130581 188325
rect 130515 188260 130516 188324
rect 130580 188260 130581 188324
rect 130515 188259 130581 188260
rect 130331 139364 130397 139365
rect 130331 139300 130332 139364
rect 130396 139300 130397 139364
rect 130331 139299 130397 139300
rect 130334 79389 130394 139299
rect 130518 81293 130578 188259
rect 130699 188188 130765 188189
rect 130699 188124 130700 188188
rect 130764 188124 130765 188188
rect 130699 188123 130765 188124
rect 130515 81292 130581 81293
rect 130515 81228 130516 81292
rect 130580 81228 130581 81292
rect 130515 81227 130581 81228
rect 130702 80613 130762 188123
rect 130699 80612 130765 80613
rect 130699 80548 130700 80612
rect 130764 80548 130765 80612
rect 130699 80547 130765 80548
rect 130331 79388 130397 79389
rect 130331 79324 130332 79388
rect 130396 79324 130397 79388
rect 130331 79323 130397 79324
rect 128123 78300 128189 78301
rect 128123 78236 128124 78300
rect 128188 78236 128189 78300
rect 128123 78235 128189 78236
rect 130886 78029 130946 195059
rect 131619 188460 131685 188461
rect 131619 188396 131620 188460
rect 131684 188396 131685 188460
rect 131619 188395 131685 188396
rect 131622 79661 131682 188395
rect 131803 139364 131869 139365
rect 131803 139300 131804 139364
rect 131868 139300 131869 139364
rect 131803 139299 131869 139300
rect 131806 80477 131866 139299
rect 131803 80476 131869 80477
rect 131803 80412 131804 80476
rect 131868 80412 131869 80476
rect 131803 80411 131869 80412
rect 131251 79660 131317 79661
rect 131251 79596 131252 79660
rect 131316 79596 131317 79660
rect 131251 79595 131317 79596
rect 131619 79660 131685 79661
rect 131619 79596 131620 79660
rect 131684 79596 131685 79660
rect 131619 79595 131685 79596
rect 130883 78028 130949 78029
rect 127571 77348 127637 77349
rect 127571 77284 127572 77348
rect 127636 77284 127637 77348
rect 127571 77283 127637 77284
rect 124075 70412 124141 70413
rect 124075 70348 124076 70412
rect 124140 70348 124141 70412
rect 124075 70347 124141 70348
rect 124078 70005 124138 70347
rect 124075 70004 124141 70005
rect 124075 69940 124076 70004
rect 124140 69940 124141 70004
rect 124075 69939 124141 69940
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 120763 31788 120829 31789
rect 120763 31724 120764 31788
rect 120828 31724 120829 31788
rect 120763 31723 120829 31724
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 130883 77964 130884 78028
rect 130948 77964 130949 78028
rect 130883 77963 130949 77964
rect 131254 68237 131314 79595
rect 131990 77893 132050 195739
rect 132171 195260 132237 195261
rect 132171 195196 132172 195260
rect 132236 195196 132237 195260
rect 132171 195195 132237 195196
rect 132174 78165 132234 195195
rect 132542 194610 132602 199819
rect 133091 199340 133157 199341
rect 133091 199276 133092 199340
rect 133156 199276 133157 199340
rect 133091 199275 133157 199276
rect 132542 194550 132970 194610
rect 132910 79933 132970 194550
rect 133094 88350 133154 199275
rect 133278 193901 133338 199822
rect 134011 199820 134012 199884
rect 134076 199882 134077 199884
rect 134563 199884 134629 199885
rect 134076 199822 134442 199882
rect 134076 199820 134077 199822
rect 134011 199819 134077 199820
rect 133643 198524 133709 198525
rect 133643 198460 133644 198524
rect 133708 198460 133709 198524
rect 133643 198459 133709 198460
rect 133459 197436 133525 197437
rect 133459 197372 133460 197436
rect 133524 197372 133525 197436
rect 133459 197371 133525 197372
rect 133275 193900 133341 193901
rect 133275 193836 133276 193900
rect 133340 193836 133341 193900
rect 133275 193835 133341 193836
rect 133094 88290 133338 88350
rect 133278 79933 133338 88290
rect 132907 79932 132973 79933
rect 132907 79868 132908 79932
rect 132972 79868 132973 79932
rect 132907 79867 132973 79868
rect 133275 79932 133341 79933
rect 133275 79868 133276 79932
rect 133340 79868 133341 79932
rect 133275 79867 133341 79868
rect 132171 78164 132237 78165
rect 132171 78100 132172 78164
rect 132236 78100 132237 78164
rect 132171 78099 132237 78100
rect 131987 77892 132053 77893
rect 131987 77828 131988 77892
rect 132052 77828 132053 77892
rect 131987 77827 132053 77828
rect 131251 68236 131317 68237
rect 131251 68172 131252 68236
rect 131316 68172 131317 68236
rect 131251 68171 131317 68172
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 133278 70410 133338 79867
rect 133462 79661 133522 197371
rect 133646 79933 133706 198459
rect 134195 197436 134261 197437
rect 134195 197372 134196 197436
rect 134260 197372 134261 197436
rect 134195 197371 134261 197372
rect 133643 79932 133709 79933
rect 133643 79868 133644 79932
rect 133708 79868 133709 79932
rect 133643 79867 133709 79868
rect 133459 79660 133525 79661
rect 133459 79596 133460 79660
rect 133524 79596 133525 79660
rect 133459 79595 133525 79596
rect 133094 70350 133338 70410
rect 133094 66877 133154 70350
rect 133091 66876 133157 66877
rect 133091 66812 133092 66876
rect 133156 66812 133157 66876
rect 133091 66811 133157 66812
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 133646 36549 133706 79867
rect 134198 79661 134258 197371
rect 134382 196210 134442 199822
rect 134563 199820 134564 199884
rect 134628 199820 134629 199884
rect 134563 199819 134629 199820
rect 135851 199884 135917 199885
rect 135851 199820 135852 199884
rect 135916 199820 135917 199884
rect 135851 199819 135917 199820
rect 136219 199884 136285 199885
rect 136219 199820 136220 199884
rect 136284 199820 136285 199884
rect 136219 199819 136285 199820
rect 137139 199884 137205 199885
rect 137139 199820 137140 199884
rect 137204 199820 137205 199884
rect 137139 199819 137205 199820
rect 137507 199884 137573 199885
rect 137507 199820 137508 199884
rect 137572 199820 137573 199884
rect 137507 199819 137573 199820
rect 137691 199884 137757 199885
rect 137691 199820 137692 199884
rect 137756 199820 137757 199884
rect 137691 199819 137757 199820
rect 138427 199884 138493 199885
rect 138427 199820 138428 199884
rect 138492 199820 138493 199884
rect 138427 199819 138493 199820
rect 134566 198750 134626 199819
rect 134566 198690 134810 198750
rect 134382 196150 134626 196210
rect 134379 189140 134445 189141
rect 134379 189076 134380 189140
rect 134444 189076 134445 189140
rect 134379 189075 134445 189076
rect 134382 80069 134442 189075
rect 134379 80068 134445 80069
rect 134379 80004 134380 80068
rect 134444 80004 134445 80068
rect 134379 80003 134445 80004
rect 134195 79660 134261 79661
rect 134195 79596 134196 79660
rect 134260 79596 134261 79660
rect 134195 79595 134261 79596
rect 134011 77756 134077 77757
rect 134011 77692 134012 77756
rect 134076 77692 134077 77756
rect 134011 77691 134077 77692
rect 133827 75988 133893 75989
rect 133827 75924 133828 75988
rect 133892 75924 133893 75988
rect 133827 75923 133893 75924
rect 133830 52461 133890 75923
rect 134014 57901 134074 77691
rect 134382 75309 134442 80003
rect 134566 79933 134626 196150
rect 134563 79932 134629 79933
rect 134563 79868 134564 79932
rect 134628 79868 134629 79932
rect 134563 79867 134629 79868
rect 134379 75308 134445 75309
rect 134379 75244 134380 75308
rect 134444 75244 134445 75308
rect 134379 75243 134445 75244
rect 134011 57900 134077 57901
rect 134011 57836 134012 57900
rect 134076 57836 134077 57900
rect 134011 57835 134077 57836
rect 133827 52460 133893 52461
rect 133827 52396 133828 52460
rect 133892 52396 133893 52460
rect 133827 52395 133893 52396
rect 133643 36548 133709 36549
rect 133643 36484 133644 36548
rect 133708 36484 133709 36548
rect 133643 36483 133709 36484
rect 134566 33829 134626 79867
rect 134750 79525 134810 198690
rect 135854 196349 135914 199819
rect 135851 196348 135917 196349
rect 135851 196284 135852 196348
rect 135916 196284 135917 196348
rect 135851 196283 135917 196284
rect 135851 196212 135917 196213
rect 135851 196148 135852 196212
rect 135916 196148 135917 196212
rect 135851 196147 135917 196148
rect 135667 80476 135733 80477
rect 135667 80412 135668 80476
rect 135732 80412 135733 80476
rect 135667 80411 135733 80412
rect 135670 80069 135730 80411
rect 135115 80068 135181 80069
rect 135115 80004 135116 80068
rect 135180 80004 135181 80068
rect 135115 80003 135181 80004
rect 135667 80068 135733 80069
rect 135667 80004 135668 80068
rect 135732 80004 135733 80068
rect 135667 80003 135733 80004
rect 134747 79524 134813 79525
rect 134747 79460 134748 79524
rect 134812 79460 134813 79524
rect 134747 79459 134813 79460
rect 134750 78573 134810 79459
rect 134747 78572 134813 78573
rect 134747 78508 134748 78572
rect 134812 78508 134813 78572
rect 134747 78507 134813 78508
rect 135118 77757 135178 80003
rect 135854 79525 135914 196147
rect 136222 196077 136282 199819
rect 136219 196076 136285 196077
rect 136219 196012 136220 196076
rect 136284 196012 136285 196076
rect 136219 196011 136285 196012
rect 137142 194989 137202 199819
rect 137510 198933 137570 199819
rect 137507 198932 137573 198933
rect 137507 198868 137508 198932
rect 137572 198868 137573 198932
rect 137507 198867 137573 198868
rect 136219 194988 136285 194989
rect 136219 194924 136220 194988
rect 136284 194924 136285 194988
rect 136219 194923 136285 194924
rect 137139 194988 137205 194989
rect 137139 194924 137140 194988
rect 137204 194924 137205 194988
rect 137139 194923 137205 194924
rect 136035 188460 136101 188461
rect 136035 188396 136036 188460
rect 136100 188396 136101 188460
rect 136035 188395 136101 188396
rect 136038 79661 136098 188395
rect 136222 79933 136282 194923
rect 137694 188730 137754 199819
rect 138430 199477 138490 199819
rect 138982 199477 139042 200363
rect 142846 199885 142906 200499
rect 148915 200020 148981 200021
rect 148915 199956 148916 200020
rect 148980 199956 148981 200020
rect 148915 199955 148981 199956
rect 141923 199884 141989 199885
rect 141923 199820 141924 199884
rect 141988 199820 141989 199884
rect 141923 199819 141989 199820
rect 142659 199884 142725 199885
rect 142659 199820 142660 199884
rect 142724 199820 142725 199884
rect 142659 199819 142725 199820
rect 142843 199884 142909 199885
rect 142843 199820 142844 199884
rect 142908 199820 142909 199884
rect 142843 199819 142909 199820
rect 144131 199884 144197 199885
rect 144131 199820 144132 199884
rect 144196 199820 144197 199884
rect 144131 199819 144197 199820
rect 148363 199884 148429 199885
rect 148363 199820 148364 199884
rect 148428 199820 148429 199884
rect 148363 199819 148429 199820
rect 140451 199748 140517 199749
rect 140451 199684 140452 199748
rect 140516 199684 140517 199748
rect 140451 199683 140517 199684
rect 138427 199476 138493 199477
rect 138427 199412 138428 199476
rect 138492 199412 138493 199476
rect 138427 199411 138493 199412
rect 138795 199476 138861 199477
rect 138795 199412 138796 199476
rect 138860 199412 138861 199476
rect 138795 199411 138861 199412
rect 138979 199476 139045 199477
rect 138979 199412 138980 199476
rect 139044 199412 139045 199476
rect 138979 199411 139045 199412
rect 138059 194988 138125 194989
rect 138059 194924 138060 194988
rect 138124 194924 138125 194988
rect 138059 194923 138125 194924
rect 137694 188670 137938 188730
rect 136587 188460 136653 188461
rect 136587 188396 136588 188460
rect 136652 188396 136653 188460
rect 136587 188395 136653 188396
rect 137507 188460 137573 188461
rect 137507 188396 137508 188460
rect 137572 188396 137573 188460
rect 137507 188395 137573 188396
rect 136403 187100 136469 187101
rect 136403 187036 136404 187100
rect 136468 187036 136469 187100
rect 136403 187035 136469 187036
rect 136219 79932 136285 79933
rect 136219 79868 136220 79932
rect 136284 79868 136285 79932
rect 136219 79867 136285 79868
rect 136035 79660 136101 79661
rect 136035 79596 136036 79660
rect 136100 79596 136101 79660
rect 136035 79595 136101 79596
rect 135483 79524 135549 79525
rect 135483 79460 135484 79524
rect 135548 79460 135549 79524
rect 135483 79459 135549 79460
rect 135851 79524 135917 79525
rect 135851 79460 135852 79524
rect 135916 79460 135917 79524
rect 135851 79459 135917 79460
rect 135115 77756 135181 77757
rect 135115 77692 135116 77756
rect 135180 77692 135181 77756
rect 135115 77691 135181 77692
rect 135299 77484 135365 77485
rect 135299 77420 135300 77484
rect 135364 77420 135365 77484
rect 135299 77419 135365 77420
rect 135302 48245 135362 77419
rect 135486 49605 135546 79459
rect 135667 78572 135733 78573
rect 135667 78508 135668 78572
rect 135732 78508 135733 78572
rect 135667 78507 135733 78508
rect 135670 59261 135730 78507
rect 135851 77756 135917 77757
rect 135851 77692 135852 77756
rect 135916 77692 135917 77756
rect 135851 77691 135917 77692
rect 135854 67421 135914 77691
rect 136222 76669 136282 79867
rect 136406 77621 136466 187035
rect 136590 79661 136650 188395
rect 137139 81700 137205 81701
rect 137139 81636 137140 81700
rect 137204 81636 137205 81700
rect 137139 81635 137205 81636
rect 137142 79933 137202 81635
rect 136771 79932 136837 79933
rect 136771 79868 136772 79932
rect 136836 79868 136837 79932
rect 136771 79867 136837 79868
rect 137139 79932 137205 79933
rect 137139 79868 137140 79932
rect 137204 79868 137205 79932
rect 137139 79867 137205 79868
rect 136587 79660 136653 79661
rect 136587 79596 136588 79660
rect 136652 79596 136653 79660
rect 136587 79595 136653 79596
rect 136774 78162 136834 79867
rect 137142 79661 137202 79867
rect 137139 79660 137205 79661
rect 137139 79596 137140 79660
rect 137204 79596 137205 79660
rect 137139 79595 137205 79596
rect 137510 79525 137570 188395
rect 137691 186284 137757 186285
rect 137691 186220 137692 186284
rect 137756 186220 137757 186284
rect 137691 186219 137757 186220
rect 137694 79933 137754 186219
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 137323 79524 137389 79525
rect 137323 79460 137324 79524
rect 137388 79460 137389 79524
rect 137323 79459 137389 79460
rect 137507 79524 137573 79525
rect 137507 79460 137508 79524
rect 137572 79460 137573 79524
rect 137507 79459 137573 79460
rect 137326 79386 137386 79459
rect 137878 79386 137938 188670
rect 138062 93870 138122 194923
rect 138427 194852 138493 194853
rect 138427 194788 138428 194852
rect 138492 194788 138493 194852
rect 138427 194787 138493 194788
rect 138430 188869 138490 194787
rect 138798 190470 138858 199411
rect 139163 199340 139229 199341
rect 139163 199276 139164 199340
rect 139228 199276 139229 199340
rect 139163 199275 139229 199276
rect 139166 196077 139226 199275
rect 140454 199205 140514 199683
rect 141926 199341 141986 199819
rect 140635 199340 140701 199341
rect 140635 199276 140636 199340
rect 140700 199276 140701 199340
rect 140635 199275 140701 199276
rect 141923 199340 141989 199341
rect 141923 199276 141924 199340
rect 141988 199276 141989 199340
rect 141923 199275 141989 199276
rect 140451 199204 140517 199205
rect 140451 199140 140452 199204
rect 140516 199140 140517 199204
rect 140451 199139 140517 199140
rect 140083 197436 140149 197437
rect 140083 197372 140084 197436
rect 140148 197372 140149 197436
rect 140083 197371 140149 197372
rect 139163 196076 139229 196077
rect 139163 196012 139164 196076
rect 139228 196012 139229 196076
rect 139163 196011 139229 196012
rect 139163 194988 139229 194989
rect 139163 194924 139164 194988
rect 139228 194924 139229 194988
rect 139163 194923 139229 194924
rect 138614 190410 138858 190470
rect 138427 188868 138493 188869
rect 138427 188804 138428 188868
rect 138492 188804 138493 188868
rect 138427 188803 138493 188804
rect 138427 188460 138493 188461
rect 138427 188396 138428 188460
rect 138492 188396 138493 188460
rect 138427 188395 138493 188396
rect 138430 93870 138490 188395
rect 138614 188053 138674 190410
rect 138795 188596 138861 188597
rect 138795 188532 138796 188596
rect 138860 188532 138861 188596
rect 138795 188531 138861 188532
rect 138611 188052 138677 188053
rect 138611 187988 138612 188052
rect 138676 187988 138677 188052
rect 138611 187987 138677 187988
rect 138062 93810 138306 93870
rect 138430 93810 138674 93870
rect 138246 81565 138306 93810
rect 138243 81564 138309 81565
rect 138243 81500 138244 81564
rect 138308 81500 138309 81564
rect 138243 81499 138309 81500
rect 138246 79933 138306 81499
rect 138243 79932 138309 79933
rect 138243 79868 138244 79932
rect 138308 79868 138309 79932
rect 138243 79867 138309 79868
rect 138243 79796 138309 79797
rect 138243 79732 138244 79796
rect 138308 79794 138309 79796
rect 138308 79734 138490 79794
rect 138308 79732 138309 79734
rect 138243 79731 138309 79732
rect 137326 79326 137938 79386
rect 136590 78102 136834 78162
rect 136403 77620 136469 77621
rect 136403 77556 136404 77620
rect 136468 77556 136469 77620
rect 136403 77555 136469 77556
rect 136219 76668 136285 76669
rect 136219 76604 136220 76668
rect 136284 76604 136285 76668
rect 136219 76603 136285 76604
rect 135851 67420 135917 67421
rect 135851 67356 135852 67420
rect 135916 67356 135917 67420
rect 135851 67355 135917 67356
rect 135667 59260 135733 59261
rect 135667 59196 135668 59260
rect 135732 59196 135733 59260
rect 135667 59195 135733 59196
rect 135483 49604 135549 49605
rect 135483 49540 135484 49604
rect 135548 49540 135549 49604
rect 135483 49539 135549 49540
rect 135299 48244 135365 48245
rect 135299 48180 135300 48244
rect 135364 48180 135365 48244
rect 135299 48179 135365 48180
rect 136590 46885 136650 78102
rect 136794 66454 137414 78000
rect 138243 77892 138309 77893
rect 138243 77828 138244 77892
rect 138308 77828 138309 77892
rect 138243 77827 138309 77828
rect 138059 77756 138125 77757
rect 138059 77692 138060 77756
rect 138124 77692 138125 77756
rect 138059 77691 138125 77692
rect 138062 75717 138122 77691
rect 138059 75716 138125 75717
rect 138059 75652 138060 75716
rect 138124 75652 138125 75716
rect 138059 75651 138125 75652
rect 138246 71229 138306 77827
rect 138430 75445 138490 79734
rect 138614 79661 138674 93810
rect 138798 79933 138858 188531
rect 139166 176670 139226 194923
rect 138982 176610 139226 176670
rect 138982 79933 139042 176610
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 139899 80204 139965 80205
rect 139899 80140 139900 80204
rect 139964 80140 139965 80204
rect 139899 80139 139965 80140
rect 138795 79932 138861 79933
rect 138795 79868 138796 79932
rect 138860 79868 138861 79932
rect 138795 79867 138861 79868
rect 138979 79932 139045 79933
rect 138979 79868 138980 79932
rect 139044 79868 139045 79932
rect 138979 79867 139045 79868
rect 138611 79660 138677 79661
rect 138611 79596 138612 79660
rect 138676 79596 138677 79660
rect 138611 79595 138677 79596
rect 138798 78437 138858 79867
rect 139531 79796 139597 79797
rect 139531 79732 139532 79796
rect 139596 79732 139597 79796
rect 139531 79731 139597 79732
rect 139347 79660 139413 79661
rect 139347 79596 139348 79660
rect 139412 79596 139413 79660
rect 139347 79595 139413 79596
rect 138795 78436 138861 78437
rect 138795 78372 138796 78436
rect 138860 78372 138861 78436
rect 138795 78371 138861 78372
rect 138427 75444 138493 75445
rect 138427 75380 138428 75444
rect 138492 75380 138493 75444
rect 138427 75379 138493 75380
rect 138243 71228 138309 71229
rect 138243 71164 138244 71228
rect 138308 71164 138309 71228
rect 138243 71163 138309 71164
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136587 46884 136653 46885
rect 136587 46820 136588 46884
rect 136652 46820 136653 46884
rect 136587 46819 136653 46820
rect 134563 33828 134629 33829
rect 134563 33764 134564 33828
rect 134628 33764 134629 33828
rect 134563 33763 134629 33764
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 139350 53821 139410 79595
rect 139534 64837 139594 79731
rect 139902 79389 139962 80139
rect 140086 80069 140146 197371
rect 140451 188596 140517 188597
rect 140451 188532 140452 188596
rect 140516 188532 140517 188596
rect 140451 188531 140517 188532
rect 140267 188460 140333 188461
rect 140267 188396 140268 188460
rect 140332 188396 140333 188460
rect 140267 188395 140333 188396
rect 140083 80068 140149 80069
rect 140083 80004 140084 80068
rect 140148 80004 140149 80068
rect 140083 80003 140149 80004
rect 140270 79933 140330 188395
rect 140267 79932 140333 79933
rect 140267 79868 140268 79932
rect 140332 79868 140333 79932
rect 140267 79867 140333 79868
rect 140454 79389 140514 188531
rect 140638 79797 140698 199275
rect 141003 191180 141069 191181
rect 141003 191116 141004 191180
rect 141068 191116 141069 191180
rect 141003 191115 141069 191116
rect 140819 190364 140885 190365
rect 140819 190300 140820 190364
rect 140884 190300 140885 190364
rect 140819 190299 140885 190300
rect 140822 80069 140882 190299
rect 140819 80068 140885 80069
rect 140819 80004 140820 80068
rect 140884 80004 140885 80068
rect 140819 80003 140885 80004
rect 141006 79930 141066 191115
rect 141294 178954 141914 198000
rect 142475 191044 142541 191045
rect 142475 190980 142476 191044
rect 142540 190980 142541 191044
rect 142475 190979 142541 190980
rect 142291 187644 142357 187645
rect 142291 187580 142292 187644
rect 142356 187580 142357 187644
rect 142291 187579 142357 187580
rect 142107 180980 142173 180981
rect 142107 180916 142108 180980
rect 142172 180916 142173 180980
rect 142107 180915 142173 180916
rect 142110 180709 142170 180915
rect 142107 180708 142173 180709
rect 142107 180644 142108 180708
rect 142172 180644 142173 180708
rect 142107 180643 142173 180644
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 142107 171324 142173 171325
rect 142107 171260 142108 171324
rect 142172 171260 142173 171324
rect 142107 171259 142173 171260
rect 142110 170917 142170 171259
rect 142107 170916 142173 170917
rect 142107 170852 142108 170916
rect 142172 170852 142173 170916
rect 142107 170851 142173 170852
rect 142107 161532 142173 161533
rect 142107 161468 142108 161532
rect 142172 161468 142173 161532
rect 142107 161467 142173 161468
rect 142110 161397 142170 161467
rect 142107 161396 142173 161397
rect 142107 161332 142108 161396
rect 142172 161332 142173 161396
rect 142107 161331 142173 161332
rect 142107 152012 142173 152013
rect 142107 151948 142108 152012
rect 142172 151948 142173 152012
rect 142107 151947 142173 151948
rect 142110 151605 142170 151947
rect 142107 151604 142173 151605
rect 142107 151540 142108 151604
rect 142172 151540 142173 151604
rect 142107 151539 142173 151540
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 142107 142356 142173 142357
rect 142107 142292 142108 142356
rect 142172 142292 142173 142356
rect 142107 142291 142173 142292
rect 142110 141810 142170 142291
rect 141926 141750 142170 141810
rect 141739 141540 141805 141541
rect 141739 141476 141740 141540
rect 141804 141476 141805 141540
rect 141739 141475 141805 141476
rect 141371 141268 141437 141269
rect 141371 141204 141372 141268
rect 141436 141204 141437 141268
rect 141371 141203 141437 141204
rect 141187 79932 141253 79933
rect 141187 79930 141188 79932
rect 141006 79870 141188 79930
rect 140635 79796 140701 79797
rect 140635 79732 140636 79796
rect 140700 79732 140701 79796
rect 140635 79731 140701 79732
rect 141006 79389 141066 79870
rect 141187 79868 141188 79870
rect 141252 79868 141253 79932
rect 141187 79867 141253 79868
rect 141374 79389 141434 141203
rect 141742 79389 141802 141475
rect 139899 79388 139965 79389
rect 139899 79324 139900 79388
rect 139964 79324 139965 79388
rect 139899 79323 139965 79324
rect 140451 79388 140517 79389
rect 140451 79324 140452 79388
rect 140516 79324 140517 79388
rect 140451 79323 140517 79324
rect 141003 79388 141069 79389
rect 141003 79324 141004 79388
rect 141068 79324 141069 79388
rect 141003 79323 141069 79324
rect 141371 79388 141437 79389
rect 141371 79324 141372 79388
rect 141436 79324 141437 79388
rect 141371 79323 141437 79324
rect 141739 79388 141805 79389
rect 141739 79324 141740 79388
rect 141804 79324 141805 79388
rect 141739 79323 141805 79324
rect 141926 78573 141986 141750
rect 142294 81701 142354 187579
rect 142478 151061 142538 190979
rect 142662 151197 142722 199819
rect 143579 188868 143645 188869
rect 143579 188804 143580 188868
rect 143644 188804 143645 188868
rect 143579 188803 143645 188804
rect 142659 151196 142725 151197
rect 142659 151132 142660 151196
rect 142724 151132 142725 151196
rect 142659 151131 142725 151132
rect 142475 151060 142541 151061
rect 142475 150996 142476 151060
rect 142540 150996 142541 151060
rect 142475 150995 142541 150996
rect 143582 146981 143642 188803
rect 144134 188189 144194 199819
rect 146891 199748 146957 199749
rect 146891 199684 146892 199748
rect 146956 199684 146957 199748
rect 146891 199683 146957 199684
rect 145603 197708 145669 197709
rect 145603 197644 145604 197708
rect 145668 197644 145669 197708
rect 145603 197643 145669 197644
rect 145235 195396 145301 195397
rect 145235 195332 145236 195396
rect 145300 195332 145301 195396
rect 145235 195331 145301 195332
rect 144131 188188 144197 188189
rect 144131 188124 144132 188188
rect 144196 188124 144197 188188
rect 144131 188123 144197 188124
rect 143579 146980 143645 146981
rect 143579 146916 143580 146980
rect 143644 146916 143645 146980
rect 143579 146915 143645 146916
rect 142291 81700 142357 81701
rect 142291 81636 142292 81700
rect 142356 81636 142357 81700
rect 142291 81635 142357 81636
rect 144683 81292 144749 81293
rect 144683 81228 144684 81292
rect 144748 81228 144749 81292
rect 144683 81227 144749 81228
rect 144499 81020 144565 81021
rect 144499 80956 144500 81020
rect 144564 80956 144565 81020
rect 144499 80955 144565 80956
rect 143579 80612 143645 80613
rect 143579 80548 143580 80612
rect 143644 80548 143645 80612
rect 143579 80547 143645 80548
rect 142843 79932 142909 79933
rect 142843 79868 142844 79932
rect 142908 79868 142909 79932
rect 142843 79867 142909 79868
rect 143211 79932 143277 79933
rect 143211 79868 143212 79932
rect 143276 79868 143277 79932
rect 143211 79867 143277 79868
rect 139899 78572 139965 78573
rect 139899 78508 139900 78572
rect 139964 78570 139965 78572
rect 141923 78572 141989 78573
rect 139964 78510 140146 78570
rect 139964 78508 139965 78510
rect 139899 78507 139965 78508
rect 139715 77756 139781 77757
rect 139715 77692 139716 77756
rect 139780 77692 139781 77756
rect 139715 77691 139781 77692
rect 139718 67285 139778 77691
rect 139899 77620 139965 77621
rect 139899 77556 139900 77620
rect 139964 77556 139965 77620
rect 139899 77555 139965 77556
rect 139902 72725 139962 77555
rect 140086 77485 140146 78510
rect 141923 78508 141924 78572
rect 141988 78570 141989 78572
rect 141988 78510 142170 78570
rect 141988 78508 141989 78510
rect 141923 78507 141989 78508
rect 141003 77620 141069 77621
rect 141003 77556 141004 77620
rect 141068 77556 141069 77620
rect 141003 77555 141069 77556
rect 140083 77484 140149 77485
rect 140083 77420 140084 77484
rect 140148 77420 140149 77484
rect 140083 77419 140149 77420
rect 139899 72724 139965 72725
rect 139899 72660 139900 72724
rect 139964 72660 139965 72724
rect 139899 72659 139965 72660
rect 139715 67284 139781 67285
rect 139715 67220 139716 67284
rect 139780 67220 139781 67284
rect 139715 67219 139781 67220
rect 141006 67149 141066 77555
rect 141294 70954 141914 78000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 142110 70413 142170 78510
rect 142659 76804 142725 76805
rect 142659 76740 142660 76804
rect 142724 76740 142725 76804
rect 142659 76739 142725 76740
rect 141003 67148 141069 67149
rect 141003 67084 141004 67148
rect 141068 67084 141069 67148
rect 141003 67083 141069 67084
rect 139531 64836 139597 64837
rect 139531 64772 139532 64836
rect 139596 64772 139597 64836
rect 139531 64771 139597 64772
rect 139347 53820 139413 53821
rect 139347 53756 139348 53820
rect 139412 53756 139413 53820
rect 139347 53755 139413 53756
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 142107 70412 142173 70413
rect 142107 70348 142108 70412
rect 142172 70348 142173 70412
rect 142107 70347 142173 70348
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 142662 3365 142722 76739
rect 142846 76669 142906 79867
rect 143027 79796 143093 79797
rect 143027 79732 143028 79796
rect 143092 79732 143093 79796
rect 143027 79731 143093 79732
rect 142843 76668 142909 76669
rect 142843 76604 142844 76668
rect 142908 76604 142909 76668
rect 142843 76603 142909 76604
rect 143030 75989 143090 79731
rect 143214 75989 143274 79867
rect 143582 79661 143642 80547
rect 144502 80069 144562 80955
rect 144499 80068 144565 80069
rect 144499 80004 144500 80068
rect 144564 80004 144565 80068
rect 144499 80003 144565 80004
rect 143763 79932 143829 79933
rect 143763 79868 143764 79932
rect 143828 79868 143829 79932
rect 143763 79867 143829 79868
rect 144499 79932 144565 79933
rect 144499 79868 144500 79932
rect 144564 79868 144565 79932
rect 144499 79867 144565 79868
rect 143579 79660 143645 79661
rect 143579 79596 143580 79660
rect 143644 79596 143645 79660
rect 143579 79595 143645 79596
rect 143579 79388 143645 79389
rect 143579 79324 143580 79388
rect 143644 79324 143645 79388
rect 143579 79323 143645 79324
rect 143027 75988 143093 75989
rect 143027 75924 143028 75988
rect 143092 75924 143093 75988
rect 143027 75923 143093 75924
rect 143211 75988 143277 75989
rect 143211 75924 143212 75988
rect 143276 75924 143277 75988
rect 143211 75923 143277 75924
rect 143582 67557 143642 79323
rect 143766 77757 143826 79867
rect 144131 78572 144197 78573
rect 144131 78508 144132 78572
rect 144196 78508 144197 78572
rect 144131 78507 144197 78508
rect 143763 77756 143829 77757
rect 143763 77692 143764 77756
rect 143828 77692 143829 77756
rect 143763 77691 143829 77692
rect 144134 75037 144194 78507
rect 144131 75036 144197 75037
rect 144131 74972 144132 75036
rect 144196 74972 144197 75036
rect 144131 74971 144197 74972
rect 143579 67556 143645 67557
rect 143579 67492 143580 67556
rect 143644 67492 143645 67556
rect 143579 67491 143645 67492
rect 144134 8941 144194 74971
rect 144315 74492 144381 74493
rect 144315 74428 144316 74492
rect 144380 74428 144381 74492
rect 144315 74427 144381 74428
rect 144318 21317 144378 74427
rect 144502 71773 144562 79867
rect 144686 79797 144746 81227
rect 145051 81156 145117 81157
rect 145051 81092 145052 81156
rect 145116 81092 145117 81156
rect 145051 81091 145117 81092
rect 144683 79796 144749 79797
rect 144683 79732 144684 79796
rect 144748 79732 144749 79796
rect 144683 79731 144749 79732
rect 145054 79389 145114 81091
rect 145051 79388 145117 79389
rect 145051 79324 145052 79388
rect 145116 79324 145117 79388
rect 145051 79323 145117 79324
rect 145238 77757 145298 195331
rect 145419 191180 145485 191181
rect 145419 191116 145420 191180
rect 145484 191116 145485 191180
rect 145419 191115 145485 191116
rect 145422 79933 145482 191115
rect 145419 79932 145485 79933
rect 145419 79868 145420 79932
rect 145484 79868 145485 79932
rect 145419 79867 145485 79868
rect 145235 77756 145301 77757
rect 145235 77692 145236 77756
rect 145300 77692 145301 77756
rect 145235 77691 145301 77692
rect 145235 76260 145301 76261
rect 145235 76196 145236 76260
rect 145300 76196 145301 76260
rect 145235 76195 145301 76196
rect 145238 75581 145298 76195
rect 145235 75580 145301 75581
rect 145235 75516 145236 75580
rect 145300 75516 145301 75580
rect 145235 75515 145301 75516
rect 144499 71772 144565 71773
rect 144499 71708 144500 71772
rect 144564 71708 144565 71772
rect 144499 71707 144565 71708
rect 145238 70410 145298 75515
rect 145422 73170 145482 79867
rect 145606 79661 145666 197643
rect 145794 183454 146414 198000
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 146339 80884 146405 80885
rect 146339 80820 146340 80884
rect 146404 80820 146405 80884
rect 146339 80819 146405 80820
rect 145971 80748 146037 80749
rect 145971 80684 145972 80748
rect 146036 80684 146037 80748
rect 145971 80683 146037 80684
rect 145603 79660 145669 79661
rect 145603 79596 145604 79660
rect 145668 79596 145669 79660
rect 145603 79595 145669 79596
rect 145974 79389 146034 80683
rect 146342 79933 146402 80819
rect 146707 80068 146773 80069
rect 146707 80004 146708 80068
rect 146772 80004 146773 80068
rect 146707 80003 146773 80004
rect 146339 79932 146405 79933
rect 146339 79868 146340 79932
rect 146404 79868 146405 79932
rect 146339 79867 146405 79868
rect 145971 79388 146037 79389
rect 145971 79324 145972 79388
rect 146036 79324 146037 79388
rect 145971 79323 146037 79324
rect 146342 78573 146402 79867
rect 146710 78709 146770 80003
rect 146894 79797 146954 199683
rect 148179 198796 148245 198797
rect 148179 198732 148180 198796
rect 148244 198732 148245 198796
rect 148179 198731 148245 198732
rect 147075 191180 147141 191181
rect 147075 191116 147076 191180
rect 147140 191116 147141 191180
rect 147075 191115 147141 191116
rect 146891 79796 146957 79797
rect 146891 79732 146892 79796
rect 146956 79732 146957 79796
rect 146891 79731 146957 79732
rect 147078 79389 147138 191115
rect 147443 184108 147509 184109
rect 147443 184044 147444 184108
rect 147508 184044 147509 184108
rect 147443 184043 147509 184044
rect 147446 93870 147506 184043
rect 147446 93810 147690 93870
rect 147630 89730 147690 93810
rect 147630 89670 147874 89730
rect 147443 79932 147509 79933
rect 147443 79868 147444 79932
rect 147508 79868 147509 79932
rect 147443 79867 147509 79868
rect 147627 79932 147693 79933
rect 147627 79868 147628 79932
rect 147692 79868 147693 79932
rect 147627 79867 147693 79868
rect 147075 79388 147141 79389
rect 147075 79324 147076 79388
rect 147140 79324 147141 79388
rect 147075 79323 147141 79324
rect 147075 79252 147141 79253
rect 147075 79188 147076 79252
rect 147140 79188 147141 79252
rect 147075 79187 147141 79188
rect 146707 78708 146773 78709
rect 146707 78644 146708 78708
rect 146772 78644 146773 78708
rect 146707 78643 146773 78644
rect 146339 78572 146405 78573
rect 146339 78508 146340 78572
rect 146404 78508 146405 78572
rect 146339 78507 146405 78508
rect 145794 75454 146414 78000
rect 146891 76668 146957 76669
rect 146891 76604 146892 76668
rect 146956 76604 146957 76668
rect 146891 76603 146957 76604
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145422 73110 145666 73170
rect 145238 70350 145482 70410
rect 144499 67556 144565 67557
rect 144499 67492 144500 67556
rect 144564 67492 144565 67556
rect 144499 67491 144565 67492
rect 144502 30973 144562 67491
rect 145422 63069 145482 70350
rect 145419 63068 145485 63069
rect 145419 63004 145420 63068
rect 145484 63004 145485 63068
rect 145419 63003 145485 63004
rect 144499 30972 144565 30973
rect 144499 30908 144500 30972
rect 144564 30908 144565 30972
rect 144499 30907 144565 30908
rect 144315 21316 144381 21317
rect 144315 21252 144316 21316
rect 144380 21252 144381 21316
rect 144315 21251 144381 21252
rect 145606 18597 145666 73110
rect 145794 39454 146414 74898
rect 146894 71773 146954 76603
rect 147078 73949 147138 79187
rect 147446 76397 147506 79867
rect 147630 77077 147690 79867
rect 147814 78709 147874 89670
rect 147995 79932 148061 79933
rect 147995 79868 147996 79932
rect 148060 79868 148061 79932
rect 147995 79867 148061 79868
rect 147998 79389 148058 79867
rect 147995 79388 148061 79389
rect 147995 79324 147996 79388
rect 148060 79324 148061 79388
rect 147995 79323 148061 79324
rect 148182 79253 148242 198731
rect 148366 80205 148426 199819
rect 148918 195261 148978 199955
rect 149651 199884 149717 199885
rect 149651 199820 149652 199884
rect 149716 199820 149717 199884
rect 149651 199819 149717 199820
rect 150019 199884 150085 199885
rect 150019 199820 150020 199884
rect 150084 199820 150085 199884
rect 150019 199819 150085 199820
rect 151307 199884 151373 199885
rect 151307 199820 151308 199884
rect 151372 199820 151373 199884
rect 151307 199819 151373 199820
rect 152595 199884 152661 199885
rect 152595 199820 152596 199884
rect 152660 199820 152661 199884
rect 152595 199819 152661 199820
rect 149654 195533 149714 199819
rect 150022 195533 150082 199819
rect 149651 195532 149717 195533
rect 149651 195468 149652 195532
rect 149716 195468 149717 195532
rect 149651 195467 149717 195468
rect 150019 195532 150085 195533
rect 150019 195468 150020 195532
rect 150084 195468 150085 195532
rect 150019 195467 150085 195468
rect 148915 195260 148981 195261
rect 148915 195196 148916 195260
rect 148980 195196 148981 195260
rect 148915 195195 148981 195196
rect 149651 195124 149717 195125
rect 149651 195060 149652 195124
rect 149716 195060 149717 195124
rect 149651 195059 149717 195060
rect 148731 194988 148797 194989
rect 148731 194924 148732 194988
rect 148796 194924 148797 194988
rect 148731 194923 148797 194924
rect 148547 80476 148613 80477
rect 148547 80412 148548 80476
rect 148612 80412 148613 80476
rect 148547 80411 148613 80412
rect 148363 80204 148429 80205
rect 148363 80140 148364 80204
rect 148428 80140 148429 80204
rect 148363 80139 148429 80140
rect 148366 79933 148426 80139
rect 148363 79932 148429 79933
rect 148363 79868 148364 79932
rect 148428 79868 148429 79932
rect 148363 79867 148429 79868
rect 148363 79660 148429 79661
rect 148363 79596 148364 79660
rect 148428 79596 148429 79660
rect 148363 79595 148429 79596
rect 148179 79252 148245 79253
rect 148179 79188 148180 79252
rect 148244 79188 148245 79252
rect 148179 79187 148245 79188
rect 147811 78708 147877 78709
rect 147811 78644 147812 78708
rect 147876 78644 147877 78708
rect 147811 78643 147877 78644
rect 147995 78028 148061 78029
rect 147995 77964 147996 78028
rect 148060 77964 148061 78028
rect 147995 77963 148061 77964
rect 147627 77076 147693 77077
rect 147627 77012 147628 77076
rect 147692 77012 147693 77076
rect 147627 77011 147693 77012
rect 147443 76396 147509 76397
rect 147443 76332 147444 76396
rect 147508 76332 147509 76396
rect 147443 76331 147509 76332
rect 147075 73948 147141 73949
rect 147075 73884 147076 73948
rect 147140 73884 147141 73948
rect 147075 73883 147141 73884
rect 146891 71772 146957 71773
rect 146891 71708 146892 71772
rect 146956 71708 146957 71772
rect 146891 71707 146957 71708
rect 147078 70410 147138 73883
rect 147630 73170 147690 77011
rect 147811 76396 147877 76397
rect 147811 76332 147812 76396
rect 147876 76332 147877 76396
rect 147811 76331 147877 76332
rect 147814 75853 147874 76331
rect 147811 75852 147877 75853
rect 147811 75788 147812 75852
rect 147876 75788 147877 75852
rect 147811 75787 147877 75788
rect 146894 70350 147138 70410
rect 147262 73110 147690 73170
rect 146894 55861 146954 70350
rect 147262 67285 147322 73110
rect 147814 71090 147874 75787
rect 147998 74085 148058 77963
rect 147995 74084 148061 74085
rect 147995 74020 147996 74084
rect 148060 74020 148061 74084
rect 147995 74019 148061 74020
rect 147446 71030 147874 71090
rect 147446 70410 147506 71030
rect 147998 70549 148058 74019
rect 148366 72589 148426 79595
rect 148550 79389 148610 80411
rect 148547 79388 148613 79389
rect 148547 79324 148548 79388
rect 148612 79324 148613 79388
rect 148547 79323 148613 79324
rect 148734 79253 148794 194923
rect 148915 191452 148981 191453
rect 148915 191388 148916 191452
rect 148980 191388 148981 191452
rect 148915 191387 148981 191388
rect 148547 79252 148613 79253
rect 148547 79188 148548 79252
rect 148612 79188 148613 79252
rect 148547 79187 148613 79188
rect 148731 79252 148797 79253
rect 148731 79188 148732 79252
rect 148796 79188 148797 79252
rect 148731 79187 148797 79188
rect 148363 72588 148429 72589
rect 148363 72524 148364 72588
rect 148428 72524 148429 72588
rect 148363 72523 148429 72524
rect 147995 70548 148061 70549
rect 147995 70484 147996 70548
rect 148060 70484 148061 70548
rect 147995 70483 148061 70484
rect 147811 70412 147877 70413
rect 147446 70350 147690 70410
rect 147630 68237 147690 70350
rect 147811 70348 147812 70412
rect 147876 70348 147877 70412
rect 148366 70410 148426 72523
rect 148550 71790 148610 79187
rect 148918 78029 148978 191387
rect 149467 191316 149533 191317
rect 149467 191252 149468 191316
rect 149532 191252 149533 191316
rect 149467 191251 149533 191252
rect 149470 80341 149530 191251
rect 149467 80340 149533 80341
rect 149467 80276 149468 80340
rect 149532 80276 149533 80340
rect 149467 80275 149533 80276
rect 149099 80204 149165 80205
rect 149099 80140 149100 80204
rect 149164 80140 149165 80204
rect 149099 80139 149165 80140
rect 149283 80204 149349 80205
rect 149283 80140 149284 80204
rect 149348 80140 149349 80204
rect 149283 80139 149349 80140
rect 149102 79253 149162 80139
rect 149099 79252 149165 79253
rect 149099 79188 149100 79252
rect 149164 79188 149165 79252
rect 149099 79187 149165 79188
rect 149099 78572 149165 78573
rect 149099 78508 149100 78572
rect 149164 78508 149165 78572
rect 149099 78507 149165 78508
rect 148915 78028 148981 78029
rect 148915 77964 148916 78028
rect 148980 77964 148981 78028
rect 148915 77963 148981 77964
rect 148550 71730 148794 71790
rect 148734 70410 148794 71730
rect 149102 71365 149162 78507
rect 149286 72997 149346 80139
rect 149654 79525 149714 195059
rect 150019 191044 150085 191045
rect 150019 190980 150020 191044
rect 150084 190980 150085 191044
rect 150019 190979 150085 190980
rect 149835 188460 149901 188461
rect 149835 188396 149836 188460
rect 149900 188396 149901 188460
rect 149835 188395 149901 188396
rect 149838 79933 149898 188395
rect 150022 81157 150082 190979
rect 150294 187954 150914 198000
rect 151123 195260 151189 195261
rect 151123 195196 151124 195260
rect 151188 195196 151189 195260
rect 151123 195195 151189 195196
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 150939 139364 151005 139365
rect 150939 139300 150940 139364
rect 151004 139300 151005 139364
rect 150939 139299 151005 139300
rect 150019 81156 150085 81157
rect 150019 81092 150020 81156
rect 150084 81092 150085 81156
rect 150019 81091 150085 81092
rect 150203 80068 150269 80069
rect 150203 80004 150204 80068
rect 150268 80004 150269 80068
rect 150203 80003 150269 80004
rect 149835 79932 149901 79933
rect 149835 79868 149836 79932
rect 149900 79868 149901 79932
rect 149835 79867 149901 79868
rect 149651 79524 149717 79525
rect 149651 79460 149652 79524
rect 149716 79460 149717 79524
rect 149651 79459 149717 79460
rect 149838 79253 149898 79867
rect 149835 79252 149901 79253
rect 149835 79188 149836 79252
rect 149900 79188 149901 79252
rect 149835 79187 149901 79188
rect 150206 78573 150266 80003
rect 150942 79661 151002 139299
rect 151126 80205 151186 195195
rect 151123 80204 151189 80205
rect 151123 80140 151124 80204
rect 151188 80140 151189 80204
rect 151123 80139 151189 80140
rect 151123 80068 151189 80069
rect 151123 80004 151124 80068
rect 151188 80004 151189 80068
rect 151123 80003 151189 80004
rect 150939 79660 151005 79661
rect 150939 79596 150940 79660
rect 151004 79596 151005 79660
rect 150939 79595 151005 79596
rect 150203 78572 150269 78573
rect 150203 78508 150204 78572
rect 150268 78508 150269 78572
rect 150203 78507 150269 78508
rect 149283 72996 149349 72997
rect 149283 72932 149284 72996
rect 149348 72932 149349 72996
rect 149283 72931 149349 72932
rect 149835 72996 149901 72997
rect 149835 72932 149836 72996
rect 149900 72932 149901 72996
rect 149835 72931 149901 72932
rect 149099 71364 149165 71365
rect 149099 71300 149100 71364
rect 149164 71300 149165 71364
rect 149099 71299 149165 71300
rect 147811 70347 147877 70348
rect 147998 70350 148426 70410
rect 148550 70350 148794 70410
rect 147627 68236 147693 68237
rect 147627 68172 147628 68236
rect 147692 68172 147693 68236
rect 147627 68171 147693 68172
rect 147259 67284 147325 67285
rect 147259 67220 147260 67284
rect 147324 67220 147325 67284
rect 147259 67219 147325 67220
rect 147814 64890 147874 70347
rect 147998 67149 148058 70350
rect 147995 67148 148061 67149
rect 147995 67084 147996 67148
rect 148060 67084 148061 67148
rect 147995 67083 148061 67084
rect 147814 64830 148242 64890
rect 146891 55860 146957 55861
rect 146891 55796 146892 55860
rect 146956 55796 146957 55860
rect 146891 55795 146957 55796
rect 148182 46341 148242 64830
rect 148179 46340 148245 46341
rect 148179 46276 148180 46340
rect 148244 46276 148245 46340
rect 148179 46275 148245 46276
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 18596 145669 18597
rect 145603 18532 145604 18596
rect 145668 18532 145669 18596
rect 145603 18531 145669 18532
rect 144131 8940 144197 8941
rect 144131 8876 144132 8940
rect 144196 8876 144197 8940
rect 144131 8875 144197 8876
rect 145794 3454 146414 38898
rect 148550 7581 148610 70350
rect 149102 64890 149162 71299
rect 149102 64830 149714 64890
rect 149654 42125 149714 64830
rect 149838 56133 149898 72931
rect 149835 56132 149901 56133
rect 149835 56068 149836 56132
rect 149900 56068 149901 56132
rect 149835 56067 149901 56068
rect 150294 43954 150914 78000
rect 151126 71637 151186 80003
rect 151310 79797 151370 199819
rect 151491 195940 151557 195941
rect 151491 195876 151492 195940
rect 151556 195876 151557 195940
rect 151491 195875 151557 195876
rect 151307 79796 151373 79797
rect 151307 79732 151308 79796
rect 151372 79732 151373 79796
rect 151307 79731 151373 79732
rect 151494 79525 151554 195875
rect 152598 195125 152658 199819
rect 153518 199613 153578 200907
rect 158115 200836 158181 200837
rect 158115 200772 158116 200836
rect 158180 200772 158181 200836
rect 158115 200771 158181 200772
rect 156275 200700 156341 200701
rect 156275 200636 156276 200700
rect 156340 200636 156341 200700
rect 156275 200635 156341 200636
rect 153699 199884 153765 199885
rect 153699 199820 153700 199884
rect 153764 199820 153765 199884
rect 153699 199819 153765 199820
rect 154435 199884 154501 199885
rect 154435 199820 154436 199884
rect 154500 199820 154501 199884
rect 154435 199819 154501 199820
rect 155539 199884 155605 199885
rect 155539 199820 155540 199884
rect 155604 199820 155605 199884
rect 155539 199819 155605 199820
rect 155723 199884 155789 199885
rect 155723 199820 155724 199884
rect 155788 199882 155789 199884
rect 155788 199822 155970 199882
rect 155788 199820 155789 199822
rect 155723 199819 155789 199820
rect 153515 199612 153581 199613
rect 153515 199548 153516 199612
rect 153580 199548 153581 199612
rect 153515 199547 153581 199548
rect 153702 198525 153762 199819
rect 153883 199612 153949 199613
rect 153883 199548 153884 199612
rect 153948 199548 153949 199612
rect 153883 199547 153949 199548
rect 153699 198524 153765 198525
rect 153699 198460 153700 198524
rect 153764 198460 153765 198524
rect 153699 198459 153765 198460
rect 153886 195938 153946 199547
rect 154067 197300 154133 197301
rect 154067 197236 154068 197300
rect 154132 197236 154133 197300
rect 154067 197235 154133 197236
rect 153702 195878 153946 195938
rect 153515 195260 153581 195261
rect 153515 195196 153516 195260
rect 153580 195196 153581 195260
rect 153515 195195 153581 195196
rect 152595 195124 152661 195125
rect 152595 195060 152596 195124
rect 152660 195060 152661 195124
rect 152595 195059 152661 195060
rect 152227 194172 152293 194173
rect 152227 194108 152228 194172
rect 152292 194108 152293 194172
rect 152227 194107 152293 194108
rect 151859 191588 151925 191589
rect 151859 191524 151860 191588
rect 151924 191524 151925 191588
rect 151859 191523 151925 191524
rect 151675 80068 151741 80069
rect 151675 80004 151676 80068
rect 151740 80004 151741 80068
rect 151675 80003 151741 80004
rect 151491 79524 151557 79525
rect 151491 79460 151492 79524
rect 151556 79460 151557 79524
rect 151491 79459 151557 79460
rect 151491 78572 151557 78573
rect 151491 78508 151492 78572
rect 151556 78508 151557 78572
rect 151491 78507 151557 78508
rect 151123 71636 151189 71637
rect 151123 71572 151124 71636
rect 151188 71572 151189 71636
rect 151123 71571 151189 71572
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 149651 42124 149717 42125
rect 149651 42060 149652 42124
rect 149716 42060 149717 42124
rect 149651 42059 149717 42060
rect 150294 7954 150914 43398
rect 151126 29613 151186 71571
rect 151494 61981 151554 78507
rect 151491 61980 151557 61981
rect 151491 61916 151492 61980
rect 151556 61916 151557 61980
rect 151491 61915 151557 61916
rect 151678 58989 151738 80003
rect 151862 79797 151922 191523
rect 151859 79796 151925 79797
rect 151859 79732 151860 79796
rect 151924 79732 151925 79796
rect 151859 79731 151925 79732
rect 152230 79525 152290 194107
rect 152595 188868 152661 188869
rect 152595 188804 152596 188868
rect 152660 188804 152661 188868
rect 152595 188803 152661 188804
rect 152411 79932 152477 79933
rect 152411 79868 152412 79932
rect 152476 79868 152477 79932
rect 152411 79867 152477 79868
rect 152227 79524 152293 79525
rect 152227 79460 152228 79524
rect 152292 79460 152293 79524
rect 152227 79459 152293 79460
rect 152414 76258 152474 79867
rect 152598 79661 152658 188803
rect 152779 187372 152845 187373
rect 152779 187308 152780 187372
rect 152844 187308 152845 187372
rect 152779 187307 152845 187308
rect 152782 79933 152842 187307
rect 152779 79932 152845 79933
rect 152779 79868 152780 79932
rect 152844 79868 152845 79932
rect 152779 79867 152845 79868
rect 152595 79660 152661 79661
rect 152595 79596 152596 79660
rect 152660 79596 152661 79660
rect 152595 79595 152661 79596
rect 153518 79525 153578 195195
rect 153702 79525 153762 195878
rect 153883 195532 153949 195533
rect 153883 195468 153884 195532
rect 153948 195468 153949 195532
rect 153883 195467 153949 195468
rect 153886 79797 153946 195467
rect 154070 82830 154130 197235
rect 154438 195261 154498 199819
rect 154619 199476 154685 199477
rect 154619 199412 154620 199476
rect 154684 199412 154685 199476
rect 154619 199411 154685 199412
rect 154435 195260 154501 195261
rect 154435 195196 154436 195260
rect 154500 195196 154501 195260
rect 154435 195195 154501 195196
rect 154070 82770 154314 82830
rect 154254 79933 154314 82770
rect 154251 79932 154317 79933
rect 154251 79868 154252 79932
rect 154316 79868 154317 79932
rect 154251 79867 154317 79868
rect 153883 79796 153949 79797
rect 153883 79732 153884 79796
rect 153948 79732 153949 79796
rect 153883 79731 153949 79732
rect 153515 79524 153581 79525
rect 153515 79460 153516 79524
rect 153580 79460 153581 79524
rect 153515 79459 153581 79460
rect 153699 79524 153765 79525
rect 153699 79460 153700 79524
rect 153764 79460 153765 79524
rect 153699 79459 153765 79460
rect 154067 78708 154133 78709
rect 154067 78644 154068 78708
rect 154132 78644 154133 78708
rect 154067 78643 154133 78644
rect 153699 77892 153765 77893
rect 153699 77828 153700 77892
rect 153764 77828 153765 77892
rect 153699 77827 153765 77828
rect 152963 76804 153029 76805
rect 152963 76740 152964 76804
rect 153028 76740 153029 76804
rect 152963 76739 153029 76740
rect 152414 76198 152842 76258
rect 152595 75988 152661 75989
rect 152595 75924 152596 75988
rect 152660 75924 152661 75988
rect 152595 75923 152661 75924
rect 152411 74628 152477 74629
rect 152411 74564 152412 74628
rect 152476 74564 152477 74628
rect 152411 74563 152477 74564
rect 152414 71501 152474 74563
rect 152411 71500 152477 71501
rect 152411 71436 152412 71500
rect 152476 71436 152477 71500
rect 152411 71435 152477 71436
rect 151675 58988 151741 58989
rect 151675 58924 151676 58988
rect 151740 58924 151741 58988
rect 151675 58923 151741 58924
rect 151123 29612 151189 29613
rect 151123 29548 151124 29612
rect 151188 29548 151189 29612
rect 151123 29547 151189 29548
rect 152414 13021 152474 71435
rect 152598 64837 152658 75923
rect 152595 64836 152661 64837
rect 152595 64772 152596 64836
rect 152660 64772 152661 64836
rect 152595 64771 152661 64772
rect 152782 63477 152842 76198
rect 152779 63476 152845 63477
rect 152779 63412 152780 63476
rect 152844 63412 152845 63476
rect 152779 63411 152845 63412
rect 152966 60621 153026 76739
rect 153702 70277 153762 77827
rect 153699 70276 153765 70277
rect 153699 70212 153700 70276
rect 153764 70212 153765 70276
rect 153699 70211 153765 70212
rect 152963 60620 153029 60621
rect 152963 60556 152964 60620
rect 153028 60556 153029 60620
rect 152963 60555 153029 60556
rect 153702 26893 153762 70211
rect 154070 59125 154130 78643
rect 154254 78165 154314 79867
rect 154622 79253 154682 199411
rect 154794 192454 155414 198000
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 154803 139364 154869 139365
rect 154803 139300 154804 139364
rect 154868 139300 154869 139364
rect 154803 139299 154869 139300
rect 155355 139364 155421 139365
rect 155355 139300 155356 139364
rect 155420 139300 155421 139364
rect 155355 139299 155421 139300
rect 154806 79661 154866 139299
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 155358 80069 155418 139299
rect 155355 80068 155421 80069
rect 155355 80004 155356 80068
rect 155420 80004 155421 80068
rect 155355 80003 155421 80004
rect 155355 79932 155421 79933
rect 155355 79868 155356 79932
rect 155420 79868 155421 79932
rect 155355 79867 155421 79868
rect 154803 79660 154869 79661
rect 154803 79596 154804 79660
rect 154868 79596 154869 79660
rect 154803 79595 154869 79596
rect 154619 79252 154685 79253
rect 154619 79188 154620 79252
rect 154684 79188 154685 79252
rect 155358 79250 155418 79867
rect 155542 79797 155602 199819
rect 155723 199748 155789 199749
rect 155723 199684 155724 199748
rect 155788 199684 155789 199748
rect 155723 199683 155789 199684
rect 155726 189957 155786 199683
rect 155910 198797 155970 199822
rect 156278 199477 156338 200635
rect 156827 199884 156893 199885
rect 156827 199820 156828 199884
rect 156892 199820 156893 199884
rect 156827 199819 156893 199820
rect 157931 199884 157997 199885
rect 157931 199820 157932 199884
rect 157996 199820 157997 199884
rect 157931 199819 157997 199820
rect 156275 199476 156341 199477
rect 156275 199412 156276 199476
rect 156340 199412 156341 199476
rect 156275 199411 156341 199412
rect 156459 199476 156525 199477
rect 156459 199412 156460 199476
rect 156524 199412 156525 199476
rect 156459 199411 156525 199412
rect 155907 198796 155973 198797
rect 155907 198732 155908 198796
rect 155972 198732 155973 198796
rect 155907 198731 155973 198732
rect 156275 198388 156341 198389
rect 156275 198324 156276 198388
rect 156340 198324 156341 198388
rect 156275 198323 156341 198324
rect 156091 195940 156157 195941
rect 156091 195876 156092 195940
rect 156156 195876 156157 195940
rect 156091 195875 156157 195876
rect 156094 191181 156154 195875
rect 156091 191180 156157 191181
rect 156091 191116 156092 191180
rect 156156 191116 156157 191180
rect 156091 191115 156157 191116
rect 155723 189956 155789 189957
rect 155723 189892 155724 189956
rect 155788 189892 155789 189956
rect 155723 189891 155789 189892
rect 155539 79796 155605 79797
rect 155539 79732 155540 79796
rect 155604 79732 155605 79796
rect 155539 79731 155605 79732
rect 155723 79796 155789 79797
rect 155723 79732 155724 79796
rect 155788 79732 155789 79796
rect 155723 79731 155789 79732
rect 155542 79389 155602 79731
rect 155539 79388 155605 79389
rect 155539 79324 155540 79388
rect 155604 79324 155605 79388
rect 155539 79323 155605 79324
rect 155358 79190 155602 79250
rect 154619 79187 154685 79188
rect 154251 78164 154317 78165
rect 154251 78100 154252 78164
rect 154316 78100 154317 78164
rect 154251 78099 154317 78100
rect 154251 76668 154317 76669
rect 154251 76604 154252 76668
rect 154316 76604 154317 76668
rect 154251 76603 154317 76604
rect 154254 61845 154314 76603
rect 154251 61844 154317 61845
rect 154251 61780 154252 61844
rect 154316 61780 154317 61844
rect 154251 61779 154317 61780
rect 154067 59124 154133 59125
rect 154067 59060 154068 59124
rect 154132 59060 154133 59124
rect 154067 59059 154133 59060
rect 154794 48454 155414 78000
rect 155542 63205 155602 79190
rect 155539 63204 155605 63205
rect 155539 63140 155540 63204
rect 155604 63140 155605 63204
rect 155539 63139 155605 63140
rect 155726 60213 155786 79731
rect 156278 79661 156338 198323
rect 156462 80205 156522 199411
rect 156830 199341 156890 199819
rect 156827 199340 156893 199341
rect 156827 199276 156828 199340
rect 156892 199276 156893 199340
rect 156827 199275 156893 199276
rect 156643 197436 156709 197437
rect 156643 197372 156644 197436
rect 156708 197372 156709 197436
rect 156643 197371 156709 197372
rect 156459 80204 156525 80205
rect 156459 80140 156460 80204
rect 156524 80140 156525 80204
rect 156459 80139 156525 80140
rect 156459 79932 156525 79933
rect 156459 79868 156460 79932
rect 156524 79868 156525 79932
rect 156459 79867 156525 79868
rect 156275 79660 156341 79661
rect 156275 79596 156276 79660
rect 156340 79596 156341 79660
rect 156275 79595 156341 79596
rect 156462 78690 156522 79867
rect 156646 79117 156706 197371
rect 157011 189276 157077 189277
rect 157011 189212 157012 189276
rect 157076 189212 157077 189276
rect 157011 189211 157077 189212
rect 157014 99390 157074 189211
rect 157014 99330 157258 99390
rect 157198 80069 157258 99330
rect 157195 80068 157261 80069
rect 157195 80004 157196 80068
rect 157260 80004 157261 80068
rect 157195 80003 157261 80004
rect 157701 79932 157767 79933
rect 157701 79868 157702 79932
rect 157766 79930 157767 79932
rect 157766 79868 157810 79930
rect 157701 79867 157810 79868
rect 157011 79796 157077 79797
rect 157011 79732 157012 79796
rect 157076 79794 157077 79796
rect 157076 79734 157258 79794
rect 157076 79732 157077 79734
rect 157011 79731 157077 79732
rect 157011 79252 157077 79253
rect 157011 79188 157012 79252
rect 157076 79188 157077 79252
rect 157011 79187 157077 79188
rect 156643 79116 156709 79117
rect 156643 79052 156644 79116
rect 156708 79052 156709 79116
rect 156643 79051 156709 79052
rect 156462 78630 156890 78690
rect 156830 75986 156890 78630
rect 156646 75926 156890 75986
rect 156646 61709 156706 75926
rect 156827 75852 156893 75853
rect 156827 75788 156828 75852
rect 156892 75788 156893 75852
rect 156827 75787 156893 75788
rect 156643 61708 156709 61709
rect 156643 61644 156644 61708
rect 156708 61644 156709 61708
rect 156643 61643 156709 61644
rect 155723 60212 155789 60213
rect 155723 60148 155724 60212
rect 155788 60148 155789 60212
rect 155723 60147 155789 60148
rect 156830 57901 156890 75787
rect 156827 57900 156893 57901
rect 156827 57836 156828 57900
rect 156892 57836 156893 57900
rect 156827 57835 156893 57836
rect 157014 53821 157074 79187
rect 157011 53820 157077 53821
rect 157011 53756 157012 53820
rect 157076 53756 157077 53820
rect 157011 53755 157077 53756
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 153699 26892 153765 26893
rect 153699 26828 153700 26892
rect 153764 26828 153765 26892
rect 153699 26827 153765 26828
rect 152411 13020 152477 13021
rect 152411 12956 152412 13020
rect 152476 12956 152477 13020
rect 152411 12955 152477 12956
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 148547 7580 148613 7581
rect 148547 7516 148548 7580
rect 148612 7516 148613 7580
rect 148547 7515 148613 7516
rect 142659 3364 142725 3365
rect 142659 3300 142660 3364
rect 142724 3300 142725 3364
rect 142659 3299 142725 3300
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 47898
rect 157198 45389 157258 79734
rect 157750 78690 157810 79867
rect 157934 78845 157994 199819
rect 158118 199749 158178 200771
rect 168603 200292 168669 200293
rect 168603 200228 168604 200292
rect 168668 200228 168669 200292
rect 168603 200227 168669 200228
rect 161427 200156 161493 200157
rect 161427 200092 161428 200156
rect 161492 200092 161493 200156
rect 161427 200091 161493 200092
rect 158299 199884 158365 199885
rect 158299 199820 158300 199884
rect 158364 199820 158365 199884
rect 158299 199819 158365 199820
rect 158667 199884 158733 199885
rect 158667 199820 158668 199884
rect 158732 199820 158733 199884
rect 158667 199819 158733 199820
rect 160875 199884 160941 199885
rect 160875 199820 160876 199884
rect 160940 199820 160941 199884
rect 160875 199819 160941 199820
rect 158115 199748 158181 199749
rect 158115 199684 158116 199748
rect 158180 199684 158181 199748
rect 158115 199683 158181 199684
rect 158115 191180 158181 191181
rect 158115 191116 158116 191180
rect 158180 191116 158181 191180
rect 158115 191115 158181 191116
rect 158118 79933 158178 191115
rect 158115 79932 158181 79933
rect 158115 79868 158116 79932
rect 158180 79868 158181 79932
rect 158115 79867 158181 79868
rect 158118 79658 158178 79867
rect 158302 79797 158362 199819
rect 158670 196077 158730 199819
rect 159035 199748 159101 199749
rect 159035 199684 159036 199748
rect 159100 199684 159101 199748
rect 159035 199683 159101 199684
rect 159771 199748 159837 199749
rect 159771 199684 159772 199748
rect 159836 199684 159837 199748
rect 159771 199683 159837 199684
rect 160323 199748 160389 199749
rect 160323 199684 160324 199748
rect 160388 199684 160389 199748
rect 160323 199683 160389 199684
rect 158851 199476 158917 199477
rect 158851 199412 158852 199476
rect 158916 199412 158917 199476
rect 158851 199411 158917 199412
rect 158667 196076 158733 196077
rect 158667 196012 158668 196076
rect 158732 196012 158733 196076
rect 158667 196011 158733 196012
rect 158483 194036 158549 194037
rect 158483 193972 158484 194036
rect 158548 193972 158549 194036
rect 158483 193971 158549 193972
rect 158299 79796 158365 79797
rect 158299 79732 158300 79796
rect 158364 79732 158365 79796
rect 158299 79731 158365 79732
rect 158486 79661 158546 193971
rect 158667 81156 158733 81157
rect 158667 81092 158668 81156
rect 158732 81092 158733 81156
rect 158667 81091 158733 81092
rect 158483 79660 158549 79661
rect 158118 79598 158362 79658
rect 158115 79524 158181 79525
rect 158115 79460 158116 79524
rect 158180 79460 158181 79524
rect 158115 79459 158181 79460
rect 157931 78844 157997 78845
rect 157931 78780 157932 78844
rect 157996 78780 157997 78844
rect 157931 78779 157997 78780
rect 157750 78630 157994 78690
rect 157934 73813 157994 78630
rect 157931 73812 157997 73813
rect 157931 73748 157932 73812
rect 157996 73748 157997 73812
rect 157931 73747 157997 73748
rect 158118 60485 158178 79459
rect 158302 79389 158362 79598
rect 158483 79596 158484 79660
rect 158548 79596 158549 79660
rect 158483 79595 158549 79596
rect 158299 79388 158365 79389
rect 158299 79324 158300 79388
rect 158364 79324 158365 79388
rect 158299 79323 158365 79324
rect 158299 79252 158365 79253
rect 158299 79188 158300 79252
rect 158364 79188 158365 79252
rect 158299 79187 158365 79188
rect 158115 60484 158181 60485
rect 158115 60420 158116 60484
rect 158180 60420 158181 60484
rect 158115 60419 158181 60420
rect 158302 58717 158362 79187
rect 158486 78165 158546 79595
rect 158670 78981 158730 81091
rect 158854 79933 158914 199411
rect 158851 79932 158917 79933
rect 158851 79868 158852 79932
rect 158916 79868 158917 79932
rect 158851 79867 158917 79868
rect 159038 79525 159098 199683
rect 159774 198389 159834 199683
rect 159771 198388 159837 198389
rect 159771 198324 159772 198388
rect 159836 198324 159837 198388
rect 159771 198323 159837 198324
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 160326 195941 160386 199683
rect 160323 195940 160389 195941
rect 160323 195876 160324 195940
rect 160388 195876 160389 195940
rect 160323 195875 160389 195876
rect 160878 191450 160938 199819
rect 161430 199477 161490 200091
rect 165659 200020 165725 200021
rect 165659 199956 165660 200020
rect 165724 199956 165725 200020
rect 165659 199955 165725 199956
rect 163083 199884 163149 199885
rect 163083 199820 163084 199884
rect 163148 199820 163149 199884
rect 163083 199819 163149 199820
rect 163267 199884 163333 199885
rect 163267 199820 163268 199884
rect 163332 199820 163333 199884
rect 163267 199819 163333 199820
rect 164371 199884 164437 199885
rect 164371 199820 164372 199884
rect 164436 199820 164437 199884
rect 164371 199819 164437 199820
rect 164555 199884 164621 199885
rect 164555 199820 164556 199884
rect 164620 199820 164621 199884
rect 164555 199819 164621 199820
rect 162899 199748 162965 199749
rect 162899 199684 162900 199748
rect 162964 199684 162965 199748
rect 162899 199683 162965 199684
rect 162902 199477 162962 199683
rect 161427 199476 161493 199477
rect 161427 199412 161428 199476
rect 161492 199412 161493 199476
rect 161427 199411 161493 199412
rect 162899 199476 162965 199477
rect 162899 199412 162900 199476
rect 162964 199412 162965 199476
rect 162899 199411 162965 199412
rect 161243 197028 161309 197029
rect 161243 196964 161244 197028
rect 161308 196964 161309 197028
rect 161243 196963 161309 196964
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 160694 191390 160938 191450
rect 159219 139364 159285 139365
rect 159219 139300 159220 139364
rect 159284 139300 159285 139364
rect 159219 139299 159285 139300
rect 159955 139364 160021 139365
rect 159955 139300 159956 139364
rect 160020 139300 160021 139364
rect 159955 139299 160021 139300
rect 159222 89730 159282 139299
rect 159222 89670 159650 89730
rect 159403 81020 159469 81021
rect 159403 80956 159404 81020
rect 159468 80956 159469 81020
rect 159403 80955 159469 80956
rect 159219 80068 159285 80069
rect 159219 80004 159220 80068
rect 159284 80004 159285 80068
rect 159219 80003 159285 80004
rect 159035 79524 159101 79525
rect 159035 79460 159036 79524
rect 159100 79460 159101 79524
rect 159035 79459 159101 79460
rect 158667 78980 158733 78981
rect 158667 78916 158668 78980
rect 158732 78916 158733 78980
rect 158667 78915 158733 78916
rect 158667 78572 158733 78573
rect 158667 78508 158668 78572
rect 158732 78508 158733 78572
rect 158667 78507 158733 78508
rect 158483 78164 158549 78165
rect 158483 78100 158484 78164
rect 158548 78100 158549 78164
rect 158483 78099 158549 78100
rect 158670 72725 158730 78507
rect 159222 78162 159282 80003
rect 159406 79117 159466 80955
rect 159590 79797 159650 89670
rect 159587 79796 159653 79797
rect 159587 79732 159588 79796
rect 159652 79732 159653 79796
rect 159587 79731 159653 79732
rect 159403 79116 159469 79117
rect 159403 79052 159404 79116
rect 159468 79052 159469 79116
rect 159403 79051 159469 79052
rect 159958 78709 160018 139299
rect 160507 80340 160573 80341
rect 160507 80276 160508 80340
rect 160572 80276 160573 80340
rect 160507 80275 160573 80276
rect 160510 79525 160570 80275
rect 160694 79797 160754 191390
rect 161059 191180 161125 191181
rect 161059 191116 161060 191180
rect 161124 191116 161125 191180
rect 161059 191115 161125 191116
rect 160875 191044 160941 191045
rect 160875 190980 160876 191044
rect 160940 190980 160941 191044
rect 160875 190979 160941 190980
rect 160691 79796 160757 79797
rect 160691 79732 160692 79796
rect 160756 79732 160757 79796
rect 160691 79731 160757 79732
rect 160507 79524 160573 79525
rect 160507 79460 160508 79524
rect 160572 79460 160573 79524
rect 160507 79459 160573 79460
rect 159955 78708 160021 78709
rect 159955 78644 159956 78708
rect 160020 78644 160021 78708
rect 159955 78643 160021 78644
rect 160694 78437 160754 79731
rect 160691 78436 160757 78437
rect 160691 78372 160692 78436
rect 160756 78372 160757 78436
rect 160691 78371 160757 78372
rect 160878 78301 160938 190979
rect 161062 80069 161122 191115
rect 161059 80068 161125 80069
rect 161059 80004 161060 80068
rect 161124 80004 161125 80068
rect 161059 80003 161125 80004
rect 161062 79525 161122 80003
rect 161059 79524 161125 79525
rect 161059 79460 161060 79524
rect 161124 79460 161125 79524
rect 161059 79459 161125 79460
rect 161246 79117 161306 196963
rect 163086 196893 163146 199819
rect 163270 199477 163330 199819
rect 163819 199748 163885 199749
rect 163819 199684 163820 199748
rect 163884 199684 163885 199748
rect 163819 199683 163885 199684
rect 163267 199476 163333 199477
rect 163267 199412 163268 199476
rect 163332 199412 163333 199476
rect 163267 199411 163333 199412
rect 163635 198252 163701 198253
rect 163635 198188 163636 198252
rect 163700 198188 163701 198252
rect 163635 198187 163701 198188
rect 163083 196892 163149 196893
rect 163083 196828 163084 196892
rect 163148 196828 163149 196892
rect 163083 196827 163149 196828
rect 162715 195940 162781 195941
rect 162715 195876 162716 195940
rect 162780 195876 162781 195940
rect 162715 195875 162781 195876
rect 162163 191180 162229 191181
rect 162163 191116 162164 191180
rect 162228 191116 162229 191180
rect 162163 191115 162229 191116
rect 161979 187508 162045 187509
rect 161979 187444 161980 187508
rect 162044 187444 162045 187508
rect 161979 187443 162045 187444
rect 161611 79796 161677 79797
rect 161611 79732 161612 79796
rect 161676 79732 161677 79796
rect 161611 79731 161677 79732
rect 161243 79116 161309 79117
rect 161243 79052 161244 79116
rect 161308 79052 161309 79116
rect 161243 79051 161309 79052
rect 161614 78706 161674 79731
rect 161982 79661 162042 187443
rect 162166 79930 162226 191115
rect 162347 154460 162413 154461
rect 162347 154396 162348 154460
rect 162412 154396 162413 154460
rect 162347 154395 162413 154396
rect 162350 93870 162410 154395
rect 162350 93810 162594 93870
rect 162534 80885 162594 93810
rect 162531 80884 162597 80885
rect 162531 80820 162532 80884
rect 162596 80820 162597 80884
rect 162531 80819 162597 80820
rect 162718 80477 162778 195875
rect 162899 195260 162965 195261
rect 162899 195196 162900 195260
rect 162964 195196 162965 195260
rect 162899 195195 162965 195196
rect 162715 80476 162781 80477
rect 162715 80412 162716 80476
rect 162780 80412 162781 80476
rect 162715 80411 162781 80412
rect 162347 79932 162413 79933
rect 162347 79930 162348 79932
rect 162166 79870 162348 79930
rect 162347 79868 162348 79870
rect 162412 79868 162413 79932
rect 162347 79867 162413 79868
rect 161979 79660 162045 79661
rect 161979 79596 161980 79660
rect 162044 79596 162045 79660
rect 161979 79595 162045 79596
rect 162163 79388 162229 79389
rect 162163 79324 162164 79388
rect 162228 79324 162229 79388
rect 162163 79323 162229 79324
rect 161062 78646 161674 78706
rect 160875 78300 160941 78301
rect 160875 78236 160876 78300
rect 160940 78236 160941 78300
rect 160875 78235 160941 78236
rect 158854 78102 159282 78162
rect 158667 72724 158733 72725
rect 158667 72660 158668 72724
rect 158732 72660 158733 72724
rect 158667 72659 158733 72660
rect 158670 70410 158730 72659
rect 158486 70350 158730 70410
rect 158299 58716 158365 58717
rect 158299 58652 158300 58716
rect 158364 58652 158365 58716
rect 158299 58651 158365 58652
rect 157195 45388 157261 45389
rect 157195 45324 157196 45388
rect 157260 45324 157261 45388
rect 157195 45323 157261 45324
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 158486 6221 158546 70350
rect 158854 53549 158914 78102
rect 159035 75988 159101 75989
rect 159035 75924 159036 75988
rect 159100 75924 159101 75988
rect 159035 75923 159101 75924
rect 158851 53548 158917 53549
rect 158851 53484 158852 53548
rect 158916 53484 158917 53548
rect 158851 53483 158917 53484
rect 159038 50693 159098 75923
rect 159294 52954 159914 78000
rect 160875 75988 160941 75989
rect 160875 75924 160876 75988
rect 160940 75924 160941 75988
rect 160875 75923 160941 75924
rect 160691 75716 160757 75717
rect 160691 75652 160692 75716
rect 160756 75652 160757 75716
rect 160691 75651 160757 75652
rect 160694 59261 160754 75651
rect 160691 59260 160757 59261
rect 160691 59196 160692 59260
rect 160756 59196 160757 59260
rect 160691 59195 160757 59196
rect 160878 55181 160938 75923
rect 160875 55180 160941 55181
rect 160875 55116 160876 55180
rect 160940 55116 160941 55180
rect 160875 55115 160941 55116
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 50692 159101 50693
rect 159035 50628 159036 50692
rect 159100 50628 159101 50692
rect 159035 50627 159101 50628
rect 159294 16954 159914 52398
rect 161062 52189 161122 78646
rect 161243 78572 161309 78573
rect 161243 78508 161244 78572
rect 161308 78508 161309 78572
rect 161243 78507 161309 78508
rect 161246 52325 161306 78507
rect 162166 67650 162226 79323
rect 162350 76941 162410 79867
rect 162902 79389 162962 195195
rect 163267 187372 163333 187373
rect 163267 187308 163268 187372
rect 163332 187308 163333 187372
rect 163267 187307 163333 187308
rect 163270 79525 163330 187307
rect 163638 80069 163698 198187
rect 163635 80068 163701 80069
rect 163635 80004 163636 80068
rect 163700 80004 163701 80068
rect 163635 80003 163701 80004
rect 163451 79796 163517 79797
rect 163451 79732 163452 79796
rect 163516 79732 163517 79796
rect 163451 79731 163517 79732
rect 163267 79524 163333 79525
rect 163267 79460 163268 79524
rect 163332 79460 163333 79524
rect 163267 79459 163333 79460
rect 162899 79388 162965 79389
rect 162899 79324 162900 79388
rect 162964 79324 162965 79388
rect 162899 79323 162965 79324
rect 162715 77620 162781 77621
rect 162715 77556 162716 77620
rect 162780 77556 162781 77620
rect 162715 77555 162781 77556
rect 162531 77076 162597 77077
rect 162531 77012 162532 77076
rect 162596 77012 162597 77076
rect 162531 77011 162597 77012
rect 162347 76940 162413 76941
rect 162347 76876 162348 76940
rect 162412 76876 162413 76940
rect 162347 76875 162413 76876
rect 162166 67590 162410 67650
rect 162350 56541 162410 67590
rect 162347 56540 162413 56541
rect 162347 56476 162348 56540
rect 162412 56476 162413 56540
rect 162347 56475 162413 56476
rect 162534 53685 162594 77011
rect 162531 53684 162597 53685
rect 162531 53620 162532 53684
rect 162596 53620 162597 53684
rect 162531 53619 162597 53620
rect 161243 52324 161309 52325
rect 161243 52260 161244 52324
rect 161308 52260 161309 52324
rect 161243 52259 161309 52260
rect 161059 52188 161125 52189
rect 161059 52124 161060 52188
rect 161124 52124 161125 52188
rect 161059 52123 161125 52124
rect 162718 50829 162778 77555
rect 163270 77213 163330 79459
rect 163267 77212 163333 77213
rect 163267 77148 163268 77212
rect 163332 77148 163333 77212
rect 163267 77147 163333 77148
rect 163267 73676 163333 73677
rect 163267 73612 163268 73676
rect 163332 73612 163333 73676
rect 163267 73611 163333 73612
rect 163270 52461 163330 73611
rect 163267 52460 163333 52461
rect 163267 52396 163268 52460
rect 163332 52396 163333 52460
rect 163267 52395 163333 52396
rect 162715 50828 162781 50829
rect 162715 50764 162716 50828
rect 162780 50764 162781 50828
rect 162715 50763 162781 50764
rect 163454 49469 163514 79731
rect 163822 78981 163882 199683
rect 164374 195125 164434 199819
rect 164371 195124 164437 195125
rect 164371 195060 164372 195124
rect 164436 195060 164437 195124
rect 164371 195059 164437 195060
rect 164558 194989 164618 199819
rect 164739 195260 164805 195261
rect 164739 195196 164740 195260
rect 164804 195196 164805 195260
rect 164739 195195 164805 195196
rect 164555 194988 164621 194989
rect 164555 194924 164556 194988
rect 164620 194924 164621 194988
rect 164555 194923 164621 194924
rect 164742 86970 164802 195195
rect 165662 194989 165722 199955
rect 168606 199885 168666 200227
rect 169891 200156 169957 200157
rect 169891 200092 169892 200156
rect 169956 200092 169957 200156
rect 169891 200091 169957 200092
rect 165843 199884 165909 199885
rect 165843 199820 165844 199884
rect 165908 199820 165909 199884
rect 165843 199819 165909 199820
rect 166579 199884 166645 199885
rect 166579 199820 166580 199884
rect 166644 199820 166645 199884
rect 166579 199819 166645 199820
rect 168603 199884 168669 199885
rect 168603 199820 168604 199884
rect 168668 199820 168669 199884
rect 168603 199819 168669 199820
rect 168787 199884 168853 199885
rect 168787 199820 168788 199884
rect 168852 199820 168853 199884
rect 168787 199819 168853 199820
rect 165846 197165 165906 199819
rect 166027 197300 166093 197301
rect 166027 197236 166028 197300
rect 166092 197236 166093 197300
rect 166027 197235 166093 197236
rect 165843 197164 165909 197165
rect 165843 197100 165844 197164
rect 165908 197100 165909 197164
rect 165843 197099 165909 197100
rect 165659 194988 165725 194989
rect 165659 194924 165660 194988
rect 165724 194924 165725 194988
rect 165659 194923 165725 194924
rect 165843 191180 165909 191181
rect 165843 191116 165844 191180
rect 165908 191116 165909 191180
rect 165843 191115 165909 191116
rect 165107 188596 165173 188597
rect 165107 188532 165108 188596
rect 165172 188532 165173 188596
rect 165107 188531 165173 188532
rect 164923 182612 164989 182613
rect 164923 182548 164924 182612
rect 164988 182548 164989 182612
rect 164923 182547 164989 182548
rect 164558 86910 164802 86970
rect 164003 79932 164069 79933
rect 164003 79868 164004 79932
rect 164068 79868 164069 79932
rect 164003 79867 164069 79868
rect 163819 78980 163885 78981
rect 163819 78916 163820 78980
rect 163884 78916 163885 78980
rect 163819 78915 163885 78916
rect 163822 78573 163882 78915
rect 163819 78572 163885 78573
rect 163819 78508 163820 78572
rect 163884 78508 163885 78572
rect 163819 78507 163885 78508
rect 164006 78434 164066 79867
rect 164558 79389 164618 86910
rect 164739 79796 164805 79797
rect 164739 79732 164740 79796
rect 164804 79732 164805 79796
rect 164739 79731 164805 79732
rect 164555 79388 164621 79389
rect 164555 79324 164556 79388
rect 164620 79324 164621 79388
rect 164555 79323 164621 79324
rect 163638 78374 164066 78434
rect 163451 49468 163517 49469
rect 163451 49404 163452 49468
rect 163516 49404 163517 49468
rect 163451 49403 163517 49404
rect 163638 48109 163698 78374
rect 164742 78162 164802 79731
rect 164926 79253 164986 182547
rect 165110 79933 165170 188531
rect 165291 185876 165357 185877
rect 165291 185812 165292 185876
rect 165356 185812 165357 185876
rect 165291 185811 165357 185812
rect 165294 79933 165354 185811
rect 165107 79932 165173 79933
rect 165107 79868 165108 79932
rect 165172 79868 165173 79932
rect 165107 79867 165173 79868
rect 165291 79932 165357 79933
rect 165291 79868 165292 79932
rect 165356 79868 165357 79932
rect 165291 79867 165357 79868
rect 164923 79252 164989 79253
rect 164923 79188 164924 79252
rect 164988 79188 164989 79252
rect 164923 79187 164989 79188
rect 165294 78437 165354 79867
rect 165846 79389 165906 191115
rect 166030 79933 166090 197235
rect 166582 195261 166642 199819
rect 166763 199748 166829 199749
rect 166763 199684 166764 199748
rect 166828 199684 166829 199748
rect 166763 199683 166829 199684
rect 167867 199748 167933 199749
rect 167867 199684 167868 199748
rect 167932 199684 167933 199748
rect 167867 199683 167933 199684
rect 166579 195260 166645 195261
rect 166579 195196 166580 195260
rect 166644 195196 166645 195260
rect 166579 195195 166645 195196
rect 166211 190092 166277 190093
rect 166211 190028 166212 190092
rect 166276 190028 166277 190092
rect 166211 190027 166277 190028
rect 166027 79932 166093 79933
rect 166027 79868 166028 79932
rect 166092 79868 166093 79932
rect 166027 79867 166093 79868
rect 165843 79388 165909 79389
rect 165843 79324 165844 79388
rect 165908 79324 165909 79388
rect 165843 79323 165909 79324
rect 166214 79253 166274 190027
rect 166766 85590 166826 199683
rect 167499 198660 167565 198661
rect 167499 198596 167500 198660
rect 167564 198596 167565 198660
rect 167499 198595 167565 198596
rect 166582 85530 166826 85590
rect 166582 79797 166642 85530
rect 167315 80204 167381 80205
rect 167315 80140 167316 80204
rect 167380 80140 167381 80204
rect 167315 80139 167381 80140
rect 166763 79932 166829 79933
rect 166763 79868 166764 79932
rect 166828 79868 166829 79932
rect 166763 79867 166829 79868
rect 166579 79796 166645 79797
rect 166579 79732 166580 79796
rect 166644 79732 166645 79796
rect 166579 79731 166645 79732
rect 166211 79252 166277 79253
rect 166211 79188 166212 79252
rect 166276 79188 166277 79252
rect 166211 79187 166277 79188
rect 166582 78845 166642 79731
rect 165475 78844 165541 78845
rect 165475 78780 165476 78844
rect 165540 78780 165541 78844
rect 165475 78779 165541 78780
rect 166579 78844 166645 78845
rect 166579 78780 166580 78844
rect 166644 78780 166645 78844
rect 166579 78779 166645 78780
rect 165291 78436 165357 78437
rect 165291 78372 165292 78436
rect 165356 78372 165357 78436
rect 165291 78371 165357 78372
rect 164742 78102 165170 78162
rect 164923 78028 164989 78029
rect 163794 57454 164414 78000
rect 164923 77964 164924 78028
rect 164988 77964 164989 78028
rect 164923 77963 164989 77964
rect 164926 67557 164986 77963
rect 164923 67556 164989 67557
rect 164923 67492 164924 67556
rect 164988 67492 164989 67556
rect 164923 67491 164989 67492
rect 165110 63341 165170 78102
rect 165291 73676 165357 73677
rect 165291 73612 165292 73676
rect 165356 73612 165357 73676
rect 165291 73611 165357 73612
rect 165107 63340 165173 63341
rect 165107 63276 165108 63340
rect 165172 63276 165173 63340
rect 165107 63275 165173 63276
rect 165294 57765 165354 73611
rect 165291 57764 165357 57765
rect 165291 57700 165292 57764
rect 165356 57700 165357 57764
rect 165291 57699 165357 57700
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 48108 163701 48109
rect 163635 48044 163636 48108
rect 163700 48044 163701 48108
rect 163635 48043 163701 48044
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 158483 6220 158549 6221
rect 158483 6156 158484 6220
rect 158548 6156 158549 6220
rect 158483 6155 158549 6156
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 56898
rect 165478 55045 165538 78779
rect 166395 78164 166461 78165
rect 166395 78100 166396 78164
rect 166460 78100 166461 78164
rect 166395 78099 166461 78100
rect 166211 75988 166277 75989
rect 166211 75924 166212 75988
rect 166276 75924 166277 75988
rect 166211 75923 166277 75924
rect 166214 62117 166274 75923
rect 166211 62116 166277 62117
rect 166211 62052 166212 62116
rect 166276 62052 166277 62116
rect 166211 62051 166277 62052
rect 165475 55044 165541 55045
rect 165475 54980 165476 55044
rect 165540 54980 165541 55044
rect 165475 54979 165541 54980
rect 166398 53277 166458 78099
rect 166579 78028 166645 78029
rect 166579 77964 166580 78028
rect 166644 77964 166645 78028
rect 166579 77963 166645 77964
rect 166395 53276 166461 53277
rect 166395 53212 166396 53276
rect 166460 53212 166461 53276
rect 166395 53211 166461 53212
rect 166582 50965 166642 77963
rect 166579 50964 166645 50965
rect 166579 50900 166580 50964
rect 166644 50900 166645 50964
rect 166579 50899 166645 50900
rect 166766 48245 166826 79867
rect 167318 76533 167378 80139
rect 167502 79933 167562 198595
rect 167683 195396 167749 195397
rect 167683 195332 167684 195396
rect 167748 195332 167749 195396
rect 167683 195331 167749 195332
rect 167686 80749 167746 195331
rect 167683 80748 167749 80749
rect 167683 80684 167684 80748
rect 167748 80684 167749 80748
rect 167683 80683 167749 80684
rect 167499 79932 167565 79933
rect 167499 79868 167500 79932
rect 167564 79868 167565 79932
rect 167499 79867 167565 79868
rect 167502 79661 167562 79867
rect 167499 79660 167565 79661
rect 167499 79596 167500 79660
rect 167564 79596 167565 79660
rect 167499 79595 167565 79596
rect 167686 79253 167746 80683
rect 167870 79661 167930 199683
rect 168051 195532 168117 195533
rect 168051 195468 168052 195532
rect 168116 195468 168117 195532
rect 168051 195467 168117 195468
rect 167867 79660 167933 79661
rect 167867 79596 167868 79660
rect 167932 79596 167933 79660
rect 167867 79595 167933 79596
rect 168054 79389 168114 195467
rect 168419 80884 168485 80885
rect 168419 80820 168420 80884
rect 168484 80820 168485 80884
rect 168419 80819 168485 80820
rect 168422 79933 168482 80819
rect 168419 79932 168485 79933
rect 168419 79868 168420 79932
rect 168484 79868 168485 79932
rect 168419 79867 168485 79868
rect 168790 79661 168850 199819
rect 169155 199748 169221 199749
rect 169155 199684 169156 199748
rect 169220 199684 169221 199748
rect 169155 199683 169221 199684
rect 169158 195533 169218 199683
rect 169523 199612 169589 199613
rect 169523 199548 169524 199612
rect 169588 199610 169589 199612
rect 169894 199610 169954 200091
rect 170811 200020 170877 200021
rect 170811 199956 170812 200020
rect 170876 199956 170877 200020
rect 170811 199955 170877 199956
rect 170443 199884 170509 199885
rect 170443 199820 170444 199884
rect 170508 199820 170509 199884
rect 170443 199819 170509 199820
rect 170075 199748 170141 199749
rect 170075 199684 170076 199748
rect 170140 199684 170141 199748
rect 170075 199683 170141 199684
rect 169588 199550 169954 199610
rect 169588 199548 169589 199550
rect 169523 199547 169589 199548
rect 169891 199476 169957 199477
rect 169891 199412 169892 199476
rect 169956 199412 169957 199476
rect 169891 199411 169957 199412
rect 169523 198116 169589 198117
rect 169523 198052 169524 198116
rect 169588 198052 169589 198116
rect 169523 198051 169589 198052
rect 169155 195532 169221 195533
rect 169155 195468 169156 195532
rect 169220 195468 169221 195532
rect 169155 195467 169221 195468
rect 169339 191180 169405 191181
rect 169339 191116 169340 191180
rect 169404 191116 169405 191180
rect 169339 191115 169405 191116
rect 168971 185876 169037 185877
rect 168971 185812 168972 185876
rect 169036 185812 169037 185876
rect 168971 185811 169037 185812
rect 168787 79660 168853 79661
rect 168787 79596 168788 79660
rect 168852 79596 168853 79660
rect 168787 79595 168853 79596
rect 168974 79389 169034 185811
rect 169155 79932 169221 79933
rect 169155 79868 169156 79932
rect 169220 79868 169221 79932
rect 169155 79867 169221 79868
rect 168051 79388 168117 79389
rect 168051 79324 168052 79388
rect 168116 79324 168117 79388
rect 168051 79323 168117 79324
rect 168971 79388 169037 79389
rect 168971 79324 168972 79388
rect 169036 79324 169037 79388
rect 168971 79323 169037 79324
rect 167683 79252 167749 79253
rect 167683 79188 167684 79252
rect 167748 79188 167749 79252
rect 167683 79187 167749 79188
rect 167315 76532 167381 76533
rect 167315 76468 167316 76532
rect 167380 76468 167381 76532
rect 167315 76467 167381 76468
rect 167315 76124 167381 76125
rect 167315 76060 167316 76124
rect 167380 76060 167381 76124
rect 167315 76059 167381 76060
rect 167318 67650 167378 76059
rect 167683 75988 167749 75989
rect 167683 75924 167684 75988
rect 167748 75924 167749 75988
rect 167683 75923 167749 75924
rect 167318 67590 167562 67650
rect 167502 49605 167562 67590
rect 167499 49604 167565 49605
rect 167499 49540 167500 49604
rect 167564 49540 167565 49604
rect 167499 49539 167565 49540
rect 166763 48244 166829 48245
rect 166763 48180 166764 48244
rect 166828 48180 166829 48244
rect 166763 48179 166829 48180
rect 167686 46885 167746 75923
rect 167867 75852 167933 75853
rect 167867 75788 167868 75852
rect 167932 75788 167933 75852
rect 167867 75787 167933 75788
rect 167683 46884 167749 46885
rect 167683 46820 167684 46884
rect 167748 46820 167749 46884
rect 167683 46819 167749 46820
rect 167870 45525 167930 75787
rect 168051 75716 168117 75717
rect 168051 75652 168052 75716
rect 168116 75652 168117 75716
rect 168051 75651 168117 75652
rect 167867 45524 167933 45525
rect 167867 45460 167868 45524
rect 167932 45460 167933 45524
rect 167867 45459 167933 45460
rect 168054 44165 168114 75651
rect 168294 61954 168914 78000
rect 169158 67650 169218 79867
rect 169342 79661 169402 191115
rect 169526 79797 169586 198051
rect 169707 80204 169773 80205
rect 169707 80140 169708 80204
rect 169772 80140 169773 80204
rect 169707 80139 169773 80140
rect 169523 79796 169589 79797
rect 169523 79732 169524 79796
rect 169588 79732 169589 79796
rect 169523 79731 169589 79732
rect 169339 79660 169405 79661
rect 169339 79596 169340 79660
rect 169404 79596 169405 79660
rect 169339 79595 169405 79596
rect 169710 70410 169770 80139
rect 169894 79797 169954 199411
rect 170078 81450 170138 199683
rect 170446 199477 170506 199819
rect 170814 199749 170874 199955
rect 170998 199749 171058 200907
rect 173755 200700 173821 200701
rect 173755 200636 173756 200700
rect 173820 200636 173821 200700
rect 173755 200635 173821 200636
rect 171363 199884 171429 199885
rect 171363 199820 171364 199884
rect 171428 199820 171429 199884
rect 171363 199819 171429 199820
rect 171915 199884 171981 199885
rect 171915 199820 171916 199884
rect 171980 199820 171981 199884
rect 171915 199819 171981 199820
rect 172099 199884 172165 199885
rect 172099 199820 172100 199884
rect 172164 199820 172165 199884
rect 172099 199819 172165 199820
rect 172651 199884 172717 199885
rect 172651 199820 172652 199884
rect 172716 199820 172717 199884
rect 172651 199819 172717 199820
rect 170811 199748 170877 199749
rect 170811 199684 170812 199748
rect 170876 199684 170877 199748
rect 170811 199683 170877 199684
rect 170995 199748 171061 199749
rect 170995 199684 170996 199748
rect 171060 199684 171061 199748
rect 170995 199683 171061 199684
rect 171366 199477 171426 199819
rect 170443 199476 170509 199477
rect 170443 199412 170444 199476
rect 170508 199412 170509 199476
rect 170443 199411 170509 199412
rect 170995 199476 171061 199477
rect 170995 199412 170996 199476
rect 171060 199412 171061 199476
rect 170995 199411 171061 199412
rect 171363 199476 171429 199477
rect 171363 199412 171364 199476
rect 171428 199412 171429 199476
rect 171363 199411 171429 199412
rect 170811 189276 170877 189277
rect 170811 189212 170812 189276
rect 170876 189212 170877 189276
rect 170811 189211 170877 189212
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 170078 81390 170322 81450
rect 170075 79932 170141 79933
rect 170075 79868 170076 79932
rect 170140 79868 170141 79932
rect 170075 79867 170141 79868
rect 169891 79796 169957 79797
rect 169891 79732 169892 79796
rect 169956 79732 169957 79796
rect 169891 79731 169957 79732
rect 170078 76125 170138 79867
rect 170262 79797 170322 81390
rect 170627 80884 170693 80885
rect 170627 80820 170628 80884
rect 170692 80820 170693 80884
rect 170627 80819 170693 80820
rect 170443 80204 170509 80205
rect 170443 80140 170444 80204
rect 170508 80140 170509 80204
rect 170443 80139 170509 80140
rect 170259 79796 170325 79797
rect 170259 79732 170260 79796
rect 170324 79732 170325 79796
rect 170259 79731 170325 79732
rect 170075 76124 170141 76125
rect 170075 76060 170076 76124
rect 170140 76060 170141 76124
rect 170075 76059 170141 76060
rect 169526 70350 169770 70410
rect 169158 67590 169402 67650
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168051 44164 168117 44165
rect 168051 44100 168052 44164
rect 168116 44100 168117 44164
rect 168051 44099 168117 44100
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 61398
rect 169342 49333 169402 67590
rect 169339 49332 169405 49333
rect 169339 49268 169340 49332
rect 169404 49268 169405 49332
rect 169339 49267 169405 49268
rect 169526 44029 169586 70350
rect 170262 66877 170322 79731
rect 170259 66876 170325 66877
rect 170259 66812 170260 66876
rect 170324 66812 170325 66876
rect 170259 66811 170325 66812
rect 170446 56405 170506 80139
rect 170630 79661 170690 80819
rect 170814 79933 170874 189211
rect 170811 79932 170877 79933
rect 170811 79868 170812 79932
rect 170876 79868 170877 79932
rect 170811 79867 170877 79868
rect 170627 79660 170693 79661
rect 170627 79596 170628 79660
rect 170692 79596 170693 79660
rect 170627 79595 170693 79596
rect 170814 79253 170874 79867
rect 170998 79253 171058 199411
rect 171918 198661 171978 199819
rect 171731 198660 171797 198661
rect 171731 198596 171732 198660
rect 171796 198596 171797 198660
rect 171731 198595 171797 198596
rect 171915 198660 171981 198661
rect 171915 198596 171916 198660
rect 171980 198596 171981 198660
rect 171915 198595 171981 198596
rect 171547 191180 171613 191181
rect 171547 191116 171548 191180
rect 171612 191116 171613 191180
rect 171547 191115 171613 191116
rect 171363 81156 171429 81157
rect 171363 81092 171364 81156
rect 171428 81092 171429 81156
rect 171363 81091 171429 81092
rect 171366 79389 171426 81091
rect 171550 79389 171610 191115
rect 171734 79933 171794 198595
rect 171915 198116 171981 198117
rect 171915 198052 171916 198116
rect 171980 198052 171981 198116
rect 171915 198051 171981 198052
rect 171731 79932 171797 79933
rect 171731 79868 171732 79932
rect 171796 79868 171797 79932
rect 171731 79867 171797 79868
rect 171731 79796 171797 79797
rect 171731 79732 171732 79796
rect 171796 79732 171797 79796
rect 171731 79731 171797 79732
rect 171363 79388 171429 79389
rect 171363 79324 171364 79388
rect 171428 79324 171429 79388
rect 171363 79323 171429 79324
rect 171547 79388 171613 79389
rect 171547 79324 171548 79388
rect 171612 79324 171613 79388
rect 171547 79323 171613 79324
rect 170811 79252 170877 79253
rect 170811 79188 170812 79252
rect 170876 79188 170877 79252
rect 170811 79187 170877 79188
rect 170995 79252 171061 79253
rect 170995 79188 170996 79252
rect 171060 79188 171061 79252
rect 170995 79187 171061 79188
rect 171550 78029 171610 79323
rect 171734 78709 171794 79731
rect 171918 79661 171978 198051
rect 172102 195533 172162 199819
rect 172283 199748 172349 199749
rect 172283 199684 172284 199748
rect 172348 199684 172349 199748
rect 172283 199683 172349 199684
rect 172099 195532 172165 195533
rect 172099 195468 172100 195532
rect 172164 195468 172165 195532
rect 172099 195467 172165 195468
rect 172286 182190 172346 199683
rect 172102 182130 172346 182190
rect 172102 79933 172162 182130
rect 172099 79932 172165 79933
rect 172099 79868 172100 79932
rect 172164 79868 172165 79932
rect 172099 79867 172165 79868
rect 171915 79660 171981 79661
rect 171915 79596 171916 79660
rect 171980 79596 171981 79660
rect 171915 79595 171981 79596
rect 171915 79252 171981 79253
rect 171915 79188 171916 79252
rect 171980 79188 171981 79252
rect 171915 79187 171981 79188
rect 171731 78708 171797 78709
rect 171731 78644 171732 78708
rect 171796 78644 171797 78708
rect 171731 78643 171797 78644
rect 171547 78028 171613 78029
rect 171547 77964 171548 78028
rect 171612 77964 171613 78028
rect 171547 77963 171613 77964
rect 171734 75989 171794 78643
rect 171731 75988 171797 75989
rect 171731 75924 171732 75988
rect 171796 75924 171797 75988
rect 171731 75923 171797 75924
rect 171918 66197 171978 79187
rect 172102 78709 172162 79867
rect 172654 79661 172714 199819
rect 173758 199477 173818 200635
rect 180747 200564 180813 200565
rect 180747 200500 180748 200564
rect 180812 200500 180813 200564
rect 180747 200499 180813 200500
rect 174310 200230 174554 200290
rect 173755 199476 173821 199477
rect 173755 199412 173756 199476
rect 173820 199412 173821 199476
rect 173755 199411 173821 199412
rect 174123 198116 174189 198117
rect 174123 198052 174124 198116
rect 174188 198052 174189 198116
rect 174123 198051 174189 198052
rect 173387 191316 173453 191317
rect 173387 191252 173388 191316
rect 173452 191252 173453 191316
rect 173387 191251 173453 191252
rect 173019 191180 173085 191181
rect 173019 191116 173020 191180
rect 173084 191116 173085 191180
rect 173019 191115 173085 191116
rect 172835 191044 172901 191045
rect 172835 190980 172836 191044
rect 172900 190980 172901 191044
rect 172835 190979 172901 190980
rect 172838 79797 172898 190979
rect 172835 79796 172901 79797
rect 172835 79732 172836 79796
rect 172900 79732 172901 79796
rect 172835 79731 172901 79732
rect 172651 79660 172717 79661
rect 172651 79596 172652 79660
rect 172716 79596 172717 79660
rect 172651 79595 172717 79596
rect 173022 79389 173082 191115
rect 173390 88350 173450 191251
rect 173206 88290 173450 88350
rect 173206 79389 173266 88290
rect 174126 81293 174186 198051
rect 174123 81292 174189 81293
rect 174123 81228 174124 81292
rect 174188 81228 174189 81292
rect 174123 81227 174189 81228
rect 174123 80068 174189 80069
rect 174123 80004 174124 80068
rect 174188 80004 174189 80068
rect 174123 80003 174189 80004
rect 173387 79932 173453 79933
rect 173387 79868 173388 79932
rect 173452 79868 173453 79932
rect 173387 79867 173453 79868
rect 173019 79388 173085 79389
rect 173019 79324 173020 79388
rect 173084 79324 173085 79388
rect 173019 79323 173085 79324
rect 173203 79388 173269 79389
rect 173203 79324 173204 79388
rect 173268 79324 173269 79388
rect 173203 79323 173269 79324
rect 172099 78708 172165 78709
rect 172099 78644 172100 78708
rect 172164 78644 172165 78708
rect 172099 78643 172165 78644
rect 173390 78301 173450 79867
rect 173571 79388 173637 79389
rect 173571 79324 173572 79388
rect 173636 79324 173637 79388
rect 173571 79323 173637 79324
rect 173387 78300 173453 78301
rect 173387 78236 173388 78300
rect 173452 78236 173453 78300
rect 173387 78235 173453 78236
rect 172099 75988 172165 75989
rect 172099 75924 172100 75988
rect 172164 75924 172165 75988
rect 172099 75923 172165 75924
rect 171915 66196 171981 66197
rect 171915 66132 171916 66196
rect 171980 66132 171981 66196
rect 171915 66131 171981 66132
rect 172102 64701 172162 75923
rect 172283 74356 172349 74357
rect 172283 74292 172284 74356
rect 172348 74292 172349 74356
rect 172283 74291 172349 74292
rect 172099 64700 172165 64701
rect 172099 64636 172100 64700
rect 172164 64636 172165 64700
rect 172099 64635 172165 64636
rect 172286 63069 172346 74291
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172283 63068 172349 63069
rect 172283 63004 172284 63068
rect 172348 63004 172349 63068
rect 172283 63003 172349 63004
rect 170443 56404 170509 56405
rect 170443 56340 170444 56404
rect 170508 56340 170509 56404
rect 170443 56339 170509 56340
rect 169523 44028 169589 44029
rect 169523 43964 169524 44028
rect 169588 43964 169589 44028
rect 169523 43963 169589 43964
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 173574 59941 173634 79323
rect 174126 76805 174186 80003
rect 174310 79797 174370 200230
rect 174494 199885 174554 200230
rect 178355 200020 178421 200021
rect 178355 199956 178356 200020
rect 178420 199956 178421 200020
rect 178355 199955 178421 199956
rect 174491 199884 174557 199885
rect 174491 199820 174492 199884
rect 174556 199820 174557 199884
rect 174491 199819 174557 199820
rect 176147 199884 176213 199885
rect 176147 199820 176148 199884
rect 176212 199820 176213 199884
rect 176147 199819 176213 199820
rect 174491 199748 174557 199749
rect 174491 199684 174492 199748
rect 174556 199684 174557 199748
rect 174491 199683 174557 199684
rect 175595 199748 175661 199749
rect 175595 199684 175596 199748
rect 175660 199684 175661 199748
rect 175595 199683 175661 199684
rect 174307 79796 174373 79797
rect 174307 79732 174308 79796
rect 174372 79732 174373 79796
rect 174307 79731 174373 79732
rect 174494 79661 174554 199683
rect 174675 196484 174741 196485
rect 174675 196420 174676 196484
rect 174740 196420 174741 196484
rect 174675 196419 174741 196420
rect 174491 79660 174557 79661
rect 174491 79596 174492 79660
rect 174556 79596 174557 79660
rect 174491 79595 174557 79596
rect 174678 79389 174738 196419
rect 175411 194852 175477 194853
rect 175411 194788 175412 194852
rect 175476 194788 175477 194852
rect 175411 194787 175477 194788
rect 174859 81292 174925 81293
rect 174859 81228 174860 81292
rect 174924 81228 174925 81292
rect 174859 81227 174925 81228
rect 174862 79933 174922 81227
rect 175227 80612 175293 80613
rect 175227 80548 175228 80612
rect 175292 80548 175293 80612
rect 175227 80547 175293 80548
rect 174859 79932 174925 79933
rect 174859 79868 174860 79932
rect 174924 79868 174925 79932
rect 174859 79867 174925 79868
rect 175230 79661 175290 80547
rect 175043 79660 175109 79661
rect 175043 79596 175044 79660
rect 175108 79596 175109 79660
rect 175043 79595 175109 79596
rect 175227 79660 175293 79661
rect 175227 79596 175228 79660
rect 175292 79596 175293 79660
rect 175227 79595 175293 79596
rect 174675 79388 174741 79389
rect 174675 79324 174676 79388
rect 174740 79324 174741 79388
rect 174675 79323 174741 79324
rect 174491 77076 174557 77077
rect 174491 77012 174492 77076
rect 174556 77012 174557 77076
rect 174491 77011 174557 77012
rect 174123 76804 174189 76805
rect 174123 76740 174124 76804
rect 174188 76740 174189 76804
rect 174123 76739 174189 76740
rect 173755 75172 173821 75173
rect 173755 75108 173756 75172
rect 173820 75108 173821 75172
rect 173755 75107 173821 75108
rect 173571 59940 173637 59941
rect 173571 59876 173572 59940
rect 173636 59876 173637 59940
rect 173571 59875 173637 59876
rect 173758 47973 173818 75107
rect 174494 57221 174554 77011
rect 175046 70410 175106 79595
rect 175414 79389 175474 194787
rect 175598 79933 175658 199683
rect 175779 191180 175845 191181
rect 175779 191116 175780 191180
rect 175844 191116 175845 191180
rect 175779 191115 175845 191116
rect 175782 93870 175842 191115
rect 176150 187781 176210 199819
rect 178171 199068 178237 199069
rect 178171 199004 178172 199068
rect 178236 199004 178237 199068
rect 178171 199003 178237 199004
rect 176515 188460 176581 188461
rect 176515 188396 176516 188460
rect 176580 188396 176581 188460
rect 176515 188395 176581 188396
rect 176883 188460 176949 188461
rect 176883 188396 176884 188460
rect 176948 188396 176949 188460
rect 176883 188395 176949 188396
rect 176147 187780 176213 187781
rect 176147 187716 176148 187780
rect 176212 187716 176213 187780
rect 176147 187715 176213 187716
rect 175782 93810 176210 93870
rect 176150 86970 176210 93810
rect 175782 86910 176210 86970
rect 175595 79932 175661 79933
rect 175595 79868 175596 79932
rect 175660 79868 175661 79932
rect 175595 79867 175661 79868
rect 175595 79796 175661 79797
rect 175595 79732 175596 79796
rect 175660 79732 175661 79796
rect 175595 79731 175661 79732
rect 175411 79388 175477 79389
rect 175411 79324 175412 79388
rect 175476 79324 175477 79388
rect 175411 79323 175477 79324
rect 175598 71637 175658 79731
rect 175782 79389 175842 86910
rect 175963 79796 176029 79797
rect 175963 79732 175964 79796
rect 176028 79732 176029 79796
rect 176331 79796 176397 79797
rect 176331 79794 176332 79796
rect 175963 79731 176029 79732
rect 176150 79734 176332 79794
rect 175779 79388 175845 79389
rect 175779 79324 175780 79388
rect 175844 79324 175845 79388
rect 175779 79323 175845 79324
rect 175966 77349 176026 79731
rect 175963 77348 176029 77349
rect 175963 77284 175964 77348
rect 176028 77284 176029 77348
rect 175963 77283 176029 77284
rect 175963 77212 176029 77213
rect 175963 77148 175964 77212
rect 176028 77148 176029 77212
rect 175963 77147 176029 77148
rect 175595 71636 175661 71637
rect 175595 71572 175596 71636
rect 175660 71572 175661 71636
rect 175595 71571 175661 71572
rect 174862 70350 175106 70410
rect 174862 64565 174922 70350
rect 174859 64564 174925 64565
rect 174859 64500 174860 64564
rect 174924 64500 174925 64564
rect 174859 64499 174925 64500
rect 175966 62797 176026 77147
rect 175963 62796 176029 62797
rect 175963 62732 175964 62796
rect 176028 62732 176029 62796
rect 175963 62731 176029 62732
rect 176150 61573 176210 79734
rect 176331 79732 176332 79734
rect 176396 79732 176397 79796
rect 176331 79731 176397 79732
rect 176518 79661 176578 188395
rect 176699 188324 176765 188325
rect 176699 188260 176700 188324
rect 176764 188260 176765 188324
rect 176699 188259 176765 188260
rect 176702 79933 176762 188259
rect 176699 79932 176765 79933
rect 176699 79868 176700 79932
rect 176764 79868 176765 79932
rect 176699 79867 176765 79868
rect 176886 79797 176946 188395
rect 177294 178954 177914 198000
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 177619 141676 177685 141677
rect 177619 141612 177620 141676
rect 177684 141612 177685 141676
rect 177619 141611 177685 141612
rect 177435 141268 177501 141269
rect 177435 141204 177436 141268
rect 177500 141204 177501 141268
rect 177435 141203 177501 141204
rect 177438 80749 177498 141203
rect 177251 80748 177317 80749
rect 177251 80684 177252 80748
rect 177316 80684 177317 80748
rect 177251 80683 177317 80684
rect 177435 80748 177501 80749
rect 177435 80684 177436 80748
rect 177500 80684 177501 80748
rect 177435 80683 177501 80684
rect 177254 80341 177314 80683
rect 177251 80340 177317 80341
rect 177251 80276 177252 80340
rect 177316 80276 177317 80340
rect 177251 80275 177317 80276
rect 177622 79933 177682 141611
rect 177619 79932 177685 79933
rect 177619 79868 177620 79932
rect 177684 79868 177685 79932
rect 177619 79867 177685 79868
rect 176883 79796 176949 79797
rect 176883 79732 176884 79796
rect 176948 79732 176949 79796
rect 176883 79731 176949 79732
rect 176515 79660 176581 79661
rect 176515 79596 176516 79660
rect 176580 79596 176581 79660
rect 176515 79595 176581 79596
rect 177067 79252 177133 79253
rect 177067 79188 177068 79252
rect 177132 79188 177133 79252
rect 177067 79187 177133 79188
rect 176515 77076 176581 77077
rect 176515 77012 176516 77076
rect 176580 77012 176581 77076
rect 176515 77011 176581 77012
rect 176331 75172 176397 75173
rect 176331 75108 176332 75172
rect 176396 75108 176397 75172
rect 176331 75107 176397 75108
rect 176147 61572 176213 61573
rect 176147 61508 176148 61572
rect 176212 61508 176213 61572
rect 176147 61507 176213 61508
rect 174491 57220 174557 57221
rect 174491 57156 174492 57220
rect 174556 57156 174557 57220
rect 174491 57155 174557 57156
rect 173755 47972 173821 47973
rect 173755 47908 173756 47972
rect 173820 47908 173821 47972
rect 173755 47907 173821 47908
rect 176334 44981 176394 75107
rect 176331 44980 176397 44981
rect 176331 44916 176332 44980
rect 176396 44916 176397 44980
rect 176331 44915 176397 44916
rect 176518 44845 176578 77011
rect 177070 50285 177130 79187
rect 178174 78437 178234 199003
rect 178358 78709 178418 199955
rect 179459 197844 179525 197845
rect 179459 197780 179460 197844
rect 179524 197780 179525 197844
rect 179459 197779 179525 197780
rect 178539 187100 178605 187101
rect 178539 187036 178540 187100
rect 178604 187036 178605 187100
rect 178539 187035 178605 187036
rect 178542 80749 178602 187035
rect 178723 140180 178789 140181
rect 178723 140116 178724 140180
rect 178788 140116 178789 140180
rect 178723 140115 178789 140116
rect 178539 80748 178605 80749
rect 178539 80684 178540 80748
rect 178604 80684 178605 80748
rect 178539 80683 178605 80684
rect 178355 78708 178421 78709
rect 178355 78644 178356 78708
rect 178420 78644 178421 78708
rect 178355 78643 178421 78644
rect 178171 78436 178237 78437
rect 178171 78372 178172 78436
rect 178236 78372 178237 78436
rect 178171 78371 178237 78372
rect 177294 70954 177914 78000
rect 178726 75037 178786 140115
rect 179462 76397 179522 197779
rect 179643 197572 179709 197573
rect 179643 197508 179644 197572
rect 179708 197508 179709 197572
rect 179643 197507 179709 197508
rect 179646 77349 179706 197507
rect 180750 195990 180810 200499
rect 180931 199612 180997 199613
rect 180931 199548 180932 199612
rect 180996 199548 180997 199612
rect 180931 199547 180997 199548
rect 180566 195930 180810 195990
rect 180566 157350 180626 195930
rect 180566 157290 180810 157350
rect 180750 147690 180810 157290
rect 180566 147630 180810 147690
rect 179827 146980 179893 146981
rect 179827 146916 179828 146980
rect 179892 146916 179893 146980
rect 179827 146915 179893 146916
rect 179643 77348 179709 77349
rect 179643 77284 179644 77348
rect 179708 77284 179709 77348
rect 179643 77283 179709 77284
rect 179830 77213 179890 146915
rect 180011 140044 180077 140045
rect 180011 139980 180012 140044
rect 180076 139980 180077 140044
rect 180011 139979 180077 139980
rect 180014 81021 180074 139979
rect 180566 89730 180626 147630
rect 180566 89670 180810 89730
rect 180011 81020 180077 81021
rect 180011 80956 180012 81020
rect 180076 80956 180077 81020
rect 180011 80955 180077 80956
rect 179827 77212 179893 77213
rect 179827 77148 179828 77212
rect 179892 77148 179893 77212
rect 179827 77147 179893 77148
rect 179459 76396 179525 76397
rect 179459 76332 179460 76396
rect 179524 76332 179525 76396
rect 179459 76331 179525 76332
rect 178723 75036 178789 75037
rect 178723 74972 178724 75036
rect 178788 74972 178789 75036
rect 178723 74971 178789 74972
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177067 50284 177133 50285
rect 177067 50220 177068 50284
rect 177132 50220 177133 50284
rect 177067 50219 177133 50220
rect 176515 44844 176581 44845
rect 176515 44780 176516 44844
rect 176580 44780 176581 44844
rect 176515 44779 176581 44780
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 179462 68373 179522 76331
rect 180750 70410 180810 89670
rect 180934 71773 180994 199547
rect 182587 199340 182653 199341
rect 182587 199276 182588 199340
rect 182652 199276 182653 199340
rect 182587 199275 182653 199276
rect 181794 183454 182414 198000
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181115 149564 181181 149565
rect 181115 149500 181116 149564
rect 181180 149500 181181 149564
rect 181115 149499 181181 149500
rect 181118 73949 181178 149499
rect 181794 147454 182414 182898
rect 181299 147252 181365 147253
rect 181299 147188 181300 147252
rect 181364 147188 181365 147252
rect 181299 147187 181365 147188
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181302 77213 181362 147187
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 181667 140044 181733 140045
rect 181667 139980 181668 140044
rect 181732 139980 181733 140044
rect 181667 139979 181733 139980
rect 181670 138821 181730 139979
rect 181667 138820 181733 138821
rect 181667 138756 181668 138820
rect 181732 138756 181733 138820
rect 181667 138755 181733 138756
rect 182590 80749 182650 199275
rect 183507 199204 183573 199205
rect 183507 199140 183508 199204
rect 183572 199140 183573 199204
rect 183507 199139 183573 199140
rect 182771 150380 182837 150381
rect 182771 150316 182772 150380
rect 182836 150316 182837 150380
rect 182771 150315 182837 150316
rect 182587 80748 182653 80749
rect 182587 80684 182588 80748
rect 182652 80684 182653 80748
rect 182587 80683 182653 80684
rect 181299 77212 181365 77213
rect 181299 77148 181300 77212
rect 181364 77148 181365 77212
rect 181299 77147 181365 77148
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181115 73948 181181 73949
rect 181115 73884 181116 73948
rect 181180 73884 181181 73948
rect 181115 73883 181181 73884
rect 180931 71772 180997 71773
rect 180931 71708 180932 71772
rect 180996 71708 180997 71772
rect 180931 71707 180997 71708
rect 180566 70350 180810 70410
rect 179459 68372 179525 68373
rect 179459 68308 179460 68372
rect 179524 68308 179525 68372
rect 179459 68307 179525 68308
rect 180566 61981 180626 70350
rect 180563 61980 180629 61981
rect 180563 61916 180564 61980
rect 180628 61916 180629 61980
rect 180563 61915 180629 61916
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 74898
rect 182774 72725 182834 150315
rect 182955 147388 183021 147389
rect 182955 147324 182956 147388
rect 183020 147324 183021 147388
rect 182955 147323 183021 147324
rect 182958 74085 183018 147323
rect 182955 74084 183021 74085
rect 182955 74020 182956 74084
rect 183020 74020 183021 74084
rect 182955 74019 183021 74020
rect 182771 72724 182837 72725
rect 182771 72660 182772 72724
rect 182836 72660 182837 72724
rect 182771 72659 182837 72660
rect 183510 70410 183570 199139
rect 183691 198932 183757 198933
rect 183691 198868 183692 198932
rect 183756 198868 183757 198932
rect 183691 198867 183757 198868
rect 183694 76261 183754 198867
rect 184979 198796 185045 198797
rect 184979 198732 184980 198796
rect 185044 198732 185045 198796
rect 184979 198731 185045 198732
rect 183875 150244 183941 150245
rect 183875 150180 183876 150244
rect 183940 150180 183941 150244
rect 183875 150179 183941 150180
rect 183691 76260 183757 76261
rect 183691 76196 183692 76260
rect 183756 76196 183757 76260
rect 183691 76195 183757 76196
rect 183694 71365 183754 76195
rect 183878 73133 183938 150179
rect 184059 149836 184125 149837
rect 184059 149772 184060 149836
rect 184124 149772 184125 149836
rect 184059 149771 184125 149772
rect 184062 74221 184122 149771
rect 184982 80341 185042 198731
rect 187003 198524 187069 198525
rect 187003 198460 187004 198524
rect 187068 198460 187069 198524
rect 187003 198459 187069 198460
rect 186294 187954 186914 198000
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186083 152556 186149 152557
rect 186083 152492 186084 152556
rect 186148 152492 186149 152556
rect 186083 152491 186149 152492
rect 185163 149972 185229 149973
rect 185163 149908 185164 149972
rect 185228 149908 185229 149972
rect 185163 149907 185229 149908
rect 184979 80340 185045 80341
rect 184979 80276 184980 80340
rect 185044 80276 185045 80340
rect 184979 80275 185045 80276
rect 184059 74220 184125 74221
rect 184059 74156 184060 74220
rect 184124 74156 184125 74220
rect 184059 74155 184125 74156
rect 183875 73132 183941 73133
rect 183875 73068 183876 73132
rect 183940 73068 183941 73132
rect 183875 73067 183941 73068
rect 185166 72997 185226 149907
rect 185347 149700 185413 149701
rect 185347 149636 185348 149700
rect 185412 149636 185413 149700
rect 185347 149635 185413 149636
rect 185350 75581 185410 149635
rect 185899 140180 185965 140181
rect 185899 140116 185900 140180
rect 185964 140116 185965 140180
rect 185899 140115 185965 140116
rect 185902 138957 185962 140115
rect 185899 138956 185965 138957
rect 185899 138892 185900 138956
rect 185964 138892 185965 138956
rect 185899 138891 185965 138892
rect 186086 138005 186146 152491
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 186083 138004 186149 138005
rect 186083 137940 186084 138004
rect 186148 137940 186149 138004
rect 186083 137939 186149 137940
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 185347 75580 185413 75581
rect 185347 75516 185348 75580
rect 185412 75516 185413 75580
rect 185347 75515 185413 75516
rect 185163 72996 185229 72997
rect 185163 72932 185164 72996
rect 185228 72932 185229 72996
rect 185163 72931 185229 72932
rect 183691 71364 183757 71365
rect 183691 71300 183692 71364
rect 183756 71300 183757 71364
rect 183691 71299 183757 71300
rect 183510 70350 183754 70410
rect 183694 58989 183754 70350
rect 183691 58988 183757 58989
rect 183691 58924 183692 58988
rect 183756 58924 183757 58988
rect 183691 58923 183757 58924
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187006 76533 187066 198459
rect 187187 195668 187253 195669
rect 187187 195604 187188 195668
rect 187252 195604 187253 195668
rect 187187 195603 187253 195604
rect 187190 79389 187250 195603
rect 187374 194853 187434 284275
rect 189027 278084 189093 278085
rect 189027 278020 189028 278084
rect 189092 278020 189093 278084
rect 189027 278019 189093 278020
rect 189030 277541 189090 278019
rect 189027 277540 189093 277541
rect 189027 277476 189028 277540
rect 189092 277476 189093 277540
rect 189027 277475 189093 277476
rect 187739 276044 187805 276045
rect 187739 275980 187740 276044
rect 187804 275980 187805 276044
rect 187739 275979 187805 275980
rect 187371 194852 187437 194853
rect 187371 194788 187372 194852
rect 187436 194788 187437 194852
rect 187371 194787 187437 194788
rect 187742 142901 187802 275979
rect 187923 262308 187989 262309
rect 187923 262244 187924 262308
rect 187988 262244 187989 262308
rect 187923 262243 187989 262244
rect 187926 144397 187986 262243
rect 188107 259996 188173 259997
rect 188107 259932 188108 259996
rect 188172 259932 188173 259996
rect 188107 259931 188173 259932
rect 187923 144396 187989 144397
rect 187923 144332 187924 144396
rect 187988 144332 187989 144396
rect 187923 144331 187989 144332
rect 188110 143309 188170 259931
rect 188291 259860 188357 259861
rect 188291 259796 188292 259860
rect 188356 259796 188357 259860
rect 188291 259795 188357 259796
rect 188107 143308 188173 143309
rect 188107 143244 188108 143308
rect 188172 143244 188173 143308
rect 188107 143243 188173 143244
rect 188294 143173 188354 259795
rect 188291 143172 188357 143173
rect 188291 143108 188292 143172
rect 188356 143108 188357 143172
rect 188291 143107 188357 143108
rect 187739 142900 187805 142901
rect 187739 142836 187740 142900
rect 187804 142836 187805 142900
rect 187739 142835 187805 142836
rect 189030 142765 189090 277475
rect 190794 264454 191414 299898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 193259 265300 193325 265301
rect 193259 265236 193260 265300
rect 193324 265236 193325 265300
rect 193259 265235 193325 265236
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 262000 191414 263898
rect 192155 262580 192221 262581
rect 192155 262516 192156 262580
rect 192220 262516 192221 262580
rect 192155 262515 192221 262516
rect 191971 262444 192037 262445
rect 191971 262380 191972 262444
rect 192036 262380 192037 262444
rect 191971 262379 192037 262380
rect 189395 260132 189461 260133
rect 189395 260068 189396 260132
rect 189460 260068 189461 260132
rect 189395 260067 189461 260068
rect 189211 198660 189277 198661
rect 189211 198596 189212 198660
rect 189276 198596 189277 198660
rect 189211 198595 189277 198596
rect 189027 142764 189093 142765
rect 189027 142700 189028 142764
rect 189092 142700 189093 142764
rect 189027 142699 189093 142700
rect 188291 141132 188357 141133
rect 188291 141068 188292 141132
rect 188356 141068 188357 141132
rect 188291 141067 188357 141068
rect 187739 139772 187805 139773
rect 187739 139708 187740 139772
rect 187804 139708 187805 139772
rect 187739 139707 187805 139708
rect 187187 79388 187253 79389
rect 187187 79324 187188 79388
rect 187252 79324 187253 79388
rect 187187 79323 187253 79324
rect 187742 79253 187802 139707
rect 188294 111893 188354 141067
rect 189027 140180 189093 140181
rect 189027 140116 189028 140180
rect 189092 140116 189093 140180
rect 189027 140115 189093 140116
rect 188659 140044 188725 140045
rect 188659 139980 188660 140044
rect 188724 139980 188725 140044
rect 188659 139979 188725 139980
rect 188662 125629 188722 139979
rect 188659 125628 188725 125629
rect 188659 125564 188660 125628
rect 188724 125564 188725 125628
rect 188659 125563 188725 125564
rect 188291 111892 188357 111893
rect 188291 111828 188292 111892
rect 188356 111828 188357 111892
rect 188291 111827 188357 111828
rect 187739 79252 187805 79253
rect 187739 79188 187740 79252
rect 187804 79188 187805 79252
rect 187739 79187 187805 79188
rect 187003 76532 187069 76533
rect 187003 76468 187004 76532
rect 187068 76468 187069 76532
rect 187003 76467 187069 76468
rect 187555 76532 187621 76533
rect 187555 76468 187556 76532
rect 187620 76468 187621 76532
rect 187555 76467 187621 76468
rect 187558 71773 187618 76467
rect 189030 75445 189090 140115
rect 189027 75444 189093 75445
rect 189027 75380 189028 75444
rect 189092 75380 189093 75444
rect 189027 75379 189093 75380
rect 187555 71772 187621 71773
rect 187555 71708 187556 71772
rect 187620 71708 187621 71772
rect 187555 71707 187621 71708
rect 189214 71093 189274 198595
rect 189398 141405 189458 260067
rect 189579 259724 189645 259725
rect 189579 259660 189580 259724
rect 189644 259660 189645 259724
rect 189579 259659 189645 259660
rect 189582 142085 189642 259659
rect 190499 198388 190565 198389
rect 190499 198324 190500 198388
rect 190564 198324 190565 198388
rect 190499 198323 190565 198324
rect 189579 142084 189645 142085
rect 189579 142020 189580 142084
rect 189644 142020 189645 142084
rect 189579 142019 189645 142020
rect 189395 141404 189461 141405
rect 189395 141340 189396 141404
rect 189460 141340 189461 141404
rect 189395 141339 189461 141340
rect 189763 140996 189829 140997
rect 189763 140932 189764 140996
rect 189828 140932 189829 140996
rect 189763 140931 189829 140932
rect 189211 71092 189277 71093
rect 189211 71028 189212 71092
rect 189276 71028 189277 71092
rect 189211 71027 189277 71028
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 189766 31789 189826 140931
rect 190315 75444 190381 75445
rect 190315 75380 190316 75444
rect 190380 75380 190381 75444
rect 190315 75379 190381 75380
rect 190318 71773 190378 75379
rect 190315 71772 190381 71773
rect 190315 71708 190316 71772
rect 190380 71708 190381 71772
rect 190315 71707 190381 71708
rect 190502 71229 190562 198323
rect 190794 192454 191414 198000
rect 191787 195532 191853 195533
rect 191787 195468 191788 195532
rect 191852 195468 191853 195532
rect 191787 195467 191853 195468
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 142000 191414 155898
rect 191603 142220 191669 142221
rect 191603 142156 191604 142220
rect 191668 142156 191669 142220
rect 191603 142155 191669 142156
rect 190683 140452 190749 140453
rect 190683 140388 190684 140452
rect 190748 140388 190749 140452
rect 190683 140387 190749 140388
rect 190686 78981 190746 140387
rect 191606 79389 191666 142155
rect 191603 79388 191669 79389
rect 191603 79324 191604 79388
rect 191668 79324 191669 79388
rect 191603 79323 191669 79324
rect 190683 78980 190749 78981
rect 190683 78916 190684 78980
rect 190748 78916 190749 78980
rect 190683 78915 190749 78916
rect 190499 71228 190565 71229
rect 190499 71164 190500 71228
rect 190564 71164 190565 71228
rect 190499 71163 190565 71164
rect 190794 48454 191414 78000
rect 191790 64157 191850 195467
rect 191974 141541 192034 262379
rect 192158 143989 192218 262515
rect 192339 262308 192405 262309
rect 192339 262244 192340 262308
rect 192404 262244 192405 262308
rect 192339 262243 192405 262244
rect 192342 144125 192402 262243
rect 193262 145757 193322 265235
rect 194731 265164 194797 265165
rect 194731 265100 194732 265164
rect 194796 265100 194797 265164
rect 194731 265099 194797 265100
rect 193443 262716 193509 262717
rect 193443 262652 193444 262716
rect 193508 262652 193509 262716
rect 193443 262651 193509 262652
rect 193259 145756 193325 145757
rect 193259 145692 193260 145756
rect 193324 145692 193325 145756
rect 193259 145691 193325 145692
rect 193446 144533 193506 262651
rect 193627 260948 193693 260949
rect 193627 260884 193628 260948
rect 193692 260884 193693 260948
rect 193627 260883 193693 260884
rect 193443 144532 193509 144533
rect 193443 144468 193444 144532
rect 193508 144468 193509 144532
rect 193443 144467 193509 144468
rect 193630 144261 193690 260883
rect 194547 198252 194613 198253
rect 194547 198188 194548 198252
rect 194612 198188 194613 198252
rect 194547 198187 194613 198188
rect 193995 146300 194061 146301
rect 193995 146236 193996 146300
rect 194060 146236 194061 146300
rect 193995 146235 194061 146236
rect 193811 146164 193877 146165
rect 193811 146100 193812 146164
rect 193876 146100 193877 146164
rect 193811 146099 193877 146100
rect 193627 144260 193693 144261
rect 193627 144196 193628 144260
rect 193692 144196 193693 144260
rect 193627 144195 193693 144196
rect 192339 144124 192405 144125
rect 192339 144060 192340 144124
rect 192404 144060 192405 144124
rect 192339 144059 192405 144060
rect 192155 143988 192221 143989
rect 192155 143924 192156 143988
rect 192220 143924 192221 143988
rect 192155 143923 192221 143924
rect 191971 141540 192037 141541
rect 191971 141476 191972 141540
rect 192036 141476 192037 141540
rect 191971 141475 192037 141476
rect 192339 140860 192405 140861
rect 192339 140796 192340 140860
rect 192404 140796 192405 140860
rect 192339 140795 192405 140796
rect 191971 139908 192037 139909
rect 191971 139844 191972 139908
rect 192036 139844 192037 139908
rect 191971 139843 192037 139844
rect 191974 79117 192034 139843
rect 191971 79116 192037 79117
rect 191971 79052 191972 79116
rect 192036 79052 192037 79116
rect 191971 79051 192037 79052
rect 191787 64156 191853 64157
rect 191787 64092 191788 64156
rect 191852 64092 191853 64156
rect 191787 64091 191853 64092
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 189763 31788 189829 31789
rect 189763 31724 189764 31788
rect 189828 31724 189829 31788
rect 189763 31723 189829 31724
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 12454 191414 47898
rect 192342 45661 192402 140795
rect 193814 65517 193874 146099
rect 193998 66197 194058 146235
rect 194550 69597 194610 198187
rect 194734 145893 194794 265099
rect 195294 232954 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 196203 265436 196269 265437
rect 196203 265372 196204 265436
rect 196268 265372 196269 265436
rect 196203 265371 196269 265372
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 196019 179348 196085 179349
rect 196019 179284 196020 179348
rect 196084 179284 196085 179348
rect 196019 179283 196085 179284
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 194731 145892 194797 145893
rect 194731 145828 194732 145892
rect 194796 145828 194797 145892
rect 194731 145827 194797 145828
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 194547 69596 194613 69597
rect 194547 69532 194548 69596
rect 194612 69532 194613 69596
rect 194547 69531 194613 69532
rect 193995 66196 194061 66197
rect 193995 66132 193996 66196
rect 194060 66132 194061 66196
rect 193995 66131 194061 66132
rect 193811 65516 193877 65517
rect 193811 65452 193812 65516
rect 193876 65452 193877 65516
rect 193811 65451 193877 65452
rect 195294 52954 195914 88398
rect 196022 68917 196082 179283
rect 196206 144805 196266 265371
rect 197491 265028 197557 265029
rect 197491 264964 197492 265028
rect 197556 264964 197557 265028
rect 197491 264963 197557 264964
rect 196571 198660 196637 198661
rect 196571 198596 196572 198660
rect 196636 198596 196637 198660
rect 196571 198595 196637 198596
rect 196203 144804 196269 144805
rect 196203 144740 196204 144804
rect 196268 144740 196269 144804
rect 196203 144739 196269 144740
rect 196574 80069 196634 198595
rect 197307 197028 197373 197029
rect 197307 196964 197308 197028
rect 197372 196964 197373 197028
rect 197307 196963 197373 196964
rect 196571 80068 196637 80069
rect 196571 80004 196572 80068
rect 196636 80004 196637 80068
rect 196571 80003 196637 80004
rect 196019 68916 196085 68917
rect 196019 68852 196020 68916
rect 196084 68852 196085 68916
rect 196019 68851 196085 68852
rect 197310 61573 197370 196963
rect 197494 144669 197554 264963
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 198779 188052 198845 188053
rect 198779 187988 198780 188052
rect 198844 187988 198845 188052
rect 198779 187987 198845 187988
rect 197859 147796 197925 147797
rect 197859 147732 197860 147796
rect 197924 147732 197925 147796
rect 197859 147731 197925 147732
rect 197491 144668 197557 144669
rect 197491 144604 197492 144668
rect 197556 144604 197557 144668
rect 197491 144603 197557 144604
rect 197862 62933 197922 147731
rect 197859 62932 197925 62933
rect 197859 62868 197860 62932
rect 197924 62868 197925 62932
rect 197859 62867 197925 62868
rect 198782 62797 198842 187987
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 200619 199748 200685 199749
rect 200619 199684 200620 199748
rect 200684 199684 200685 199748
rect 200619 199683 200685 199684
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199331 146300 199397 146301
rect 199331 146236 199332 146300
rect 199396 146236 199397 146300
rect 199331 146235 199397 146236
rect 199334 70413 199394 146235
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199331 70412 199397 70413
rect 199331 70348 199332 70412
rect 199396 70348 199397 70412
rect 199331 70347 199397 70348
rect 198779 62796 198845 62797
rect 198779 62732 198780 62796
rect 198844 62732 198845 62796
rect 198779 62731 198845 62732
rect 197307 61572 197373 61573
rect 197307 61508 197308 61572
rect 197372 61508 197373 61572
rect 197307 61507 197373 61508
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 192339 45660 192405 45661
rect 192339 45596 192340 45660
rect 192404 45596 192405 45660
rect 192339 45595 192405 45596
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 200622 56541 200682 199683
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 201723 150380 201789 150381
rect 201723 150316 201724 150380
rect 201788 150316 201789 150380
rect 201723 150315 201789 150316
rect 203011 150380 203077 150381
rect 203011 150316 203012 150380
rect 203076 150316 203077 150380
rect 203011 150315 203077 150316
rect 201539 150108 201605 150109
rect 201539 150044 201540 150108
rect 201604 150044 201605 150108
rect 201539 150043 201605 150044
rect 200803 138140 200869 138141
rect 200803 138076 200804 138140
rect 200868 138076 200869 138140
rect 200803 138075 200869 138076
rect 200806 67557 200866 138075
rect 201542 74357 201602 150043
rect 201726 77621 201786 150315
rect 202827 147116 202893 147117
rect 202827 147052 202828 147116
rect 202892 147052 202893 147116
rect 202827 147051 202893 147052
rect 202830 84210 202890 147051
rect 203014 93870 203074 150315
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 203014 93810 203258 93870
rect 202830 84150 203074 84210
rect 201723 77620 201789 77621
rect 201723 77556 201724 77620
rect 201788 77556 201789 77620
rect 201723 77555 201789 77556
rect 201539 74356 201605 74357
rect 201539 74292 201540 74356
rect 201604 74292 201605 74356
rect 201539 74291 201605 74292
rect 200803 67556 200869 67557
rect 200803 67492 200804 67556
rect 200868 67492 200869 67556
rect 200803 67491 200869 67492
rect 200619 56540 200685 56541
rect 200619 56476 200620 56540
rect 200684 56476 200685 56540
rect 200619 56475 200685 56476
rect 203014 47973 203074 84150
rect 203198 78029 203258 93810
rect 203195 78028 203261 78029
rect 203195 77964 203196 78028
rect 203260 77964 203261 78028
rect 203195 77963 203261 77964
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 203011 47972 203077 47973
rect 203011 47908 203012 47972
rect 203076 47908 203077 47972
rect 203011 47907 203077 47908
rect 204115 47972 204181 47973
rect 204115 47908 204116 47972
rect 204180 47908 204181 47972
rect 204115 47907 204181 47908
rect 204118 47565 204178 47907
rect 204115 47564 204181 47565
rect 204115 47500 204116 47564
rect 204180 47500 204181 47564
rect 204115 47499 204181 47500
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 1066 0 68854 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 68854 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
